library IEEE;use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity ROM is
generic(
   width : natural := 24
);
port(
   dir  : in std_logic_vector(width-1 downto 0);
   data : out std_logic_vector(width-1 downto 0)
);
end ROM;
architecture Behavioral of ROM is
type srom is array (0 to 2**width-1) of integer range 2**width - 1 downto 0;
signal srom_1 : srom;
begin
data <= std_logic_vector(to_signed(srom_1(to_integer(unsigned(dir))),width));
srom_1(0) <= 8388607;
srom_1(1) <= 8962711;
srom_1(2) <= 9534124;
srom_1(3) <= 10100165;
srom_1(4) <= 10658180;
srom_1(5) <= 11205552;
srom_1(6) <= 11739714;
srom_1(7) <= 12258162;
srom_1(8) <= 12758464;
srom_1(9) <= 13238274;
srom_1(10) <= 13695343;
srom_1(11) <= 14127527;
srom_1(12) <= 14532798;
srom_1(13) <= 14909258;
srom_1(14) <= 15255140;
srom_1(15) <= 15568822;
srom_1(16) <= 15848834;
srom_1(17) <= 16093863;
srom_1(18) <= 16302758;
srom_1(19) <= 16474542;
srom_1(20) <= 16608408;
srom_1(21) <= 16703728;
srom_1(22) <= 16760056;
srom_1(23) <= 16777128;
srom_1(24) <= 16754862;
srom_1(25) <= 16693365;
srom_1(26) <= 16592923;
srom_1(27) <= 16454009;
srom_1(28) <= 16277273;
srom_1(29) <= 16063545;
srom_1(30) <= 15813826;
srom_1(31) <= 15529288;
srom_1(32) <= 15211265;
srom_1(33) <= 14861247;
srom_1(34) <= 14480878;
srom_1(35) <= 14071940;
srom_1(36) <= 13636350;
srom_1(37) <= 13176152;
srom_1(38) <= 12693504;
srom_1(39) <= 12190668;
srom_1(40) <= 11670004;
srom_1(41) <= 11133951;
srom_1(42) <= 10585025;
srom_1(43) <= 10025799;
srom_1(44) <= 9458896;
srom_1(45) <= 8886974;
srom_1(46) <= 8312715;
srom_1(47) <= 7738811;
srom_1(48) <= 7167955;
srom_1(49) <= 6602823;
srom_1(50) <= 6046065;
srom_1(51) <= 5500292;
srom_1(52) <= 4968063;
srom_1(53) <= 4451875;
srom_1(54) <= 3954147;
srom_1(55) <= 3477213;
srom_1(56) <= 3023311;
srom_1(57) <= 2594569;
srom_1(58) <= 2192997;
srom_1(59) <= 1820478;
srom_1(60) <= 1478760;
srom_1(61) <= 1169444;
srom_1(62) <= 893981;
srom_1(63) <= 653663;
srom_1(64) <= 449617;
srom_1(65) <= 282800;
srom_1(66) <= 153993;
srom_1(67) <= 63802;
srom_1(68) <= 12648;
srom_1(69) <= 772;
srom_1(70) <= 28229;
srom_1(71) <= 94892;
srom_1(72) <= 200446;
srom_1(73) <= 344397;
srom_1(74) <= 526070;
srom_1(75) <= 744614;
srom_1(76) <= 999003;
srom_1(77) <= 1288044;
srom_1(78) <= 1610382;
srom_1(79) <= 1964506;
srom_1(80) <= 2348754;
srom_1(81) <= 2761326;
srom_1(82) <= 3200285;
srom_1(83) <= 3663575;
srom_1(84) <= 4149022;
srom_1(85) <= 4654349;
srom_1(86) <= 5177188;
srom_1(87) <= 5715086;
srom_1(88) <= 6265522;
srom_1(89) <= 6825913;
srom_1(90) <= 7393632;
srom_1(91) <= 7966017;
srom_1(92) <= 8540384;
srom_1(93) <= 9114039;
srom_1(94) <= 9684292;
srom_1(95) <= 10248469;
srom_1(96) <= 10803925;
srom_1(97) <= 11348054;
srom_1(98) <= 11878306;
srom_1(99) <= 12392193;
srom_1(100) <= 12887306;
srom_1(101) <= 13361323;
srom_1(102) <= 13812021;
srom_1(103) <= 14237287;
srom_1(104) <= 14635126;
srom_1(105) <= 15003674;
srom_1(106) <= 15341201;
srom_1(107) <= 15646125;
srom_1(108) <= 15917016;
srom_1(109) <= 16152604;
srom_1(110) <= 16351783;
srom_1(111) <= 16513621;
srom_1(112) <= 16637358;
srom_1(113) <= 16722413;
srom_1(114) <= 16768388;
srom_1(115) <= 16775068;
srom_1(116) <= 16742421;
srom_1(117) <= 16670599;
srom_1(118) <= 16559941;
srom_1(119) <= 16410964;
srom_1(120) <= 16224368;
srom_1(121) <= 16001027;
srom_1(122) <= 15741989;
srom_1(123) <= 15448469;
srom_1(124) <= 15121842;
srom_1(125) <= 14763641;
srom_1(126) <= 14375545;
srom_1(127) <= 13959375;
srom_1(128) <= 13517081;
srom_1(129) <= 13050738;
srom_1(130) <= 12562532;
srom_1(131) <= 12054754;
srom_1(132) <= 11529783;
srom_1(133) <= 10990083;
srom_1(134) <= 10438184;
srom_1(135) <= 9876673;
srom_1(136) <= 9308184;
srom_1(137) <= 8735383;
srom_1(138) <= 8160956;
srom_1(139) <= 7587597;
srom_1(140) <= 7017993;
srom_1(141) <= 6454817;
srom_1(142) <= 5900709;
srom_1(143) <= 5358268;
srom_1(144) <= 4830037;
srom_1(145) <= 4318494;
srom_1(146) <= 3826036;
srom_1(147) <= 3354974;
srom_1(148) <= 2907517;
srom_1(149) <= 2485762;
srom_1(150) <= 2091687;
srom_1(151) <= 1727141;
srom_1(152) <= 1393833;
srom_1(153) <= 1093326;
srom_1(154) <= 827029;
srom_1(155) <= 596191;
srom_1(156) <= 401894;
srom_1(157) <= 245049;
srom_1(158) <= 126393;
srom_1(159) <= 46480;
srom_1(160) <= 5687;
srom_1(161) <= 4205;
srom_1(162) <= 42039;
srom_1(163) <= 119014;
srom_1(164) <= 234767;
srom_1(165) <= 388757;
srom_1(166) <= 580261;
srom_1(167) <= 808380;
srom_1(168) <= 1072046;
srom_1(169) <= 1370022;
srom_1(170) <= 1700911;
srom_1(171) <= 2063160;
srom_1(172) <= 2455071;
srom_1(173) <= 2874807;
srom_1(174) <= 3320399;
srom_1(175) <= 3789758;
srom_1(176) <= 4280682;
srom_1(177) <= 4790870;
srom_1(178) <= 5317928;
srom_1(179) <= 5859386;
srom_1(180) <= 6412705;
srom_1(181) <= 6975289;
srom_1(182) <= 7544501;
srom_1(183) <= 8117671;
srom_1(184) <= 8692111;
srom_1(185) <= 9265128;
srom_1(186) <= 9834035;
srom_1(187) <= 10396164;
srom_1(188) <= 10948879;
srom_1(189) <= 11489588;
srom_1(190) <= 12015755;
srom_1(191) <= 12524913;
srom_1(192) <= 13014675;
srom_1(193) <= 13482743;
srom_1(194) <= 13926923;
srom_1(195) <= 14345133;
srom_1(196) <= 14735410;
srom_1(197) <= 15095924;
srom_1(198) <= 15424986;
srom_1(199) <= 15721052;
srom_1(200) <= 15982733;
srom_1(201) <= 16208803;
srom_1(202) <= 16398201;
srom_1(203) <= 16550040;
srom_1(204) <= 16663607;
srom_1(205) <= 16738369;
srom_1(206) <= 16773977;
srom_1(207) <= 16770263;
srom_1(208) <= 16727244;
srom_1(209) <= 16645122;
srom_1(210) <= 16524283;
srom_1(211) <= 16365293;
srom_1(212) <= 16168898;
srom_1(213) <= 15936018;
srom_1(214) <= 15667745;
srom_1(215) <= 15365338;
srom_1(216) <= 15030215;
srom_1(217) <= 14663947;
srom_1(218) <= 14268252;
srom_1(219) <= 13844986;
srom_1(220) <= 13396132;
srom_1(221) <= 12923796;
srom_1(222) <= 12430194;
srom_1(223) <= 11917639;
srom_1(224) <= 11388535;
srom_1(225) <= 10845363;
srom_1(226) <= 10290671;
srom_1(227) <= 9727059;
srom_1(228) <= 9157171;
srom_1(229) <= 8583679;
srom_1(230) <= 8009272;
srom_1(231) <= 7436644;
srom_1(232) <= 6868480;
srom_1(233) <= 6307445;
srom_1(234) <= 5756168;
srom_1(235) <= 5217236;
srom_1(236) <= 4693176;
srom_1(237) <= 4186445;
srom_1(238) <= 3699419;
srom_1(239) <= 3234383;
srom_1(240) <= 2793516;
srom_1(241) <= 2378887;
srom_1(242) <= 1992439;
srom_1(243) <= 1635985;
srom_1(244) <= 1311197;
srom_1(245) <= 1019597;
srom_1(246) <= 762553;
srom_1(247) <= 541269;
srom_1(248) <= 356785;
srom_1(249) <= 209965;
srom_1(250) <= 101497;
srom_1(251) <= 31891;
srom_1(252) <= 1471;
srom_1(253) <= 10382;
srom_1(254) <= 58582;
srom_1(255) <= 145843;
srom_1(256) <= 271758;
srom_1(257) <= 435736;
srom_1(258) <= 637007;
srom_1(259) <= 874628;
srom_1(260) <= 1147485;
srom_1(261) <= 1454298;
srom_1(262) <= 1793628;
srom_1(263) <= 2163885;
srom_1(264) <= 2563331;
srom_1(265) <= 2990094;
srom_1(266) <= 3442172;
srom_1(267) <= 3917446;
srom_1(268) <= 4413687;
srom_1(269) <= 4928568;
srom_1(270) <= 5459674;
srom_1(271) <= 6004514;
srom_1(272) <= 6560535;
srom_1(273) <= 7125128;
srom_1(274) <= 7695646;
srom_1(275) <= 8269413;
srom_1(276) <= 8843739;
srom_1(277) <= 9415931;
srom_1(278) <= 9983306;
srom_1(279) <= 10543202;
srom_1(280) <= 11092995;
srom_1(281) <= 11630106;
srom_1(282) <= 12152016;
srom_1(283) <= 12656279;
srom_1(284) <= 13140529;
srom_1(285) <= 13602496;
srom_1(286) <= 14040012;
srom_1(287) <= 14451028;
srom_1(288) <= 14833615;
srom_1(289) <= 15185978;
srom_1(290) <= 15506467;
srom_1(291) <= 15793578;
srom_1(292) <= 16045964;
srom_1(293) <= 16262442;
srom_1(294) <= 16441997;
srom_1(295) <= 16583787;
srom_1(296) <= 16687147;
srom_1(297) <= 16751592;
srom_1(298) <= 16776820;
srom_1(299) <= 16762713;
srom_1(300) <= 16709337;
srom_1(301) <= 16616942;
srom_1(302) <= 16485962;
srom_1(303) <= 16317010;
srom_1(304) <= 16110880;
srom_1(305) <= 15868537;
srom_1(306) <= 15591118;
srom_1(307) <= 15279924;
srom_1(308) <= 14936414;
srom_1(309) <= 14562199;
srom_1(310) <= 14159035;
srom_1(311) <= 13728810;
srom_1(312) <= 13273544;
srom_1(313) <= 12795371;
srom_1(314) <= 12296532;
srom_1(315) <= 11779368;
srom_1(316) <= 11246304;
srom_1(317) <= 10699839;
srom_1(318) <= 10142536;
srom_1(319) <= 9577008;
srom_1(320) <= 9005907;
srom_1(321) <= 8431911;
srom_1(322) <= 7857713;
srom_1(323) <= 7286003;
srom_1(324) <= 6719465;
srom_1(325) <= 6160753;
srom_1(326) <= 5612489;
srom_1(327) <= 5077243;
srom_1(328) <= 4557525;
srom_1(329) <= 4055772;
srom_1(330) <= 3574338;
srom_1(331) <= 3115479;
srom_1(332) <= 2681348;
srom_1(333) <= 2273979;
srom_1(334) <= 1895285;
srom_1(335) <= 1547040;
srom_1(336) <= 1230877;
srom_1(337) <= 948280;
srom_1(338) <= 700573;
srom_1(339) <= 488917;
srom_1(340) <= 314306;
srom_1(341) <= 177558;
srom_1(342) <= 79315;
srom_1(343) <= 20036;
srom_1(344) <= 1;
srom_1(345) <= 19303;
srom_1(346) <= 77851;
srom_1(347) <= 175372;
srom_1(348) <= 311407;
srom_1(349) <= 485318;
srom_1(350) <= 696291;
srom_1(351) <= 943336;
srom_1(352) <= 1225295;
srom_1(353) <= 1540844;
srom_1(354) <= 1888505;
srom_1(355) <= 2266648;
srom_1(356) <= 2673498;
srom_1(357) <= 3107148;
srom_1(358) <= 3565565;
srom_1(359) <= 4046599;
srom_1(360) <= 4547994;
srom_1(361) <= 5067399;
srom_1(362) <= 5602378;
srom_1(363) <= 6150423;
srom_1(364) <= 6708963;
srom_1(365) <= 7275380;
srom_1(366) <= 7847017;
srom_1(367) <= 8421194;
srom_1(368) <= 8995218;
srom_1(369) <= 9566398;
srom_1(370) <= 10132054;
srom_1(371) <= 10689535;
srom_1(372) <= 11236226;
srom_1(373) <= 11769563;
srom_1(374) <= 12287046;
srom_1(375) <= 12786248;
srom_1(376) <= 13264828;
srom_1(377) <= 13720541;
srom_1(378) <= 14151251;
srom_1(379) <= 14554939;
srom_1(380) <= 14929710;
srom_1(381) <= 15273807;
srom_1(382) <= 15585618;
srom_1(383) <= 15863679;
srom_1(384) <= 16106688;
srom_1(385) <= 16313503;
srom_1(386) <= 16483156;
srom_1(387) <= 16614851;
srom_1(388) <= 16707970;
srom_1(389) <= 16762076;
srom_1(390) <= 16776917;
srom_1(391) <= 16752422;
srom_1(392) <= 16688706;
srom_1(393) <= 16586068;
srom_1(394) <= 16444990;
srom_1(395) <= 16266132;
srom_1(396) <= 16050334;
srom_1(397) <= 15798607;
srom_1(398) <= 15512132;
srom_1(399) <= 15192253;
srom_1(400) <= 14840469;
srom_1(401) <= 14458430;
srom_1(402) <= 14047928;
srom_1(403) <= 13610887;
srom_1(404) <= 13149357;
srom_1(405) <= 12665502;
srom_1(406) <= 12161591;
srom_1(407) <= 11639988;
srom_1(408) <= 11103138;
srom_1(409) <= 10553558;
srom_1(410) <= 9993826;
srom_1(411) <= 9426567;
srom_1(412) <= 8854440;
srom_1(413) <= 8280129;
srom_1(414) <= 7706327;
srom_1(415) <= 7135724;
srom_1(416) <= 6570996;
srom_1(417) <= 6014791;
srom_1(418) <= 5469719;
srom_1(419) <= 4938334;
srom_1(420) <= 4423128;
srom_1(421) <= 3926518;
srom_1(422) <= 3450832;
srom_1(423) <= 2998301;
srom_1(424) <= 2571047;
srom_1(425) <= 2171074;
srom_1(426) <= 1800257;
srom_1(427) <= 1460335;
srom_1(428) <= 1152902;
srom_1(429) <= 879399;
srom_1(430) <= 641110;
srom_1(431) <= 439151;
srom_1(432) <= 274471;
srom_1(433) <= 147840;
srom_1(434) <= 59853;
srom_1(435) <= 10922;
srom_1(436) <= 1277;
srom_1(437) <= 30964;
srom_1(438) <= 99842;
srom_1(439) <= 207589;
srom_1(440) <= 353699;
srom_1(441) <= 537489;
srom_1(442) <= 758094;
srom_1(443) <= 1014482;
srom_1(444) <= 1305449;
srom_1(445) <= 1629632;
srom_1(446) <= 1985510;
srom_1(447) <= 2371415;
srom_1(448) <= 2785536;
srom_1(449) <= 3225932;
srom_1(450) <= 3690537;
srom_1(451) <= 4177173;
srom_1(452) <= 4683558;
srom_1(453) <= 5207317;
srom_1(454) <= 5745995;
srom_1(455) <= 6297064;
srom_1(456) <= 6857942;
srom_1(457) <= 7425997;
srom_1(458) <= 7998567;
srom_1(459) <= 8572965;
srom_1(460) <= 9146499;
srom_1(461) <= 9716479;
srom_1(462) <= 10280232;
srom_1(463) <= 10835114;
srom_1(464) <= 11378524;
srom_1(465) <= 11907913;
srom_1(466) <= 12420799;
srom_1(467) <= 12914777;
srom_1(468) <= 13387530;
srom_1(469) <= 13836841;
srom_1(470) <= 14260604;
srom_1(471) <= 14656830;
srom_1(472) <= 15023663;
srom_1(473) <= 15359382;
srom_1(474) <= 15662413;
srom_1(475) <= 15931334;
srom_1(476) <= 16164884;
srom_1(477) <= 16361970;
srom_1(478) <= 16521665;
srom_1(479) <= 16643221;
srom_1(480) <= 16726069;
srom_1(481) <= 16769819;
srom_1(482) <= 16774268;
srom_1(483) <= 16739393;
srom_1(484) <= 16665358;
srom_1(485) <= 16552510;
srom_1(486) <= 16401380;
srom_1(487) <= 16212674;
srom_1(488) <= 15987279;
srom_1(489) <= 15726252;
srom_1(490) <= 15430815;
srom_1(491) <= 15102355;
srom_1(492) <= 14742412;
srom_1(493) <= 14352674;
srom_1(494) <= 13934968;
srom_1(495) <= 13491254;
srom_1(496) <= 13023611;
srom_1(497) <= 12534233;
srom_1(498) <= 12025415;
srom_1(499) <= 11499543;
srom_1(500) <= 10959082;
srom_1(501) <= 10406568;
srom_1(502) <= 9844591;
srom_1(503) <= 9275786;
srom_1(504) <= 8702821;
srom_1(505) <= 8128382;
srom_1(506) <= 7555164;
srom_1(507) <= 6985854;
srom_1(508) <= 6423122;
srom_1(509) <= 5869607;
srom_1(510) <= 5327904;
srom_1(511) <= 4800554;
srom_1(512) <= 4290029;
srom_1(513) <= 3798725;
srom_1(514) <= 3328943;
srom_1(515) <= 2882888;
srom_1(516) <= 2462652;
srom_1(517) <= 2070204;
srom_1(518) <= 1707386;
srom_1(519) <= 1375898;
srom_1(520) <= 1077294;
srom_1(521) <= 812977;
srom_1(522) <= 584184;
srom_1(523) <= 391988;
srom_1(524) <= 237292;
srom_1(525) <= 120819;
srom_1(526) <= 43118;
srom_1(527) <= 4551;
srom_1(528) <= 5300;
srom_1(529) <= 45361;
srom_1(530) <= 124546;
srom_1(531) <= 242484;
srom_1(532) <= 398623;
srom_1(533) <= 592229;
srom_1(534) <= 822395;
srom_1(535) <= 1088042;
srom_1(536) <= 1387923;
srom_1(537) <= 1720633;
srom_1(538) <= 2084612;
srom_1(539) <= 2478152;
srom_1(540) <= 2899408;
srom_1(541) <= 3346405;
srom_1(542) <= 3817047;
srom_1(543) <= 4309126;
srom_1(544) <= 4820335;
srom_1(545) <= 5348277;
srom_1(546) <= 5890477;
srom_1(547) <= 6444390;
srom_1(548) <= 7007421;
srom_1(549) <= 7576929;
srom_1(550) <= 8150243;
srom_1(551) <= 8724675;
srom_1(552) <= 9297531;
srom_1(553) <= 9866125;
srom_1(554) <= 10427790;
srom_1(555) <= 10979892;
srom_1(556) <= 11519844;
srom_1(557) <= 12045111;
srom_1(558) <= 12553232;
srom_1(559) <= 13041824;
srom_1(560) <= 13508595;
srom_1(561) <= 13951357;
srom_1(562) <= 14368033;
srom_1(563) <= 14756670;
srom_1(564) <= 15115445;
srom_1(565) <= 15442675;
srom_1(566) <= 15736826;
srom_1(567) <= 15996519;
srom_1(568) <= 16220536;
srom_1(569) <= 16407826;
srom_1(570) <= 16557511;
srom_1(571) <= 16668889;
srom_1(572) <= 16741439;
srom_1(573) <= 16774819;
srom_1(574) <= 16768873;
srom_1(575) <= 16723629;
srom_1(576) <= 16639300;
srom_1(577) <= 16516280;
srom_1(578) <= 16355147;
srom_1(579) <= 16156655;
srom_1(580) <= 15921737;
srom_1(581) <= 15651494;
srom_1(582) <= 15347192;
srom_1(583) <= 15010259;
srom_1(584) <= 14642275;
srom_1(585) <= 14244965;
srom_1(586) <= 13820193;
srom_1(587) <= 13369950;
srom_1(588) <= 12896348;
srom_1(589) <= 12401607;
srom_1(590) <= 11888048;
srom_1(591) <= 11358080;
srom_1(592) <= 10814186;
srom_1(593) <= 10258918;
srom_1(594) <= 9694879;
srom_1(595) <= 9124715;
srom_1(596) <= 8551099;
srom_1(597) <= 7976721;
srom_1(598) <= 7404274;
srom_1(599) <= 6836444;
srom_1(600) <= 6275891;
srom_1(601) <= 5725247;
srom_1(602) <= 5187091;
srom_1(603) <= 4663949;
srom_1(604) <= 4158273;
srom_1(605) <= 3672434;
srom_1(606) <= 3208711;
srom_1(607) <= 2769278;
srom_1(608) <= 2356197;
srom_1(609) <= 1971403;
srom_1(610) <= 1616702;
srom_1(611) <= 1293756;
srom_1(612) <= 1004081;
srom_1(613) <= 749034;
srom_1(614) <= 529812;
srom_1(615) <= 347443;
srom_1(616) <= 202781;
srom_1(617) <= 96506;
srom_1(618) <= 29115;
srom_1(619) <= 924;
srom_1(620) <= 12066;
srom_1(621) <= 62489;
srom_1(622) <= 151956;
srom_1(623) <= 280047;
srom_1(624) <= 446162;
srom_1(625) <= 649522;
srom_1(626) <= 889173;
srom_1(627) <= 1163992;
srom_1(628) <= 1472689;
srom_1(629) <= 1813817;
srom_1(630) <= 2185777;
srom_1(631) <= 2586824;
srom_1(632) <= 3015077;
srom_1(633) <= 3468529;
srom_1(634) <= 3945053;
srom_1(635) <= 4442414;
srom_1(636) <= 4958280;
srom_1(637) <= 5490233;
srom_1(638) <= 6035776;
srom_1(639) <= 6592353;
srom_1(640) <= 7157353;
srom_1(641) <= 7728127;
srom_1(642) <= 8301998;
srom_1(643) <= 8876276;
srom_1(644) <= 9448266;
srom_1(645) <= 10015287;
srom_1(646) <= 10574680;
srom_1(647) <= 11123822;
srom_1(648) <= 11660138;
srom_1(649) <= 12181112;
srom_1(650) <= 12684302;
srom_1(651) <= 13167348;
srom_1(652) <= 13627985;
srom_1(653) <= 14064052;
srom_1(654) <= 14473506;
srom_1(655) <= 14854425;
srom_1(656) <= 15205024;
srom_1(657) <= 15523658;
srom_1(658) <= 15808833;
srom_1(659) <= 16059213;
srom_1(660) <= 16273622;
srom_1(661) <= 16451056;
srom_1(662) <= 16590683;
srom_1(663) <= 16691847;
srom_1(664) <= 16754074;
srom_1(665) <= 16777072;
srom_1(666) <= 16760735;
srom_1(667) <= 16705137;
srom_1(668) <= 16610540;
srom_1(669) <= 16477388;
srom_1(670) <= 16306305;
srom_1(671) <= 16098093;
srom_1(672) <= 15853729;
srom_1(673) <= 15574358;
srom_1(674) <= 15261290;
srom_1(675) <= 14915995;
srom_1(676) <= 14540090;
srom_1(677) <= 14135338;
srom_1(678) <= 13703639;
srom_1(679) <= 13247015;
srom_1(680) <= 12767608;
srom_1(681) <= 12267667;
srom_1(682) <= 11749536;
srom_1(683) <= 11215644;
srom_1(684) <= 10668495;
srom_1(685) <= 10110655;
srom_1(686) <= 9544740;
srom_1(687) <= 8973403;
srom_1(688) <= 8399324;
srom_1(689) <= 7825194;
srom_1(690) <= 7253707;
srom_1(691) <= 6687541;
srom_1(692) <= 6129353;
srom_1(693) <= 5581759;
srom_1(694) <= 5047327;
srom_1(695) <= 4528563;
srom_1(696) <= 4027901;
srom_1(697) <= 3547687;
srom_1(698) <= 3090174;
srom_1(699) <= 2657508;
srom_1(700) <= 2251716;
srom_1(701) <= 1874703;
srom_1(702) <= 1528235;
srom_1(703) <= 1213938;
srom_1(704) <= 933285;
srom_1(705) <= 687593;
srom_1(706) <= 478014;
srom_1(707) <= 305530;
srom_1(708) <= 170951;
srom_1(709) <= 74907;
srom_1(710) <= 17849;
srom_1(711) <= 44;
srom_1(712) <= 21576;
srom_1(713) <= 82343;
srom_1(714) <= 182062;
srom_1(715) <= 320264;
srom_1(716) <= 496302;
srom_1(717) <= 709349;
srom_1(718) <= 958406;
srom_1(719) <= 1242307;
srom_1(720) <= 1559719;
srom_1(721) <= 1909154;
srom_1(722) <= 2288973;
srom_1(723) <= 2697396;
srom_1(724) <= 3132506;
srom_1(725) <= 3592264;
srom_1(726) <= 4074514;
srom_1(727) <= 4576995;
srom_1(728) <= 5097349;
srom_1(729) <= 5633137;
srom_1(730) <= 6181846;
srom_1(731) <= 6740904;
srom_1(732) <= 7307688;
srom_1(733) <= 7879541;
srom_1(734) <= 8453782;
srom_1(735) <= 9027716;
srom_1(736) <= 9598654;
srom_1(737) <= 10163917;
srom_1(738) <= 10720855;
srom_1(739) <= 11266857;
srom_1(740) <= 11799361;
srom_1(741) <= 12315872;
srom_1(742) <= 12813965;
srom_1(743) <= 13291307;
srom_1(744) <= 13745659;
srom_1(745) <= 14174889;
srom_1(746) <= 14576986;
srom_1(747) <= 14950063;
srom_1(748) <= 15292371;
srom_1(749) <= 15602305;
srom_1(750) <= 15878412;
srom_1(751) <= 16119396;
srom_1(752) <= 16324128;
srom_1(753) <= 16491647;
srom_1(754) <= 16621169;
srom_1(755) <= 16712085;
srom_1(756) <= 16763970;
srom_1(757) <= 16776580;
srom_1(758) <= 16749855;
srom_1(759) <= 16683922;
srom_1(760) <= 16579089;
srom_1(761) <= 16435849;
srom_1(762) <= 16254872;
srom_1(763) <= 16037007;
srom_1(764) <= 15783276;
srom_1(765) <= 15494870;
srom_1(766) <= 15173139;
srom_1(767) <= 14819594;
srom_1(768) <= 14435891;
srom_1(769) <= 14023831;
srom_1(770) <= 13585345;
srom_1(771) <= 13122490;
srom_1(772) <= 12637436;
srom_1(773) <= 12132457;
srom_1(774) <= 11609923;
srom_1(775) <= 11072283;
srom_1(776) <= 10522058;
srom_1(777) <= 9961828;
srom_1(778) <= 9394222;
srom_1(779) <= 8821899;
srom_1(780) <= 8247545;
srom_1(781) <= 7673852;
srom_1(782) <= 7103511;
srom_1(783) <= 6539196;
srom_1(784) <= 5983554;
srom_1(785) <= 5439189;
srom_1(786) <= 4908656;
srom_1(787) <= 4394441;
srom_1(788) <= 3898957;
srom_1(789) <= 3424525;
srom_1(790) <= 2973372;
srom_1(791) <= 2547613;
srom_1(792) <= 2149245;
srom_1(793) <= 1780135;
srom_1(794) <= 1442014;
srom_1(795) <= 1136468;
srom_1(796) <= 864930;
srom_1(797) <= 628674;
srom_1(798) <= 428806;
srom_1(799) <= 266264;
srom_1(800) <= 141811;
srom_1(801) <= 56030;
srom_1(802) <= 9323;
srom_1(803) <= 1910;
srom_1(804) <= 33824;
srom_1(805) <= 104917;
srom_1(806) <= 214855;
srom_1(807) <= 363123;
srom_1(808) <= 549025;
srom_1(809) <= 771689;
srom_1(810) <= 1030072;
srom_1(811) <= 1322962;
srom_1(812) <= 1648984;
srom_1(813) <= 2006611;
srom_1(814) <= 2394166;
srom_1(815) <= 2809830;
srom_1(816) <= 3251656;
srom_1(817) <= 3717570;
srom_1(818) <= 4205388;
srom_1(819) <= 4712823;
srom_1(820) <= 5237495;
srom_1(821) <= 5776943;
srom_1(822) <= 6328639;
srom_1(823) <= 6889994;
srom_1(824) <= 7458377;
srom_1(825) <= 8031122;
srom_1(826) <= 8605543;
srom_1(827) <= 9178948;
srom_1(828) <= 9748645;
srom_1(829) <= 10311966;
srom_1(830) <= 10866267;
srom_1(831) <= 11408949;
srom_1(832) <= 11937468;
srom_1(833) <= 12449345;
srom_1(834) <= 12942180;
srom_1(835) <= 13413662;
srom_1(836) <= 13861579;
srom_1(837) <= 14283832;
srom_1(838) <= 14678440;
srom_1(839) <= 15043553;
srom_1(840) <= 15377458;
srom_1(841) <= 15678591;
srom_1(842) <= 15945538;
srom_1(843) <= 16177048;
srom_1(844) <= 16372035;
srom_1(845) <= 16529586;
srom_1(846) <= 16648960;
srom_1(847) <= 16729599;
srom_1(848) <= 16771124;
srom_1(849) <= 16773341;
srom_1(850) <= 16736239;
srom_1(851) <= 16659991;
srom_1(852) <= 16544957;
srom_1(853) <= 16391674;
srom_1(854) <= 16200863;
srom_1(855) <= 15973417;
srom_1(856) <= 15710403;
srom_1(857) <= 15413055;
srom_1(858) <= 15082767;
srom_1(859) <= 14721087;
srom_1(860) <= 14329712;
srom_1(861) <= 13910478;
srom_1(862) <= 13465349;
srom_1(863) <= 12996414;
srom_1(864) <= 12505872;
srom_1(865) <= 11996022;
srom_1(866) <= 11469256;
srom_1(867) <= 10928043;
srom_1(868) <= 10374922;
srom_1(869) <= 9812487;
srom_1(870) <= 9243374;
srom_1(871) <= 8670254;
srom_1(872) <= 8095812;
srom_1(873) <= 7522744;
srom_1(874) <= 6953736;
srom_1(875) <= 6391456;
srom_1(876) <= 5838542;
srom_1(877) <= 5297586;
srom_1(878) <= 4771125;
srom_1(879) <= 4261627;
srom_1(880) <= 3771482;
srom_1(881) <= 3302989;
srom_1(882) <= 2858344;
srom_1(883) <= 2439632;
srom_1(884) <= 2048816;
srom_1(885) <= 1687731;
srom_1(886) <= 1358068;
srom_1(887) <= 1061373;
srom_1(888) <= 799039;
srom_1(889) <= 572294;
srom_1(890) <= 382203;
srom_1(891) <= 229657;
srom_1(892) <= 115371;
srom_1(893) <= 39881;
srom_1(894) <= 3541;
srom_1(895) <= 6521;
srom_1(896) <= 48808;
srom_1(897) <= 130203;
srom_1(898) <= 250325;
srom_1(899) <= 408609;
srom_1(900) <= 604315;
srom_1(901) <= 836524;
srom_1(902) <= 1104147;
srom_1(903) <= 1405930;
srom_1(904) <= 1740457;
srom_1(905) <= 2106159;
srom_1(906) <= 2501321;
srom_1(907) <= 2924092;
srom_1(908) <= 3372487;
srom_1(909) <= 3844404;
srom_1(910) <= 4337631;
srom_1(911) <= 4849855;
srom_1(912) <= 5378672;
srom_1(913) <= 5921605;
srom_1(914) <= 6476106;
srom_1(915) <= 7039575;
srom_1(916) <= 7609370;
srom_1(917) <= 8182820;
srom_1(918) <= 8757234;
srom_1(919) <= 9329920;
srom_1(920) <= 9898192;
srom_1(921) <= 10459385;
srom_1(922) <= 11010867;
srom_1(923) <= 11550052;
srom_1(924) <= 12074413;
srom_1(925) <= 12581489;
srom_1(926) <= 13068904;
srom_1(927) <= 13534371;
srom_1(928) <= 13975707;
srom_1(929) <= 14390844;
srom_1(930) <= 14777835;
srom_1(931) <= 15134864;
srom_1(932) <= 15460257;
srom_1(933) <= 15752489;
srom_1(934) <= 16010190;
srom_1(935) <= 16232150;
srom_1(936) <= 16417329;
srom_1(937) <= 16564859;
srom_1(938) <= 16674047;
srom_1(939) <= 16744382;
srom_1(940) <= 16775534;
srom_1(941) <= 16767357;
srom_1(942) <= 16719889;
srom_1(943) <= 16633353;
srom_1(944) <= 16508154;
srom_1(945) <= 16344880;
srom_1(946) <= 16144296;
srom_1(947) <= 15907343;
srom_1(948) <= 15635132;
srom_1(949) <= 15328940;
srom_1(950) <= 14990202;
srom_1(951) <= 14620507;
srom_1(952) <= 14221589;
srom_1(953) <= 13795317;
srom_1(954) <= 13343692;
srom_1(955) <= 12868831;
srom_1(956) <= 12372960;
srom_1(957) <= 11858405;
srom_1(958) <= 11327579;
srom_1(959) <= 10782972;
srom_1(960) <= 10227136;
srom_1(961) <= 9662679;
srom_1(962) <= 9092247;
srom_1(963) <= 8518516;
srom_1(964) <= 7944175;
srom_1(965) <= 7371919;
srom_1(966) <= 6804430;
srom_1(967) <= 6244370;
srom_1(968) <= 5694365;
srom_1(969) <= 5156994;
srom_1(970) <= 4634778;
srom_1(971) <= 4130164;
srom_1(972) <= 3645520;
srom_1(973) <= 3183117;
srom_1(974) <= 2745125;
srom_1(975) <= 2333597;
srom_1(976) <= 1950463;
srom_1(977) <= 1597520;
srom_1(978) <= 1276423;
srom_1(979) <= 988677;
srom_1(980) <= 735632;
srom_1(981) <= 518474;
srom_1(982) <= 338222;
srom_1(983) <= 195721;
srom_1(984) <= 91639;
srom_1(985) <= 26465;
srom_1(986) <= 504;
srom_1(987) <= 13877;
srom_1(988) <= 66522;
srom_1(989) <= 158193;
srom_1(990) <= 288458;
srom_1(991) <= 456708;
srom_1(992) <= 662154;
srom_1(993) <= 903831;
srom_1(994) <= 1180607;
srom_1(995) <= 1491184;
srom_1(996) <= 1834105;
srom_1(997) <= 2207763;
srom_1(998) <= 2610404;
srom_1(999) <= 3040142;
srom_1(1000) <= 3494960;
srom_1(1001) <= 3972727;
srom_1(1002) <= 4471201;
srom_1(1003) <= 4988045;
srom_1(1004) <= 5520835;
srom_1(1005) <= 6067074;
srom_1(1006) <= 6624199;
srom_1(1007) <= 7189597;
srom_1(1008) <= 7760619;
srom_1(1009) <= 8334585;
srom_1(1010) <= 8908804;
srom_1(1011) <= 9480585;
srom_1(1012) <= 10047244;
srom_1(1013) <= 10606126;
srom_1(1014) <= 11154608;
srom_1(1015) <= 11690121;
srom_1(1016) <= 12210151;
srom_1(1017) <= 12712260;
srom_1(1018) <= 13194095;
srom_1(1019) <= 13653395;
srom_1(1020) <= 14088007;
srom_1(1021) <= 14495892;
srom_1(1022) <= 14875138;
srom_1(1023) <= 15223966;
srom_1(1024) <= 15540741;
srom_1(1025) <= 15823977;
srom_1(1026) <= 16072346;
srom_1(1027) <= 16284684;
srom_1(1028) <= 16459994;
srom_1(1029) <= 16597455;
srom_1(1030) <= 16696421;
srom_1(1031) <= 16756429;
srom_1(1032) <= 16777198;
srom_1(1033) <= 16758630;
srom_1(1034) <= 16700812;
srom_1(1035) <= 16604015;
srom_1(1036) <= 16468693;
srom_1(1037) <= 16295481;
srom_1(1038) <= 16085190;
srom_1(1039) <= 15838808;
srom_1(1040) <= 15557489;
srom_1(1041) <= 15242553;
srom_1(1042) <= 14895477;
srom_1(1043) <= 14517887;
srom_1(1044) <= 14111555;
srom_1(1045) <= 13678387;
srom_1(1046) <= 13220412;
srom_1(1047) <= 12739780;
srom_1(1048) <= 12238744;
srom_1(1049) <= 11719653;
srom_1(1050) <= 11184941;
srom_1(1051) <= 10637117;
srom_1(1052) <= 10078748;
srom_1(1053) <= 9512454;
srom_1(1054) <= 8940890;
srom_1(1055) <= 8366736;
srom_1(1056) <= 7792684;
srom_1(1057) <= 7221427;
srom_1(1058) <= 6655643;
srom_1(1059) <= 6097986;
srom_1(1060) <= 5551070;
srom_1(1061) <= 5017461;
srom_1(1062) <= 4499660;
srom_1(1063) <= 4000095;
srom_1(1064) <= 3521110;
srom_1(1065) <= 3064950;
srom_1(1066) <= 2633754;
srom_1(1067) <= 2229545;
srom_1(1068) <= 1854218;
srom_1(1069) <= 1509533;
srom_1(1070) <= 1197107;
srom_1(1071) <= 918403;
srom_1(1072) <= 674730;
srom_1(1073) <= 467230;
srom_1(1074) <= 296876;
srom_1(1075) <= 164467;
srom_1(1076) <= 70624;
srom_1(1077) <= 15787;
srom_1(1078) <= 213;
srom_1(1079) <= 23975;
srom_1(1080) <= 86961;
srom_1(1081) <= 188877;
srom_1(1082) <= 329244;
srom_1(1083) <= 507404;
srom_1(1084) <= 722522;
srom_1(1085) <= 973588;
srom_1(1086) <= 1259427;
srom_1(1087) <= 1578696;
srom_1(1088) <= 1929900;
srom_1(1089) <= 2311390;
srom_1(1090) <= 2721379;
srom_1(1091) <= 3157943;
srom_1(1092) <= 3619036;
srom_1(1093) <= 4102495;
srom_1(1094) <= 4606053;
srom_1(1095) <= 5127348;
srom_1(1096) <= 5663937;
srom_1(1097) <= 6213303;
srom_1(1098) <= 6772869;
srom_1(1099) <= 7340012;
srom_1(1100) <= 7912073;
srom_1(1101) <= 8486368;
srom_1(1102) <= 9060204;
srom_1(1103) <= 9630892;
srom_1(1104) <= 10195753;
srom_1(1105) <= 10752141;
srom_1(1106) <= 11297445;
srom_1(1107) <= 11829108;
srom_1(1108) <= 12344638;
srom_1(1109) <= 12841616;
srom_1(1110) <= 13317713;
srom_1(1111) <= 13770696;
srom_1(1112) <= 14198440;
srom_1(1113) <= 14598940;
srom_1(1114) <= 14970317;
srom_1(1115) <= 15310830;
srom_1(1116) <= 15618883;
srom_1(1117) <= 15893031;
srom_1(1118) <= 16131988;
srom_1(1119) <= 16334633;
srom_1(1120) <= 16500017;
srom_1(1121) <= 16627363;
srom_1(1122) <= 16716075;
srom_1(1123) <= 16765737;
srom_1(1124) <= 16776116;
srom_1(1125) <= 16747162;
srom_1(1126) <= 16679013;
srom_1(1127) <= 16571987;
srom_1(1128) <= 16426586;
srom_1(1129) <= 16243493;
srom_1(1130) <= 16023565;
srom_1(1131) <= 15767834;
srom_1(1132) <= 15477499;
srom_1(1133) <= 15153923;
srom_1(1134) <= 14798621;
srom_1(1135) <= 14413261;
srom_1(1136) <= 13999648;
srom_1(1137) <= 13559724;
srom_1(1138) <= 13095551;
srom_1(1139) <= 12609305;
srom_1(1140) <= 12103267;
srom_1(1141) <= 11579810;
srom_1(1142) <= 11041387;
srom_1(1143) <= 10490526;
srom_1(1144) <= 9929807;
srom_1(1145) <= 9361861;
srom_1(1146) <= 8789352;
srom_1(1147) <= 8214963;
srom_1(1148) <= 7641388;
srom_1(1149) <= 7071317;
srom_1(1150) <= 6507424;
srom_1(1151) <= 5952352;
srom_1(1152) <= 5408705;
srom_1(1153) <= 4879031;
srom_1(1154) <= 4365815;
srom_1(1155) <= 3871463;
srom_1(1156) <= 3398293;
srom_1(1157) <= 2948525;
srom_1(1158) <= 2524268;
srom_1(1159) <= 2127510;
srom_1(1160) <= 1760112;
srom_1(1161) <= 1423798;
srom_1(1162) <= 1120145;
srom_1(1163) <= 850575;
srom_1(1164) <= 616354;
srom_1(1165) <= 418580;
srom_1(1166) <= 258180;
srom_1(1167) <= 135906;
srom_1(1168) <= 52332;
srom_1(1169) <= 7850;
srom_1(1170) <= 2668;
srom_1(1171) <= 36811;
srom_1(1172) <= 110118;
srom_1(1173) <= 222245;
srom_1(1174) <= 372668;
srom_1(1175) <= 560680;
srom_1(1176) <= 785400;
srom_1(1177) <= 1045774;
srom_1(1178) <= 1340581;
srom_1(1179) <= 1668438;
srom_1(1180) <= 2027809;
srom_1(1181) <= 2417008;
srom_1(1182) <= 2834209;
srom_1(1183) <= 3277457;
srom_1(1184) <= 3744673;
srom_1(1185) <= 4233666;
srom_1(1186) <= 4742143;
srom_1(1187) <= 5267720;
srom_1(1188) <= 5807931;
srom_1(1189) <= 6360244;
srom_1(1190) <= 6922069;
srom_1(1191) <= 7490771;
srom_1(1192) <= 8063683;
srom_1(1193) <= 8638119;
srom_1(1194) <= 9211384;
srom_1(1195) <= 9780792;
srom_1(1196) <= 10343671;
srom_1(1197) <= 10897382;
srom_1(1198) <= 11439328;
srom_1(1199) <= 11966969;
srom_1(1200) <= 12477829;
srom_1(1201) <= 12969514;
srom_1(1202) <= 13439717;
srom_1(1203) <= 13886234;
srom_1(1204) <= 14306971;
srom_1(1205) <= 14699954;
srom_1(1206) <= 15063342;
srom_1(1207) <= 15395429;
srom_1(1208) <= 15694658;
srom_1(1209) <= 15959628;
srom_1(1210) <= 16189094;
srom_1(1211) <= 16381981;
srom_1(1212) <= 16537384;
srom_1(1213) <= 16654574;
srom_1(1214) <= 16733003;
srom_1(1215) <= 16772302;
srom_1(1216) <= 16772287;
srom_1(1217) <= 16732959;
srom_1(1218) <= 16654500;
srom_1(1219) <= 16537280;
srom_1(1220) <= 16381848;
srom_1(1221) <= 16188933;
srom_1(1222) <= 15959440;
srom_1(1223) <= 15694444;
srom_1(1224) <= 15395189;
srom_1(1225) <= 15063077;
srom_1(1226) <= 14699667;
srom_1(1227) <= 14306661;
srom_1(1228) <= 13885904;
srom_1(1229) <= 13439369;
srom_1(1230) <= 12969148;
srom_1(1231) <= 12477448;
srom_1(1232) <= 11966574;
srom_1(1233) <= 11438922;
srom_1(1234) <= 10896965;
srom_1(1235) <= 10343246;
srom_1(1236) <= 9780361;
srom_1(1237) <= 9210950;
srom_1(1238) <= 8637682;
srom_1(1239) <= 8063246;
srom_1(1240) <= 7490337;
srom_1(1241) <= 6921639;
srom_1(1242) <= 6359820;
srom_1(1243) <= 5807516;
srom_1(1244) <= 5267314;
srom_1(1245) <= 4741750;
srom_1(1246) <= 4233287;
srom_1(1247) <= 3744310;
srom_1(1248) <= 3277111;
srom_1(1249) <= 2833882;
srom_1(1250) <= 2416701;
srom_1(1251) <= 2027524;
srom_1(1252) <= 1668177;
srom_1(1253) <= 1340344;
srom_1(1254) <= 1045562;
srom_1(1255) <= 785215;
srom_1(1256) <= 560523;
srom_1(1257) <= 372539;
srom_1(1258) <= 222145;
srom_1(1259) <= 110047;
srom_1(1260) <= 36770;
srom_1(1261) <= 2657;
srom_1(1262) <= 7869;
srom_1(1263) <= 52381;
srom_1(1264) <= 135985;
srom_1(1265) <= 258288;
srom_1(1266) <= 418716;
srom_1(1267) <= 616519;
srom_1(1268) <= 850767;
srom_1(1269) <= 1120363;
srom_1(1270) <= 1424042;
srom_1(1271) <= 1760380;
srom_1(1272) <= 2127800;
srom_1(1273) <= 2524580;
srom_1(1274) <= 2948858;
srom_1(1275) <= 3398645;
srom_1(1276) <= 3871831;
srom_1(1277) <= 4366198;
srom_1(1278) <= 4879427;
srom_1(1279) <= 5409113;
srom_1(1280) <= 5952770;
srom_1(1281) <= 6507850;
srom_1(1282) <= 7071749;
srom_1(1283) <= 7641823;
srom_1(1284) <= 8215399;
srom_1(1285) <= 8789788;
srom_1(1286) <= 9362295;
srom_1(1287) <= 9930236;
srom_1(1288) <= 10490948;
srom_1(1289) <= 11041802;
srom_1(1290) <= 11580213;
srom_1(1291) <= 12103658;
srom_1(1292) <= 12609682;
srom_1(1293) <= 13095912;
srom_1(1294) <= 13560068;
srom_1(1295) <= 13999973;
srom_1(1296) <= 14413564;
srom_1(1297) <= 14798903;
srom_1(1298) <= 15154181;
srom_1(1299) <= 15477733;
srom_1(1300) <= 15768042;
srom_1(1301) <= 16023746;
srom_1(1302) <= 16243646;
srom_1(1303) <= 16426711;
srom_1(1304) <= 16572083;
srom_1(1305) <= 16679080;
srom_1(1306) <= 16747199;
srom_1(1307) <= 16776123;
srom_1(1308) <= 16765714;
srom_1(1309) <= 16716023;
srom_1(1310) <= 16627281;
srom_1(1311) <= 16499905;
srom_1(1312) <= 16334493;
srom_1(1313) <= 16131820;
srom_1(1314) <= 15892836;
srom_1(1315) <= 15618662;
srom_1(1316) <= 15310584;
srom_1(1317) <= 14970046;
srom_1(1318) <= 14598646;
srom_1(1319) <= 14198125;
srom_1(1320) <= 13770361;
srom_1(1321) <= 13317360;
srom_1(1322) <= 12841246;
srom_1(1323) <= 12344253;
srom_1(1324) <= 11828710;
srom_1(1325) <= 11297035;
srom_1(1326) <= 10751722;
srom_1(1327) <= 10195327;
srom_1(1328) <= 9630460;
srom_1(1329) <= 9059769;
srom_1(1330) <= 8485931;
srom_1(1331) <= 7911637;
srom_1(1332) <= 7339579;
srom_1(1333) <= 6772441;
srom_1(1334) <= 6212881;
srom_1(1335) <= 5663524;
srom_1(1336) <= 5126946;
srom_1(1337) <= 4605663;
srom_1(1338) <= 4102120;
srom_1(1339) <= 3618677;
srom_1(1340) <= 3157602;
srom_1(1341) <= 2721057;
srom_1(1342) <= 2311089;
srom_1(1343) <= 1929621;
srom_1(1344) <= 1578441;
srom_1(1345) <= 1259197;
srom_1(1346) <= 973384;
srom_1(1347) <= 722344;
srom_1(1348) <= 507254;
srom_1(1349) <= 329123;
srom_1(1350) <= 188785;
srom_1(1351) <= 86898;
srom_1(1352) <= 23942;
srom_1(1353) <= 210;
srom_1(1354) <= 15814;
srom_1(1355) <= 70681;
srom_1(1356) <= 164554;
srom_1(1357) <= 296992;
srom_1(1358) <= 467374;
srom_1(1359) <= 674902;
srom_1(1360) <= 918602;
srom_1(1361) <= 1197331;
srom_1(1362) <= 1509783;
srom_1(1363) <= 1854492;
srom_1(1364) <= 2229842;
srom_1(1365) <= 2634072;
srom_1(1366) <= 3065287;
srom_1(1367) <= 3521465;
srom_1(1368) <= 4000467;
srom_1(1369) <= 4500046;
srom_1(1370) <= 5017861;
srom_1(1371) <= 5551481;
srom_1(1372) <= 6098406;
srom_1(1373) <= 6656071;
srom_1(1374) <= 7221860;
srom_1(1375) <= 7793120;
srom_1(1376) <= 8367172;
srom_1(1377) <= 8941326;
srom_1(1378) <= 9512887;
srom_1(1379) <= 10079176;
srom_1(1380) <= 10637537;
srom_1(1381) <= 11185353;
srom_1(1382) <= 11720053;
srom_1(1383) <= 12239132;
srom_1(1384) <= 12740153;
srom_1(1385) <= 13220769;
srom_1(1386) <= 13678726;
srom_1(1387) <= 14111875;
srom_1(1388) <= 14518185;
srom_1(1389) <= 14895752;
srom_1(1390) <= 15242805;
srom_1(1391) <= 15557716;
srom_1(1392) <= 15839009;
srom_1(1393) <= 16085364;
srom_1(1394) <= 16295626;
srom_1(1395) <= 16468810;
srom_1(1396) <= 16604103;
srom_1(1397) <= 16700870;
srom_1(1398) <= 16758659;
srom_1(1399) <= 16777197;
srom_1(1400) <= 16756399;
srom_1(1401) <= 16696361;
srom_1(1402) <= 16597365;
srom_1(1403) <= 16459875;
srom_1(1404) <= 16284537;
srom_1(1405) <= 16072171;
srom_1(1406) <= 15823775;
srom_1(1407) <= 15540513;
srom_1(1408) <= 15223713;
srom_1(1409) <= 14874861;
srom_1(1410) <= 14495592;
srom_1(1411) <= 14087686;
srom_1(1412) <= 13653055;
srom_1(1413) <= 13193737;
srom_1(1414) <= 12711886;
srom_1(1415) <= 12209762;
srom_1(1416) <= 11689719;
srom_1(1417) <= 11154196;
srom_1(1418) <= 10605705;
srom_1(1419) <= 10046816;
srom_1(1420) <= 9480152;
srom_1(1421) <= 8908369;
srom_1(1422) <= 8334148;
srom_1(1423) <= 7760183;
srom_1(1424) <= 7189165;
srom_1(1425) <= 6623772;
srom_1(1426) <= 6066654;
srom_1(1427) <= 5520425;
srom_1(1428) <= 4987646;
srom_1(1429) <= 4470815;
srom_1(1430) <= 3972356;
srom_1(1431) <= 3494606;
srom_1(1432) <= 3039806;
srom_1(1433) <= 2610088;
srom_1(1434) <= 2207468;
srom_1(1435) <= 1833833;
srom_1(1436) <= 1490935;
srom_1(1437) <= 1180384;
srom_1(1438) <= 903634;
srom_1(1439) <= 661984;
srom_1(1440) <= 456566;
srom_1(1441) <= 288345;
srom_1(1442) <= 158108;
srom_1(1443) <= 66467;
srom_1(1444) <= 13852;
srom_1(1445) <= 508;
srom_1(1446) <= 26500;
srom_1(1447) <= 91704;
srom_1(1448) <= 195815;
srom_1(1449) <= 338345;
srom_1(1450) <= 518625;
srom_1(1451) <= 735811;
srom_1(1452) <= 988883;
srom_1(1453) <= 1276654;
srom_1(1454) <= 1597777;
srom_1(1455) <= 1950743;
srom_1(1456) <= 2333899;
srom_1(1457) <= 2745448;
srom_1(1458) <= 3183460;
srom_1(1459) <= 3645880;
srom_1(1460) <= 4130540;
srom_1(1461) <= 4635168;
srom_1(1462) <= 5157397;
srom_1(1463) <= 5694779;
srom_1(1464) <= 6244792;
srom_1(1465) <= 6804859;
srom_1(1466) <= 7372352;
srom_1(1467) <= 7944611;
srom_1(1468) <= 8518953;
srom_1(1469) <= 9092682;
srom_1(1470) <= 9663111;
srom_1(1471) <= 10227562;
srom_1(1472) <= 10783390;
srom_1(1473) <= 11327988;
srom_1(1474) <= 11858803;
srom_1(1475) <= 12373344;
srom_1(1476) <= 12869200;
srom_1(1477) <= 13344044;
srom_1(1478) <= 13795651;
srom_1(1479) <= 14221903;
srom_1(1480) <= 14620800;
srom_1(1481) <= 14990472;
srom_1(1482) <= 15329185;
srom_1(1483) <= 15635352;
srom_1(1484) <= 15907537;
srom_1(1485) <= 16144462;
srom_1(1486) <= 16345018;
srom_1(1487) <= 16508264;
srom_1(1488) <= 16633433;
srom_1(1489) <= 16719940;
srom_1(1490) <= 16767378;
srom_1(1491) <= 16775525;
srom_1(1492) <= 16744343;
srom_1(1493) <= 16673979;
srom_1(1494) <= 16564761;
srom_1(1495) <= 16417202;
srom_1(1496) <= 16231995;
srom_1(1497) <= 16010007;
srom_1(1498) <= 15752280;
srom_1(1499) <= 15460022;
srom_1(1500) <= 15134604;
srom_1(1501) <= 14777552;
srom_1(1502) <= 14390539;
srom_1(1503) <= 13975382;
srom_1(1504) <= 13534026;
srom_1(1505) <= 13068541;
srom_1(1506) <= 12581111;
srom_1(1507) <= 12074020;
srom_1(1508) <= 11549648;
srom_1(1509) <= 11010452;
srom_1(1510) <= 10458961;
srom_1(1511) <= 9897762;
srom_1(1512) <= 9329486;
srom_1(1513) <= 8756798;
srom_1(1514) <= 8182383;
srom_1(1515) <= 7608936;
srom_1(1516) <= 7039144;
srom_1(1517) <= 6475680;
srom_1(1518) <= 5921187;
srom_1(1519) <= 5378265;
srom_1(1520) <= 4849459;
srom_1(1521) <= 4337249;
srom_1(1522) <= 3844037;
srom_1(1523) <= 3372137;
srom_1(1524) <= 2923760;
srom_1(1525) <= 2501010;
srom_1(1526) <= 2105869;
srom_1(1527) <= 1740190;
srom_1(1528) <= 1405688;
srom_1(1529) <= 1103931;
srom_1(1530) <= 836334;
srom_1(1531) <= 604152;
srom_1(1532) <= 408475;
srom_1(1533) <= 250219;
srom_1(1534) <= 130126;
srom_1(1535) <= 48761;
srom_1(1536) <= 6504;
srom_1(1537) <= 3553;
srom_1(1538) <= 39923;
srom_1(1539) <= 115443;
srom_1(1540) <= 229758;
srom_1(1541) <= 382334;
srom_1(1542) <= 572453;
srom_1(1543) <= 799225;
srom_1(1544) <= 1061586;
srom_1(1545) <= 1358306;
srom_1(1546) <= 1687993;
srom_1(1547) <= 2049102;
srom_1(1548) <= 2439939;
srom_1(1549) <= 2858672;
srom_1(1550) <= 3303336;
srom_1(1551) <= 3771847;
srom_1(1552) <= 4262007;
srom_1(1553) <= 4771519;
srom_1(1554) <= 5297992;
srom_1(1555) <= 5838958;
srom_1(1556) <= 6391880;
srom_1(1557) <= 6954166;
srom_1(1558) <= 7523178;
srom_1(1559) <= 8096249;
srom_1(1560) <= 8670690;
srom_1(1561) <= 9243809;
srom_1(1562) <= 9812917;
srom_1(1563) <= 10375346;
srom_1(1564) <= 10928459;
srom_1(1565) <= 11469662;
srom_1(1566) <= 11996416;
srom_1(1567) <= 12506252;
srom_1(1568) <= 12996779;
srom_1(1569) <= 13465697;
srom_1(1570) <= 13910807;
srom_1(1571) <= 14330021;
srom_1(1572) <= 14721373;
srom_1(1573) <= 15083030;
srom_1(1574) <= 15413293;
srom_1(1575) <= 15710616;
srom_1(1576) <= 15973603;
srom_1(1577) <= 16201022;
srom_1(1578) <= 16391805;
srom_1(1579) <= 16545059;
srom_1(1580) <= 16660064;
srom_1(1581) <= 16736282;
srom_1(1582) <= 16773354;
srom_1(1583) <= 16771108;
srom_1(1584) <= 16729553;
srom_1(1585) <= 16648884;
srom_1(1586) <= 16529480;
srom_1(1587) <= 16371901;
srom_1(1588) <= 16176886;
srom_1(1589) <= 15945348;
srom_1(1590) <= 15678375;
srom_1(1591) <= 15377217;
srom_1(1592) <= 15043287;
srom_1(1593) <= 14678151;
srom_1(1594) <= 14283521;
srom_1(1595) <= 13861248;
srom_1(1596) <= 13413312;
srom_1(1597) <= 12941813;
srom_1(1598) <= 12448963;
srom_1(1599) <= 11937072;
srom_1(1600) <= 11408542;
srom_1(1601) <= 10865849;
srom_1(1602) <= 10311541;
srom_1(1603) <= 9748215;
srom_1(1604) <= 9178513;
srom_1(1605) <= 8605107;
srom_1(1606) <= 8030686;
srom_1(1607) <= 7457943;
srom_1(1608) <= 6889564;
srom_1(1609) <= 6328215;
srom_1(1610) <= 5776528;
srom_1(1611) <= 5237090;
srom_1(1612) <= 4712430;
srom_1(1613) <= 4205010;
srom_1(1614) <= 3717207;
srom_1(1615) <= 3251310;
srom_1(1616) <= 2809504;
srom_1(1617) <= 2393860;
srom_1(1618) <= 2006328;
srom_1(1619) <= 1648724;
srom_1(1620) <= 1322726;
srom_1(1621) <= 1029863;
srom_1(1622) <= 771507;
srom_1(1623) <= 548870;
srom_1(1624) <= 362996;
srom_1(1625) <= 214757;
srom_1(1626) <= 104848;
srom_1(1627) <= 33785;
srom_1(1628) <= 1900;
srom_1(1629) <= 9344;
srom_1(1630) <= 56080;
srom_1(1631) <= 141891;
srom_1(1632) <= 266373;
srom_1(1633) <= 428944;
srom_1(1634) <= 628839;
srom_1(1635) <= 865124;
srom_1(1636) <= 1136688;
srom_1(1637) <= 1442259;
srom_1(1638) <= 1780404;
srom_1(1639) <= 2149537;
srom_1(1640) <= 2547927;
srom_1(1641) <= 2973706;
srom_1(1642) <= 3424877;
srom_1(1643) <= 3899325;
srom_1(1644) <= 4394825;
srom_1(1645) <= 4909053;
srom_1(1646) <= 5439598;
srom_1(1647) <= 5983972;
srom_1(1648) <= 6539622;
srom_1(1649) <= 7103942;
srom_1(1650) <= 7674287;
srom_1(1651) <= 8247981;
srom_1(1652) <= 8822335;
srom_1(1653) <= 9394655;
srom_1(1654) <= 9962257;
srom_1(1655) <= 10522480;
srom_1(1656) <= 11072696;
srom_1(1657) <= 11610326;
srom_1(1658) <= 12132848;
srom_1(1659) <= 12637812;
srom_1(1660) <= 13122850;
srom_1(1661) <= 13585688;
srom_1(1662) <= 14024154;
srom_1(1663) <= 14436194;
srom_1(1664) <= 14819874;
srom_1(1665) <= 15173396;
srom_1(1666) <= 15495102;
srom_1(1667) <= 15783483;
srom_1(1668) <= 16037186;
srom_1(1669) <= 16255023;
srom_1(1670) <= 16435972;
srom_1(1671) <= 16579184;
srom_1(1672) <= 16683987;
srom_1(1673) <= 16749890;
srom_1(1674) <= 16776585;
srom_1(1675) <= 16763945;
srom_1(1676) <= 16712031;
srom_1(1677) <= 16621085;
srom_1(1678) <= 16491534;
srom_1(1679) <= 16323986;
srom_1(1680) <= 16119226;
srom_1(1681) <= 15878215;
srom_1(1682) <= 15602082;
srom_1(1683) <= 15292123;
srom_1(1684) <= 14949791;
srom_1(1685) <= 14576691;
srom_1(1686) <= 14174573;
srom_1(1687) <= 13745323;
srom_1(1688) <= 13290953;
srom_1(1689) <= 12813594;
srom_1(1690) <= 12315486;
srom_1(1691) <= 11798962;
srom_1(1692) <= 11266447;
srom_1(1693) <= 10720436;
srom_1(1694) <= 10163490;
srom_1(1695) <= 9598222;
srom_1(1696) <= 9027281;
srom_1(1697) <= 8453345;
srom_1(1698) <= 7879105;
srom_1(1699) <= 7307255;
srom_1(1700) <= 6740476;
srom_1(1701) <= 6181425;
srom_1(1702) <= 5632724;
srom_1(1703) <= 5096947;
srom_1(1704) <= 4576606;
srom_1(1705) <= 4074140;
srom_1(1706) <= 3591906;
srom_1(1707) <= 3132166;
srom_1(1708) <= 2697075;
srom_1(1709) <= 2288673;
srom_1(1710) <= 1908876;
srom_1(1711) <= 1559465;
srom_1(1712) <= 1242078;
srom_1(1713) <= 958204;
srom_1(1714) <= 709173;
srom_1(1715) <= 496154;
srom_1(1716) <= 320145;
srom_1(1717) <= 181972;
srom_1(1718) <= 82282;
srom_1(1719) <= 21544;
srom_1(1720) <= 42;
srom_1(1721) <= 17877;
srom_1(1722) <= 74965;
srom_1(1723) <= 171039;
srom_1(1724) <= 305647;
srom_1(1725) <= 478159;
srom_1(1726) <= 687767;
srom_1(1727) <= 933486;
srom_1(1728) <= 1214164;
srom_1(1729) <= 1528486;
srom_1(1730) <= 1874978;
srom_1(1731) <= 2252014;
srom_1(1732) <= 2657827;
srom_1(1733) <= 3090513;
srom_1(1734) <= 3548044;
srom_1(1735) <= 4028274;
srom_1(1736) <= 4528951;
srom_1(1737) <= 5047727;
srom_1(1738) <= 5582170;
srom_1(1739) <= 6129773;
srom_1(1740) <= 6687969;
srom_1(1741) <= 7254139;
srom_1(1742) <= 7825630;
srom_1(1743) <= 8399760;
srom_1(1744) <= 8973838;
srom_1(1745) <= 9545172;
srom_1(1746) <= 10111082;
srom_1(1747) <= 10668915;
srom_1(1748) <= 11216055;
srom_1(1749) <= 11749936;
srom_1(1750) <= 12268054;
srom_1(1751) <= 12767981;
srom_1(1752) <= 13247371;
srom_1(1753) <= 13703977;
srom_1(1754) <= 14135657;
srom_1(1755) <= 14540387;
srom_1(1756) <= 14916269;
srom_1(1757) <= 15261541;
srom_1(1758) <= 15574583;
srom_1(1759) <= 15853928;
srom_1(1760) <= 16098265;
srom_1(1761) <= 16306449;
srom_1(1762) <= 16477504;
srom_1(1763) <= 16610627;
srom_1(1764) <= 16705194;
srom_1(1765) <= 16760762;
srom_1(1766) <= 16777070;
srom_1(1767) <= 16754041;
srom_1(1768) <= 16691784;
srom_1(1769) <= 16590591;
srom_1(1770) <= 16450936;
srom_1(1771) <= 16273473;
srom_1(1772) <= 16059036;
srom_1(1773) <= 15808630;
srom_1(1774) <= 15523428;
srom_1(1775) <= 15204769;
srom_1(1776) <= 14854147;
srom_1(1777) <= 14473205;
srom_1(1778) <= 14063731;
srom_1(1779) <= 13627644;
srom_1(1780) <= 13166989;
srom_1(1781) <= 12683927;
srom_1(1782) <= 12180723;
srom_1(1783) <= 11659736;
srom_1(1784) <= 11123410;
srom_1(1785) <= 10574259;
srom_1(1786) <= 10014859;
srom_1(1787) <= 9447833;
srom_1(1788) <= 8875840;
srom_1(1789) <= 8301562;
srom_1(1790) <= 7727692;
srom_1(1791) <= 7156921;
srom_1(1792) <= 6591927;
srom_1(1793) <= 6035357;
srom_1(1794) <= 5489823;
srom_1(1795) <= 4957882;
srom_1(1796) <= 4442029;
srom_1(1797) <= 3944683;
srom_1(1798) <= 3468176;
srom_1(1799) <= 3014742;
srom_1(1800) <= 2586509;
srom_1(1801) <= 2185483;
srom_1(1802) <= 1813546;
srom_1(1803) <= 1472442;
srom_1(1804) <= 1163770;
srom_1(1805) <= 888977;
srom_1(1806) <= 649354;
srom_1(1807) <= 446022;
srom_1(1808) <= 279935;
srom_1(1809) <= 151873;
srom_1(1810) <= 62436;
srom_1(1811) <= 12043;
srom_1(1812) <= 931;
srom_1(1813) <= 29151;
srom_1(1814) <= 96572;
srom_1(1815) <= 202877;
srom_1(1816) <= 347567;
srom_1(1817) <= 529965;
srom_1(1818) <= 749215;
srom_1(1819) <= 1004288;
srom_1(1820) <= 1293989;
srom_1(1821) <= 1616959;
srom_1(1822) <= 1971684;
srom_1(1823) <= 2356500;
srom_1(1824) <= 2769602;
srom_1(1825) <= 3209054;
srom_1(1826) <= 3672795;
srom_1(1827) <= 4158650;
srom_1(1828) <= 4664340;
srom_1(1829) <= 5187495;
srom_1(1830) <= 5725661;
srom_1(1831) <= 6276314;
srom_1(1832) <= 6836873;
srom_1(1833) <= 7404708;
srom_1(1834) <= 7977157;
srom_1(1835) <= 8551535;
srom_1(1836) <= 9125150;
srom_1(1837) <= 9695310;
srom_1(1838) <= 10259343;
srom_1(1839) <= 10814604;
srom_1(1840) <= 11358488;
srom_1(1841) <= 11888445;
srom_1(1842) <= 12401991;
srom_1(1843) <= 12896716;
srom_1(1844) <= 13370301;
srom_1(1845) <= 13820525;
srom_1(1846) <= 14245277;
srom_1(1847) <= 14642566;
srom_1(1848) <= 15010527;
srom_1(1849) <= 15347436;
srom_1(1850) <= 15651712;
srom_1(1851) <= 15921929;
srom_1(1852) <= 16156820;
srom_1(1853) <= 16355283;
srom_1(1854) <= 16516388;
srom_1(1855) <= 16639379;
srom_1(1856) <= 16723678;
srom_1(1857) <= 16768892;
srom_1(1858) <= 16774808;
srom_1(1859) <= 16741398;
srom_1(1860) <= 16668819;
srom_1(1861) <= 16557412;
srom_1(1862) <= 16407697;
srom_1(1863) <= 16220379;
srom_1(1864) <= 15996335;
srom_1(1865) <= 15736615;
srom_1(1866) <= 15442438;
srom_1(1867) <= 15115184;
srom_1(1868) <= 14756386;
srom_1(1869) <= 14367727;
srom_1(1870) <= 13951030;
srom_1(1871) <= 13508250;
srom_1(1872) <= 13041461;
srom_1(1873) <= 12552853;
srom_1(1874) <= 12044718;
srom_1(1875) <= 11519438;
srom_1(1876) <= 10979477;
srom_1(1877) <= 10427366;
srom_1(1878) <= 9865695;
srom_1(1879) <= 9297097;
srom_1(1880) <= 8724239;
srom_1(1881) <= 8149807;
srom_1(1882) <= 7576495;
srom_1(1883) <= 7006991;
srom_1(1884) <= 6443966;
srom_1(1885) <= 5890060;
srom_1(1886) <= 5347870;
srom_1(1887) <= 4819940;
srom_1(1888) <= 4308744;
srom_1(1889) <= 3816681;
srom_1(1890) <= 3346056;
srom_1(1891) <= 2899078;
srom_1(1892) <= 2477842;
srom_1(1893) <= 2084324;
srom_1(1894) <= 1720368;
srom_1(1895) <= 1387683;
srom_1(1896) <= 1087827;
srom_1(1897) <= 822207;
srom_1(1898) <= 592068;
srom_1(1899) <= 398490;
srom_1(1900) <= 242380;
srom_1(1901) <= 124471;
srom_1(1902) <= 45315;
srom_1(1903) <= 5284;
srom_1(1904) <= 4565;
srom_1(1905) <= 43162;
srom_1(1906) <= 120893;
srom_1(1907) <= 237395;
srom_1(1908) <= 392120;
srom_1(1909) <= 584344;
srom_1(1910) <= 813164;
srom_1(1911) <= 1077509;
srom_1(1912) <= 1376137;
srom_1(1913) <= 1707650;
srom_1(1914) <= 2070491;
srom_1(1915) <= 2462961;
srom_1(1916) <= 2883218;
srom_1(1917) <= 3329292;
srom_1(1918) <= 3799090;
srom_1(1919) <= 4290410;
srom_1(1920) <= 4800949;
srom_1(1921) <= 5328310;
srom_1(1922) <= 5870023;
srom_1(1923) <= 6423546;
srom_1(1924) <= 6986284;
srom_1(1925) <= 7555598;
srom_1(1926) <= 8128819;
srom_1(1927) <= 8703257;
srom_1(1928) <= 9276220;
srom_1(1929) <= 9845021;
srom_1(1930) <= 10406992;
srom_1(1931) <= 10959498;
srom_1(1932) <= 11499949;
srom_1(1933) <= 12025809;
srom_1(1934) <= 12534613;
srom_1(1935) <= 13023975;
srom_1(1936) <= 13491600;
srom_1(1937) <= 13935296;
srom_1(1938) <= 14352981;
srom_1(1939) <= 14742697;
srom_1(1940) <= 15102617;
srom_1(1941) <= 15431052;
srom_1(1942) <= 15726463;
srom_1(1943) <= 15987464;
srom_1(1944) <= 16212832;
srom_1(1945) <= 16401509;
srom_1(1946) <= 16552611;
srom_1(1947) <= 16665429;
srom_1(1948) <= 16739434;
srom_1(1949) <= 16774279;
srom_1(1950) <= 16769801;
srom_1(1951) <= 16726021;
srom_1(1952) <= 16643143;
srom_1(1953) <= 16521558;
srom_1(1954) <= 16361834;
srom_1(1955) <= 16164721;
srom_1(1956) <= 15931143;
srom_1(1957) <= 15662195;
srom_1(1958) <= 15359139;
srom_1(1959) <= 15023396;
srom_1(1960) <= 14656540;
srom_1(1961) <= 14260292;
srom_1(1962) <= 13836509;
srom_1(1963) <= 13387179;
srom_1(1964) <= 12914409;
srom_1(1965) <= 12420416;
srom_1(1966) <= 11907517;
srom_1(1967) <= 11378116;
srom_1(1968) <= 10834696;
srom_1(1969) <= 10279806;
srom_1(1970) <= 9716047;
srom_1(1971) <= 9146064;
srom_1(1972) <= 8572528;
srom_1(1973) <= 7998130;
srom_1(1974) <= 7425563;
srom_1(1975) <= 6857513;
srom_1(1976) <= 6296641;
srom_1(1977) <= 5745580;
srom_1(1978) <= 5206913;
srom_1(1979) <= 4683166;
srom_1(1980) <= 4176795;
srom_1(1981) <= 3690175;
srom_1(1982) <= 3225587;
srom_1(1983) <= 2785211;
srom_1(1984) <= 2371110;
srom_1(1985) <= 1985228;
srom_1(1986) <= 1629374;
srom_1(1987) <= 1305215;
srom_1(1988) <= 1014274;
srom_1(1989) <= 757913;
srom_1(1990) <= 537335;
srom_1(1991) <= 353574;
srom_1(1992) <= 207492;
srom_1(1993) <= 99775;
srom_1(1994) <= 30926;
srom_1(1995) <= 1270;
srom_1(1996) <= 10945;
srom_1(1997) <= 59905;
srom_1(1998) <= 147921;
srom_1(1999) <= 274581;
srom_1(2000) <= 439291;
srom_1(2001) <= 641277;
srom_1(2002) <= 879594;
srom_1(2003) <= 1153122;
srom_1(2004) <= 1460581;
srom_1(2005) <= 1800527;
srom_1(2006) <= 2171367;
srom_1(2007) <= 2571362;
srom_1(2008) <= 2998636;
srom_1(2009) <= 3451185;
srom_1(2010) <= 3926888;
srom_1(2011) <= 4423513;
srom_1(2012) <= 4938732;
srom_1(2013) <= 5470128;
srom_1(2014) <= 6015210;
srom_1(2015) <= 6571422;
srom_1(2016) <= 7136155;
srom_1(2017) <= 7706762;
srom_1(2018) <= 8280566;
srom_1(2019) <= 8854876;
srom_1(2020) <= 9427000;
srom_1(2021) <= 9994255;
srom_1(2022) <= 10553980;
srom_1(2023) <= 11103551;
srom_1(2024) <= 11640390;
srom_1(2025) <= 12161981;
srom_1(2026) <= 12665878;
srom_1(2027) <= 13149716;
srom_1(2028) <= 13611229;
srom_1(2029) <= 14048250;
srom_1(2030) <= 14458732;
srom_1(2031) <= 14840748;
srom_1(2032) <= 15192509;
srom_1(2033) <= 15512363;
srom_1(2034) <= 15798812;
srom_1(2035) <= 16050512;
srom_1(2036) <= 16266282;
srom_1(2037) <= 16445111;
srom_1(2038) <= 16586161;
srom_1(2039) <= 16688769;
srom_1(2040) <= 16752455;
srom_1(2041) <= 16776921;
srom_1(2042) <= 16762050;
srom_1(2043) <= 16707914;
srom_1(2044) <= 16614765;
srom_1(2045) <= 16483041;
srom_1(2046) <= 16313360;
srom_1(2047) <= 16106516;
srom_1(2048) <= 15863481;
srom_1(2049) <= 15585394;
srom_1(2050) <= 15273558;
srom_1(2051) <= 14929436;
srom_1(2052) <= 14554643;
srom_1(2053) <= 14150934;
srom_1(2054) <= 13720204;
srom_1(2055) <= 13264472;
srom_1(2056) <= 12785876;
srom_1(2057) <= 12286659;
srom_1(2058) <= 11769163;
srom_1(2059) <= 11235815;
srom_1(2060) <= 10689115;
srom_1(2061) <= 10131627;
srom_1(2062) <= 9565965;
srom_1(2063) <= 8994783;
srom_1(2064) <= 8420758;
srom_1(2065) <= 7846582;
srom_1(2066) <= 7274947;
srom_1(2067) <= 6708536;
srom_1(2068) <= 6150002;
srom_1(2069) <= 5601966;
srom_1(2070) <= 5066998;
srom_1(2071) <= 4547606;
srom_1(2072) <= 4046225;
srom_1(2073) <= 3565208;
srom_1(2074) <= 3106809;
srom_1(2075) <= 2673178;
srom_1(2076) <= 2266349;
srom_1(2077) <= 1888229;
srom_1(2078) <= 1540592;
srom_1(2079) <= 1225067;
srom_1(2080) <= 943135;
srom_1(2081) <= 696117;
srom_1(2082) <= 485172;
srom_1(2083) <= 311289;
srom_1(2084) <= 175283;
srom_1(2085) <= 77792;
srom_1(2086) <= 19273;
srom_1(2087) <= 2;
srom_1(2088) <= 20067;
srom_1(2089) <= 79375;
srom_1(2090) <= 177648;
srom_1(2091) <= 314425;
srom_1(2092) <= 489064;
srom_1(2093) <= 700747;
srom_1(2094) <= 948482;
srom_1(2095) <= 1231105;
srom_1(2096) <= 1547293;
srom_1(2097) <= 1895562;
srom_1(2098) <= 2274278;
srom_1(2099) <= 2681668;
srom_1(2100) <= 3115818;
srom_1(2101) <= 3574695;
srom_1(2102) <= 4056146;
srom_1(2103) <= 4557913;
srom_1(2104) <= 5077644;
srom_1(2105) <= 5612901;
srom_1(2106) <= 6161174;
srom_1(2107) <= 6719893;
srom_1(2108) <= 7286436;
srom_1(2109) <= 7858148;
srom_1(2110) <= 8432348;
srom_1(2111) <= 9006342;
srom_1(2112) <= 9577440;
srom_1(2113) <= 10142963;
srom_1(2114) <= 10700259;
srom_1(2115) <= 11246715;
srom_1(2116) <= 11779768;
srom_1(2117) <= 12296919;
srom_1(2118) <= 12795742;
srom_1(2119) <= 13273899;
srom_1(2120) <= 13729147;
srom_1(2121) <= 14159352;
srom_1(2122) <= 14562495;
srom_1(2123) <= 14936687;
srom_1(2124) <= 15280173;
srom_1(2125) <= 15591342;
srom_1(2126) <= 15868734;
srom_1(2127) <= 16111050;
srom_1(2128) <= 16317153;
srom_1(2129) <= 16486076;
srom_1(2130) <= 16617027;
srom_1(2131) <= 16709392;
srom_1(2132) <= 16762739;
srom_1(2133) <= 16776816;
srom_1(2134) <= 16751558;
srom_1(2135) <= 16687083;
srom_1(2136) <= 16583694;
srom_1(2137) <= 16441875;
srom_1(2138) <= 16262291;
srom_1(2139) <= 16045785;
srom_1(2140) <= 15793372;
srom_1(2141) <= 15506236;
srom_1(2142) <= 15185723;
srom_1(2143) <= 14833335;
srom_1(2144) <= 14450726;
srom_1(2145) <= 14039690;
srom_1(2146) <= 13602154;
srom_1(2147) <= 13140169;
srom_1(2148) <= 12655903;
srom_1(2149) <= 12151626;
srom_1(2150) <= 11629703;
srom_1(2151) <= 11092582;
srom_1(2152) <= 10542780;
srom_1(2153) <= 9982877;
srom_1(2154) <= 9415498;
srom_1(2155) <= 8843303;
srom_1(2156) <= 8268976;
srom_1(2157) <= 7695210;
srom_1(2158) <= 7124696;
srom_1(2159) <= 6560109;
srom_1(2160) <= 6004096;
srom_1(2161) <= 5459265;
srom_1(2162) <= 4928170;
srom_1(2163) <= 4413303;
srom_1(2164) <= 3917077;
srom_1(2165) <= 3441820;
srom_1(2166) <= 2989760;
srom_1(2167) <= 2563017;
srom_1(2168) <= 2163592;
srom_1(2169) <= 1793359;
srom_1(2170) <= 1454052;
srom_1(2171) <= 1147265;
srom_1(2172) <= 874434;
srom_1(2173) <= 636840;
srom_1(2174) <= 435597;
srom_1(2175) <= 271648;
srom_1(2176) <= 145762;
srom_1(2177) <= 58530;
srom_1(2178) <= 10361;
srom_1(2179) <= 1480;
srom_1(2180) <= 31929;
srom_1(2181) <= 101565;
srom_1(2182) <= 210062;
srom_1(2183) <= 356911;
srom_1(2184) <= 541424;
srom_1(2185) <= 762734;
srom_1(2186) <= 1019805;
srom_1(2187) <= 1311431;
srom_1(2188) <= 1636244;
srom_1(2189) <= 1992722;
srom_1(2190) <= 2379191;
srom_1(2191) <= 2793841;
srom_1(2192) <= 3234727;
srom_1(2193) <= 3699781;
srom_1(2194) <= 4186823;
srom_1(2195) <= 4693568;
srom_1(2196) <= 5217641;
srom_1(2197) <= 5756583;
srom_1(2198) <= 6307868;
srom_1(2199) <= 6868910;
srom_1(2200) <= 7437078;
srom_1(2201) <= 8009709;
srom_1(2202) <= 8584116;
srom_1(2203) <= 9157606;
srom_1(2204) <= 9727491;
srom_1(2205) <= 10291096;
srom_1(2206) <= 10845781;
srom_1(2207) <= 11388943;
srom_1(2208) <= 11918035;
srom_1(2209) <= 12430576;
srom_1(2210) <= 12924164;
srom_1(2211) <= 13396482;
srom_1(2212) <= 13845317;
srom_1(2213) <= 14268564;
srom_1(2214) <= 14664237;
srom_1(2215) <= 15030482;
srom_1(2216) <= 15365581;
srom_1(2217) <= 15667962;
srom_1(2218) <= 15936208;
srom_1(2219) <= 16169061;
srom_1(2220) <= 16365428;
srom_1(2221) <= 16524390;
srom_1(2222) <= 16645199;
srom_1(2223) <= 16727291;
srom_1(2224) <= 16770280;
srom_1(2225) <= 16773965;
srom_1(2226) <= 16738327;
srom_1(2227) <= 16663535;
srom_1(2228) <= 16549939;
srom_1(2229) <= 16398072;
srom_1(2230) <= 16208645;
srom_1(2231) <= 15982548;
srom_1(2232) <= 15720840;
srom_1(2233) <= 15424748;
srom_1(2234) <= 15095662;
srom_1(2235) <= 14735124;
srom_1(2236) <= 14344825;
srom_1(2237) <= 13926595;
srom_1(2238) <= 13482396;
srom_1(2239) <= 13014310;
srom_1(2240) <= 12524533;
srom_1(2241) <= 12015361;
srom_1(2242) <= 11489182;
srom_1(2243) <= 10948463;
srom_1(2244) <= 10395740;
srom_1(2245) <= 9833605;
srom_1(2246) <= 9264694;
srom_1(2247) <= 8691675;
srom_1(2248) <= 8117234;
srom_1(2249) <= 7544066;
srom_1(2250) <= 6974858;
srom_1(2251) <= 6412280;
srom_1(2252) <= 5858970;
srom_1(2253) <= 5317522;
srom_1(2254) <= 4790475;
srom_1(2255) <= 4280301;
srom_1(2256) <= 3789393;
srom_1(2257) <= 3320051;
srom_1(2258) <= 2874478;
srom_1(2259) <= 2454763;
srom_1(2260) <= 2062873;
srom_1(2261) <= 1700647;
srom_1(2262) <= 1369783;
srom_1(2263) <= 1071833;
srom_1(2264) <= 808193;
srom_1(2265) <= 580101;
srom_1(2266) <= 388626;
srom_1(2267) <= 234665;
srom_1(2268) <= 118940;
srom_1(2269) <= 41996;
srom_1(2270) <= 4191;
srom_1(2271) <= 5703;
srom_1(2272) <= 46526;
srom_1(2273) <= 126468;
srom_1(2274) <= 245154;
srom_1(2275) <= 402027;
srom_1(2276) <= 596352;
srom_1(2277) <= 827218;
srom_1(2278) <= 1093542;
srom_1(2279) <= 1394074;
srom_1(2280) <= 1727407;
srom_1(2281) <= 2091976;
srom_1(2282) <= 2486072;
srom_1(2283) <= 2907847;
srom_1(2284) <= 3355323;
srom_1(2285) <= 3826403;
srom_1(2286) <= 4318875;
srom_1(2287) <= 4830433;
srom_1(2288) <= 5358675;
srom_1(2289) <= 5901126;
srom_1(2290) <= 6455242;
srom_1(2291) <= 7018424;
srom_1(2292) <= 7588031;
srom_1(2293) <= 8161393;
srom_1(2294) <= 8735820;
srom_1(2295) <= 9308618;
srom_1(2296) <= 9877103;
srom_1(2297) <= 10438607;
srom_1(2298) <= 10990498;
srom_1(2299) <= 11530188;
srom_1(2300) <= 12055146;
srom_1(2301) <= 12562911;
srom_1(2302) <= 13051101;
srom_1(2303) <= 13517426;
srom_1(2304) <= 13959701;
srom_1(2305) <= 14375851;
srom_1(2306) <= 14763925;
srom_1(2307) <= 15122103;
srom_1(2308) <= 15448705;
srom_1(2309) <= 15742199;
srom_1(2310) <= 16001211;
srom_1(2311) <= 16224524;
srom_1(2312) <= 16411092;
srom_1(2313) <= 16560040;
srom_1(2314) <= 16670669;
srom_1(2315) <= 16742460;
srom_1(2316) <= 16775078;
srom_1(2317) <= 16768368;
srom_1(2318) <= 16722363;
srom_1(2319) <= 16637278;
srom_1(2320) <= 16513512;
srom_1(2321) <= 16351646;
srom_1(2322) <= 16152438;
srom_1(2323) <= 15916823;
srom_1(2324) <= 15645906;
srom_1(2325) <= 15340957;
srom_1(2326) <= 15003405;
srom_1(2327) <= 14634835;
srom_1(2328) <= 14236974;
srom_1(2329) <= 13811688;
srom_1(2330) <= 13360971;
srom_1(2331) <= 12886937;
srom_1(2332) <= 12391809;
srom_1(2333) <= 11877908;
srom_1(2334) <= 11347645;
srom_1(2335) <= 10803506;
srom_1(2336) <= 10248043;
srom_1(2337) <= 9683860;
srom_1(2338) <= 9113604;
srom_1(2339) <= 8539947;
srom_1(2340) <= 7965581;
srom_1(2341) <= 7393198;
srom_1(2342) <= 6825484;
srom_1(2343) <= 6265099;
srom_1(2344) <= 5714672;
srom_1(2345) <= 5176785;
srom_1(2346) <= 4653958;
srom_1(2347) <= 4148645;
srom_1(2348) <= 3663214;
srom_1(2349) <= 3199942;
srom_1(2350) <= 2761002;
srom_1(2351) <= 2348451;
srom_1(2352) <= 1964225;
srom_1(2353) <= 1610125;
srom_1(2354) <= 1287812;
srom_1(2355) <= 998796;
srom_1(2356) <= 744434;
srom_1(2357) <= 525918;
srom_1(2358) <= 344273;
srom_1(2359) <= 200351;
srom_1(2360) <= 94826;
srom_1(2361) <= 28194;
srom_1(2362) <= 766;
srom_1(2363) <= 12672;
srom_1(2364) <= 63855;
srom_1(2365) <= 154076;
srom_1(2366) <= 282912;
srom_1(2367) <= 449758;
srom_1(2368) <= 653832;
srom_1(2369) <= 894177;
srom_1(2370) <= 1169666;
srom_1(2371) <= 1479007;
srom_1(2372) <= 1820750;
srom_1(2373) <= 2193291;
srom_1(2374) <= 2594885;
srom_1(2375) <= 3023647;
srom_1(2376) <= 3477567;
srom_1(2377) <= 3954517;
srom_1(2378) <= 4452260;
srom_1(2379) <= 4968462;
srom_1(2380) <= 5500702;
srom_1(2381) <= 6046484;
srom_1(2382) <= 6603250;
srom_1(2383) <= 7168387;
srom_1(2384) <= 7739247;
srom_1(2385) <= 8313151;
srom_1(2386) <= 8887410;
srom_1(2387) <= 9459329;
srom_1(2388) <= 10026228;
srom_1(2389) <= 10585447;
srom_1(2390) <= 11134364;
srom_1(2391) <= 11670406;
srom_1(2392) <= 12191058;
srom_1(2393) <= 12693879;
srom_1(2394) <= 13176511;
srom_1(2395) <= 13636691;
srom_1(2396) <= 14072261;
srom_1(2397) <= 14481178;
srom_1(2398) <= 14861525;
srom_1(2399) <= 15211519;
srom_1(2400) <= 15529517;
srom_1(2401) <= 15814029;
srom_1(2402) <= 16063721;
srom_1(2403) <= 16277422;
srom_1(2404) <= 16454129;
srom_1(2405) <= 16593014;
srom_1(2406) <= 16693426;
srom_1(2407) <= 16754894;
srom_1(2408) <= 16777130;
srom_1(2409) <= 16760028;
srom_1(2410) <= 16703671;
srom_1(2411) <= 16608321;
srom_1(2412) <= 16474426;
srom_1(2413) <= 16302614;
srom_1(2414) <= 16093690;
srom_1(2415) <= 15848635;
srom_1(2416) <= 15568597;
srom_1(2417) <= 15254889;
srom_1(2418) <= 14908983;
srom_1(2419) <= 14532501;
srom_1(2420) <= 14127208;
srom_1(2421) <= 13695005;
srom_1(2422) <= 13237918;
srom_1(2423) <= 12758091;
srom_1(2424) <= 12257774;
srom_1(2425) <= 11739314;
srom_1(2426) <= 11205140;
srom_1(2427) <= 10657759;
srom_1(2428) <= 10099737;
srom_1(2429) <= 9533691;
srom_1(2430) <= 8962276;
srom_1(2431) <= 8388170;
srom_1(2432) <= 7814066;
srom_1(2433) <= 7242657;
srom_1(2434) <= 6676621;
srom_1(2435) <= 6118613;
srom_1(2436) <= 5571250;
srom_1(2437) <= 5037099;
srom_1(2438) <= 4518664;
srom_1(2439) <= 4018376;
srom_1(2440) <= 3538582;
srom_1(2441) <= 3081532;
srom_1(2442) <= 2649368;
srom_1(2443) <= 2244117;
srom_1(2444) <= 1867680;
srom_1(2445) <= 1521822;
srom_1(2446) <= 1208165;
srom_1(2447) <= 928179;
srom_1(2448) <= 683178;
srom_1(2449) <= 474310;
srom_1(2450) <= 302555;
srom_1(2451) <= 168718;
srom_1(2452) <= 73427;
srom_1(2453) <= 17129;
srom_1(2454) <= 87;
srom_1(2455) <= 22383;
srom_1(2456) <= 83910;
srom_1(2457) <= 184381;
srom_1(2458) <= 323324;
srom_1(2459) <= 500088;
srom_1(2460) <= 713844;
srom_1(2461) <= 963590;
srom_1(2462) <= 1248154;
srom_1(2463) <= 1566203;
srom_1(2464) <= 1916243;
srom_1(2465) <= 2296635;
srom_1(2466) <= 2705595;
srom_1(2467) <= 3141204;
srom_1(2468) <= 3601419;
srom_1(2469) <= 4084084;
srom_1(2470) <= 4586934;
srom_1(2471) <= 5107611;
srom_1(2472) <= 5643674;
srom_1(2473) <= 6192609;
srom_1(2474) <= 6751842;
srom_1(2475) <= 7318750;
srom_1(2476) <= 7890675;
srom_1(2477) <= 8464935;
srom_1(2478) <= 9038837;
srom_1(2479) <= 9609690;
srom_1(2480) <= 10174817;
srom_1(2481) <= 10731567;
srom_1(2482) <= 11277331;
srom_1(2483) <= 11809548;
srom_1(2484) <= 12325724;
srom_1(2485) <= 12823437;
srom_1(2486) <= 13300354;
srom_1(2487) <= 13754237;
srom_1(2488) <= 14182960;
srom_1(2489) <= 14584510;
srom_1(2490) <= 14957006;
srom_1(2491) <= 15298701;
srom_1(2492) <= 15607992;
srom_1(2493) <= 15883428;
srom_1(2494) <= 16123719;
srom_1(2495) <= 16327737;
srom_1(2496) <= 16494526;
srom_1(2497) <= 16623303;
srom_1(2498) <= 16713465;
srom_1(2499) <= 16764589;
srom_1(2500) <= 16776435;
srom_1(2501) <= 16748948;
srom_1(2502) <= 16682256;
srom_1(2503) <= 16576672;
srom_1(2504) <= 16432692;
srom_1(2505) <= 16250990;
srom_1(2506) <= 16032419;
srom_1(2507) <= 15778003;
srom_1(2508) <= 15488936;
srom_1(2509) <= 15166573;
srom_1(2510) <= 14812426;
srom_1(2511) <= 14428156;
srom_1(2512) <= 14015563;
srom_1(2513) <= 13576585;
srom_1(2514) <= 13113277;
srom_1(2515) <= 12627815;
srom_1(2516) <= 12122473;
srom_1(2517) <= 11599622;
srom_1(2518) <= 11061713;
srom_1(2519) <= 10511269;
srom_1(2520) <= 9950871;
srom_1(2521) <= 9383147;
srom_1(2522) <= 8810760;
srom_1(2523) <= 8236393;
srom_1(2524) <= 7662739;
srom_1(2525) <= 7092490;
srom_1(2526) <= 6528318;
srom_1(2527) <= 5972870;
srom_1(2528) <= 5428750;
srom_1(2529) <= 4898510;
srom_1(2530) <= 4384637;
srom_1(2531) <= 3889539;
srom_1(2532) <= 3415539;
srom_1(2533) <= 2964859;
srom_1(2534) <= 2539613;
srom_1(2535) <= 2141795;
srom_1(2536) <= 1773271;
srom_1(2537) <= 1435768;
srom_1(2538) <= 1130869;
srom_1(2539) <= 860004;
srom_1(2540) <= 624444;
srom_1(2541) <= 425292;
srom_1(2542) <= 263483;
srom_1(2543) <= 139776;
srom_1(2544) <= 54750;
srom_1(2545) <= 8805;
srom_1(2546) <= 2155;
srom_1(2547) <= 34832;
srom_1(2548) <= 106683;
srom_1(2549) <= 217371;
srom_1(2550) <= 366376;
srom_1(2551) <= 553001;
srom_1(2552) <= 776369;
srom_1(2553) <= 1035434;
srom_1(2554) <= 1328980;
srom_1(2555) <= 1655631;
srom_1(2556) <= 2013856;
srom_1(2557) <= 2401974;
srom_1(2558) <= 2818165;
srom_1(2559) <= 3260478;
srom_1(2560) <= 3726839;
srom_1(2561) <= 4215060;
srom_1(2562) <= 4722852;
srom_1(2563) <= 5247834;
srom_1(2564) <= 5787545;
srom_1(2565) <= 6339453;
srom_1(2566) <= 6900970;
srom_1(2567) <= 7469463;
srom_1(2568) <= 8042266;
srom_1(2569) <= 8616693;
srom_1(2570) <= 9190051;
srom_1(2571) <= 9759650;
srom_1(2572) <= 10322821;
srom_1(2573) <= 10876921;
srom_1(2574) <= 11419352;
srom_1(2575) <= 11947571;
srom_1(2576) <= 12459101;
srom_1(2577) <= 12951543;
srom_1(2578) <= 13422588;
srom_1(2579) <= 13870027;
srom_1(2580) <= 14291762;
srom_1(2581) <= 14685814;
srom_1(2582) <= 15050337;
srom_1(2583) <= 15383621;
srom_1(2584) <= 15684102;
srom_1(2585) <= 15950373;
srom_1(2586) <= 16181184;
srom_1(2587) <= 16375453;
srom_1(2588) <= 16532268;
srom_1(2589) <= 16650896;
srom_1(2590) <= 16730778;
srom_1(2591) <= 16771542;
srom_1(2592) <= 16772995;
srom_1(2593) <= 16735130;
srom_1(2594) <= 16658126;
srom_1(2595) <= 16542343;
srom_1(2596) <= 16388325;
srom_1(2597) <= 16196793;
srom_1(2598) <= 15968646;
srom_1(2599) <= 15704953;
srom_1(2600) <= 15406952;
srom_1(2601) <= 15076039;
srom_1(2602) <= 14713766;
srom_1(2603) <= 14321833;
srom_1(2604) <= 13902077;
srom_1(2605) <= 13456466;
srom_1(2606) <= 12987090;
srom_1(2607) <= 12496150;
srom_1(2608) <= 11985949;
srom_1(2609) <= 11458878;
srom_1(2610) <= 10917410;
srom_1(2611) <= 10364084;
srom_1(2612) <= 9801494;
srom_1(2613) <= 9232278;
srom_1(2614) <= 8659106;
srom_1(2615) <= 8084666;
srom_1(2616) <= 7511650;
srom_1(2617) <= 6942748;
srom_1(2618) <= 6380625;
srom_1(2619) <= 5827918;
srom_1(2620) <= 5287220;
srom_1(2621) <= 4761065;
srom_1(2622) <= 4251920;
srom_1(2623) <= 3762174;
srom_1(2624) <= 3294123;
srom_1(2625) <= 2849962;
srom_1(2626) <= 2431773;
srom_1(2627) <= 2041518;
srom_1(2628) <= 1681027;
srom_1(2629) <= 1351989;
srom_1(2630) <= 1055949;
srom_1(2631) <= 794294;
srom_1(2632) <= 568252;
srom_1(2633) <= 378882;
srom_1(2634) <= 227072;
srom_1(2635) <= 113535;
srom_1(2636) <= 38802;
srom_1(2637) <= 3224;
srom_1(2638) <= 6968;
srom_1(2639) <= 50017;
srom_1(2640) <= 132168;
srom_1(2641) <= 253036;
srom_1(2642) <= 412055;
srom_1(2643) <= 608479;
srom_1(2644) <= 841386;
srom_1(2645) <= 1109685;
srom_1(2646) <= 1412117;
srom_1(2647) <= 1747264;
srom_1(2648) <= 2113555;
srom_1(2649) <= 2509272;
srom_1(2650) <= 2932559;
srom_1(2651) <= 3381431;
srom_1(2652) <= 3853784;
srom_1(2653) <= 4347402;
srom_1(2654) <= 4859970;
srom_1(2655) <= 5389086;
srom_1(2656) <= 5932267;
srom_1(2657) <= 6486967;
srom_1(2658) <= 7050585;
srom_1(2659) <= 7620476;
srom_1(2660) <= 8193970;
srom_1(2661) <= 8768377;
srom_1(2662) <= 9341003;
srom_1(2663) <= 9909162;
srom_1(2664) <= 10470191;
srom_1(2665) <= 11021459;
srom_1(2666) <= 11560381;
srom_1(2667) <= 12084429;
srom_1(2668) <= 12591146;
srom_1(2669) <= 13078156;
srom_1(2670) <= 13543175;
srom_1(2671) <= 13984022;
srom_1(2672) <= 14398631;
srom_1(2673) <= 14785056;
srom_1(2674) <= 15141487;
srom_1(2675) <= 15466251;
srom_1(2676) <= 15757825;
srom_1(2677) <= 16014842;
srom_1(2678) <= 16236098;
srom_1(2679) <= 16420554;
srom_1(2680) <= 16567345;
srom_1(2681) <= 16675784;
srom_1(2682) <= 16745361;
srom_1(2683) <= 16775750;
srom_1(2684) <= 16766809;
srom_1(2685) <= 16718580;
srom_1(2686) <= 16631289;
srom_1(2687) <= 16505344;
srom_1(2688) <= 16341338;
srom_1(2689) <= 16140039;
srom_1(2690) <= 15902391;
srom_1(2691) <= 15629507;
srom_1(2692) <= 15322669;
srom_1(2693) <= 14983315;
srom_1(2694) <= 14613035;
srom_1(2695) <= 14213568;
srom_1(2696) <= 13786785;
srom_1(2697) <= 13334688;
srom_1(2698) <= 12859397;
srom_1(2699) <= 12363141;
srom_1(2700) <= 11848247;
srom_1(2701) <= 11317130;
srom_1(2702) <= 10772280;
srom_1(2703) <= 10216252;
srom_1(2704) <= 9651654;
srom_1(2705) <= 9081132;
srom_1(2706) <= 8507363;
srom_1(2707) <= 7933038;
srom_1(2708) <= 7360848;
srom_1(2709) <= 6793479;
srom_1(2710) <= 6233589;
srom_1(2711) <= 5683805;
srom_1(2712) <= 5146704;
srom_1(2713) <= 4624806;
srom_1(2714) <= 4120558;
srom_1(2715) <= 3636324;
srom_1(2716) <= 3174375;
srom_1(2717) <= 2736878;
srom_1(2718) <= 2325883;
srom_1(2719) <= 1943319;
srom_1(2720) <= 1590979;
srom_1(2721) <= 1270515;
srom_1(2722) <= 983430;
srom_1(2723) <= 731071;
srom_1(2724) <= 514621;
srom_1(2725) <= 335094;
srom_1(2726) <= 193333;
srom_1(2727) <= 90003;
srom_1(2728) <= 25587;
srom_1(2729) <= 389;
srom_1(2730) <= 14526;
srom_1(2731) <= 67931;
srom_1(2732) <= 160356;
srom_1(2733) <= 291365;
srom_1(2734) <= 460345;
srom_1(2735) <= 666504;
srom_1(2736) <= 908874;
srom_1(2737) <= 1186319;
srom_1(2738) <= 1497538;
srom_1(2739) <= 1841072;
srom_1(2740) <= 2215309;
srom_1(2741) <= 2618495;
srom_1(2742) <= 3048739;
srom_1(2743) <= 3504024;
srom_1(2744) <= 3982214;
srom_1(2745) <= 4481067;
srom_1(2746) <= 4998244;
srom_1(2747) <= 5531320;
srom_1(2748) <= 6077794;
srom_1(2749) <= 6635104;
srom_1(2750) <= 7200638;
srom_1(2751) <= 7771742;
srom_1(2752) <= 8345738;
srom_1(2753) <= 8919936;
srom_1(2754) <= 9491642;
srom_1(2755) <= 10058176;
srom_1(2756) <= 10616881;
srom_1(2757) <= 11165136;
srom_1(2758) <= 11700371;
srom_1(2759) <= 12220076;
srom_1(2760) <= 12721815;
srom_1(2761) <= 13203233;
srom_1(2762) <= 13662074;
srom_1(2763) <= 14096186;
srom_1(2764) <= 14503532;
srom_1(2765) <= 14882204;
srom_1(2766) <= 15230426;
srom_1(2767) <= 15546563;
srom_1(2768) <= 15829135;
srom_1(2769) <= 16076815;
srom_1(2770) <= 16288443;
srom_1(2771) <= 16463025;
srom_1(2772) <= 16599744;
srom_1(2773) <= 16697958;
srom_1(2774) <= 16757207;
srom_1(2775) <= 16777212;
srom_1(2776) <= 16757880;
srom_1(2777) <= 16699302;
srom_1(2778) <= 16601753;
srom_1(2779) <= 16465688;
srom_1(2780) <= 16291748;
srom_1(2781) <= 16080747;
srom_1(2782) <= 15833675;
srom_1(2783) <= 15551691;
srom_1(2784) <= 15236117;
srom_1(2785) <= 14888432;
srom_1(2786) <= 14510267;
srom_1(2787) <= 14103395;
srom_1(2788) <= 13669726;
srom_1(2789) <= 13211291;
srom_1(2790) <= 12730240;
srom_1(2791) <= 12228831;
srom_1(2792) <= 11709413;
srom_1(2793) <= 11174423;
srom_1(2794) <= 10626369;
srom_1(2795) <= 10067822;
srom_1(2796) <= 9501400;
srom_1(2797) <= 8929760;
srom_1(2798) <= 8355582;
srom_1(2799) <= 7781559;
srom_1(2800) <= 7210383;
srom_1(2801) <= 6644732;
srom_1(2802) <= 6087258;
srom_1(2803) <= 5540577;
srom_1(2804) <= 5007250;
srom_1(2805) <= 4489780;
srom_1(2806) <= 3990593;
srom_1(2807) <= 3512030;
srom_1(2808) <= 3056335;
srom_1(2809) <= 2625644;
srom_1(2810) <= 2221978;
srom_1(2811) <= 1847230;
srom_1(2812) <= 1503156;
srom_1(2813) <= 1191371;
srom_1(2814) <= 913335;
srom_1(2815) <= 670354;
srom_1(2816) <= 463567;
srom_1(2817) <= 293943;
srom_1(2818) <= 162277;
srom_1(2819) <= 69187;
srom_1(2820) <= 15110;
srom_1(2821) <= 300;
srom_1(2822) <= 24825;
srom_1(2823) <= 88570;
srom_1(2824) <= 191237;
srom_1(2825) <= 332345;
srom_1(2826) <= 511231;
srom_1(2827) <= 727057;
srom_1(2828) <= 978811;
srom_1(2829) <= 1265311;
srom_1(2830) <= 1585215;
srom_1(2831) <= 1937023;
srom_1(2832) <= 2319084;
srom_1(2833) <= 2729608;
srom_1(2834) <= 3166668;
srom_1(2835) <= 3628216;
srom_1(2836) <= 4112087;
srom_1(2837) <= 4616012;
srom_1(2838) <= 5137628;
srom_1(2839) <= 5674489;
srom_1(2840) <= 6224077;
srom_1(2841) <= 6783816;
srom_1(2842) <= 7351080;
srom_1(2843) <= 7923209;
srom_1(2844) <= 8497521;
srom_1(2845) <= 9071322;
srom_1(2846) <= 9641921;
srom_1(2847) <= 10206643;
srom_1(2848) <= 10762840;
srom_1(2849) <= 11307904;
srom_1(2850) <= 11839277;
srom_1(2851) <= 12354470;
srom_1(2852) <= 12851065;
srom_1(2853) <= 13326734;
srom_1(2854) <= 13779246;
srom_1(2855) <= 14206480;
srom_1(2856) <= 14606432;
srom_1(2857) <= 14977226;
srom_1(2858) <= 15317125;
srom_1(2859) <= 15624532;
srom_1(2860) <= 15898009;
srom_1(2861) <= 16136270;
srom_1(2862) <= 16338201;
srom_1(2863) <= 16502853;
srom_1(2864) <= 16629455;
srom_1(2865) <= 16717412;
srom_1(2866) <= 16766313;
srom_1(2867) <= 16775928;
srom_1(2868) <= 16746212;
srom_1(2869) <= 16677304;
srom_1(2870) <= 16569528;
srom_1(2871) <= 16423388;
srom_1(2872) <= 16239571;
srom_1(2873) <= 16018937;
srom_1(2874) <= 15762523;
srom_1(2875) <= 15471530;
srom_1(2876) <= 15147322;
srom_1(2877) <= 14791421;
srom_1(2878) <= 14405494;
srom_1(2879) <= 13991352;
srom_1(2880) <= 13550937;
srom_1(2881) <= 13086314;
srom_1(2882) <= 12599662;
srom_1(2883) <= 12093263;
srom_1(2884) <= 11569492;
srom_1(2885) <= 11030804;
srom_1(2886) <= 10479726;
srom_1(2887) <= 9918842;
srom_1(2888) <= 9350782;
srom_1(2889) <= 8778210;
srom_1(2890) <= 8203812;
srom_1(2891) <= 7630279;
srom_1(2892) <= 7060303;
srom_1(2893) <= 6496556;
srom_1(2894) <= 5941681;
srom_1(2895) <= 5398281;
srom_1(2896) <= 4868903;
srom_1(2897) <= 4356031;
srom_1(2898) <= 3862068;
srom_1(2899) <= 3389332;
srom_1(2900) <= 2940040;
srom_1(2901) <= 2516298;
srom_1(2902) <= 2120092;
srom_1(2903) <= 1753282;
srom_1(2904) <= 1417588;
srom_1(2905) <= 1114583;
srom_1(2906) <= 845688;
srom_1(2907) <= 612165;
srom_1(2908) <= 415108;
srom_1(2909) <= 255441;
srom_1(2910) <= 133914;
srom_1(2911) <= 51096;
srom_1(2912) <= 7375;
srom_1(2913) <= 2957;
srom_1(2914) <= 37862;
srom_1(2915) <= 111926;
srom_1(2916) <= 224803;
srom_1(2917) <= 375962;
srom_1(2918) <= 564696;
srom_1(2919) <= 790119;
srom_1(2920) <= 1051173;
srom_1(2921) <= 1346635;
srom_1(2922) <= 1675120;
srom_1(2923) <= 2035086;
srom_1(2924) <= 2424846;
srom_1(2925) <= 2842573;
srom_1(2926) <= 3286306;
srom_1(2927) <= 3753966;
srom_1(2928) <= 4243359;
srom_1(2929) <= 4752191;
srom_1(2930) <= 5278076;
srom_1(2931) <= 5818546;
srom_1(2932) <= 6371069;
srom_1(2933) <= 6933052;
srom_1(2934) <= 7501861;
srom_1(2935) <= 8074828;
srom_1(2936) <= 8649267;
srom_1(2937) <= 9222484;
srom_1(2938) <= 9791790;
srom_1(2939) <= 10354516;
srom_1(2940) <= 10908023;
srom_1(2941) <= 11449716;
srom_1(2942) <= 11977054;
srom_1(2943) <= 12487565;
srom_1(2944) <= 12978854;
srom_1(2945) <= 13448618;
srom_1(2946) <= 13894654;
srom_1(2947) <= 14314870;
srom_1(2948) <= 14707296;
srom_1(2949) <= 15070091;
srom_1(2950) <= 15401555;
srom_1(2951) <= 15700133;
srom_1(2952) <= 15964424;
srom_1(2953) <= 16193189;
srom_1(2954) <= 16385357;
srom_1(2955) <= 16540024;
srom_1(2956) <= 16656467;
srom_1(2957) <= 16734140;
srom_1(2958) <= 16772677;
srom_1(2959) <= 16771898;
srom_1(2960) <= 16731807;
srom_1(2961) <= 16652592;
srom_1(2962) <= 16534624;
srom_1(2963) <= 16378457;
srom_1(2964) <= 16184823;
srom_1(2965) <= 15954629;
srom_1(2966) <= 15688956;
srom_1(2967) <= 15389049;
srom_1(2968) <= 15056315;
srom_1(2969) <= 14692313;
srom_1(2970) <= 14298751;
srom_1(2971) <= 13877475;
srom_1(2972) <= 13430459;
srom_1(2973) <= 12959800;
srom_1(2974) <= 12467706;
srom_1(2975) <= 11956483;
srom_1(2976) <= 11428529;
srom_1(2977) <= 10886320;
srom_1(2978) <= 10332398;
srom_1(2979) <= 9769361;
srom_1(2980) <= 9199849;
srom_1(2981) <= 8626533;
srom_1(2982) <= 8052101;
srom_1(2983) <= 7479248;
srom_1(2984) <= 6910658;
srom_1(2985) <= 6349000;
srom_1(2986) <= 5796905;
srom_1(2987) <= 5256964;
srom_1(2988) <= 4731709;
srom_1(2989) <= 4223601;
srom_1(2990) <= 3735025;
srom_1(2991) <= 3268272;
srom_1(2992) <= 2825529;
srom_1(2993) <= 2408873;
srom_1(2994) <= 2020259;
srom_1(2995) <= 1661507;
srom_1(2996) <= 1334302;
srom_1(2997) <= 1040176;
srom_1(2998) <= 780510;
srom_1(2999) <= 556521;
srom_1(3000) <= 369259;
srom_1(3001) <= 219603;
srom_1(3002) <= 108254;
srom_1(3003) <= 35734;
srom_1(3004) <= 2384;
srom_1(3005) <= 8360;
srom_1(3006) <= 53633;
srom_1(3007) <= 137992;
srom_1(3008) <= 261041;
srom_1(3009) <= 422203;
srom_1(3010) <= 620722;
srom_1(3011) <= 855668;
srom_1(3012) <= 1125938;
srom_1(3013) <= 1430265;
srom_1(3014) <= 1767222;
srom_1(3015) <= 2135229;
srom_1(3016) <= 2532561;
srom_1(3017) <= 2957353;
srom_1(3018) <= 3407615;
srom_1(3019) <= 3881234;
srom_1(3020) <= 4375989;
srom_1(3021) <= 4889561;
srom_1(3022) <= 5419542;
srom_1(3023) <= 5963445;
srom_1(3024) <= 6518721;
srom_1(3025) <= 7082765;
srom_1(3026) <= 7652933;
srom_1(3027) <= 8226551;
srom_1(3028) <= 8800928;
srom_1(3029) <= 9373372;
srom_1(3030) <= 9941199;
srom_1(3031) <= 10501744;
srom_1(3032) <= 11052380;
srom_1(3033) <= 11590525;
srom_1(3034) <= 12113655;
srom_1(3035) <= 12619317;
srom_1(3036) <= 13105140;
srom_1(3037) <= 13568846;
srom_1(3038) <= 14008259;
srom_1(3039) <= 14421320;
srom_1(3040) <= 14806091;
srom_1(3041) <= 15160769;
srom_1(3042) <= 15483690;
srom_1(3043) <= 15773339;
srom_1(3044) <= 16028359;
srom_1(3045) <= 16247553;
srom_1(3046) <= 16429894;
srom_1(3047) <= 16574527;
srom_1(3048) <= 16680773;
srom_1(3049) <= 16748135;
srom_1(3050) <= 16776295;
srom_1(3051) <= 16765123;
srom_1(3052) <= 16714671;
srom_1(3053) <= 16625174;
srom_1(3054) <= 16497054;
srom_1(3055) <= 16330910;
srom_1(3056) <= 16127523;
srom_1(3057) <= 15887844;
srom_1(3058) <= 15612999;
srom_1(3059) <= 15304277;
srom_1(3060) <= 14963125;
srom_1(3061) <= 14591142;
srom_1(3062) <= 14190074;
srom_1(3063) <= 13761800;
srom_1(3064) <= 13308330;
srom_1(3065) <= 12831789;
srom_1(3066) <= 12334413;
srom_1(3067) <= 11818534;
srom_1(3068) <= 11286571;
srom_1(3069) <= 10741018;
srom_1(3070) <= 10184433;
srom_1(3071) <= 9619428;
srom_1(3072) <= 9048651;
srom_1(3073) <= 8474778;
srom_1(3074) <= 7900502;
srom_1(3075) <= 7328514;
srom_1(3076) <= 6761497;
srom_1(3077) <= 6202111;
srom_1(3078) <= 5652978;
srom_1(3079) <= 5116673;
srom_1(3080) <= 4595711;
srom_1(3081) <= 4092536;
srom_1(3082) <= 3609506;
srom_1(3083) <= 3148887;
srom_1(3084) <= 2712839;
srom_1(3085) <= 2303407;
srom_1(3086) <= 1922510;
srom_1(3087) <= 1571935;
srom_1(3088) <= 1253325;
srom_1(3089) <= 968176;
srom_1(3090) <= 717823;
srom_1(3091) <= 503442;
srom_1(3092) <= 326036;
srom_1(3093) <= 186439;
srom_1(3094) <= 85304;
srom_1(3095) <= 23107;
srom_1(3096) <= 138;
srom_1(3097) <= 16506;
srom_1(3098) <= 72133;
srom_1(3099) <= 166759;
srom_1(3100) <= 299940;
srom_1(3101) <= 471052;
srom_1(3102) <= 679292;
srom_1(3103) <= 923683;
srom_1(3104) <= 1203080;
srom_1(3105) <= 1516173;
srom_1(3106) <= 1861493;
srom_1(3107) <= 2237420;
srom_1(3108) <= 2642193;
srom_1(3109) <= 3073912;
srom_1(3110) <= 3530554;
srom_1(3111) <= 4009977;
srom_1(3112) <= 4509933;
srom_1(3113) <= 5028077;
srom_1(3114) <= 5561980;
srom_1(3115) <= 6109138;
srom_1(3116) <= 6666985;
srom_1(3117) <= 7232906;
srom_1(3118) <= 7804246;
srom_1(3119) <= 8378326;
srom_1(3120) <= 8952455;
srom_1(3121) <= 9523939;
srom_1(3122) <= 10090099;
srom_1(3123) <= 10648281;
srom_1(3124) <= 11195866;
srom_1(3125) <= 11730287;
srom_1(3126) <= 12249038;
srom_1(3127) <= 12749685;
srom_1(3128) <= 13229882;
srom_1(3129) <= 13687377;
srom_1(3130) <= 14120024;
srom_1(3131) <= 14525795;
srom_1(3132) <= 14902786;
srom_1(3133) <= 15249229;
srom_1(3134) <= 15563501;
srom_1(3135) <= 15844128;
srom_1(3136) <= 16089793;
srom_1(3137) <= 16299344;
srom_1(3138) <= 16471799;
srom_1(3139) <= 16606350;
srom_1(3140) <= 16702364;
srom_1(3141) <= 16759393;
srom_1(3142) <= 16777168;
srom_1(3143) <= 16755606;
srom_1(3144) <= 16694808;
srom_1(3145) <= 16595060;
srom_1(3146) <= 16456829;
srom_1(3147) <= 16280763;
srom_1(3148) <= 16067689;
srom_1(3149) <= 15818604;
srom_1(3150) <= 15534677;
srom_1(3151) <= 15217241;
srom_1(3152) <= 14867782;
srom_1(3153) <= 14487940;
srom_1(3154) <= 14079497;
srom_1(3155) <= 13644367;
srom_1(3156) <= 13184590;
srom_1(3157) <= 12702324;
srom_1(3158) <= 12199829;
srom_1(3159) <= 11679462;
srom_1(3160) <= 11143664;
srom_1(3161) <= 10594945;
srom_1(3162) <= 10035881;
srom_1(3163) <= 9469092;
srom_1(3164) <= 8897236;
srom_1(3165) <= 8322995;
srom_1(3166) <= 7749061;
srom_1(3167) <= 7178127;
srom_1(3168) <= 6612869;
srom_1(3169) <= 6055938;
srom_1(3170) <= 5509946;
srom_1(3171) <= 4977453;
srom_1(3172) <= 4460956;
srom_1(3173) <= 3962877;
srom_1(3174) <= 3485551;
srom_1(3175) <= 3031218;
srom_1(3176) <= 2602008;
srom_1(3177) <= 2199932;
srom_1(3178) <= 1826878;
srom_1(3179) <= 1484594;
srom_1(3180) <= 1174685;
srom_1(3181) <= 898605;
srom_1(3182) <= 657648;
srom_1(3183) <= 452944;
srom_1(3184) <= 285453;
srom_1(3185) <= 155960;
srom_1(3186) <= 65073;
srom_1(3187) <= 13219;
srom_1(3188) <= 639;
srom_1(3189) <= 27393;
srom_1(3190) <= 93356;
srom_1(3191) <= 198218;
srom_1(3192) <= 341488;
srom_1(3193) <= 522493;
srom_1(3194) <= 740385;
srom_1(3195) <= 994143;
srom_1(3196) <= 1282575;
srom_1(3197) <= 1604331;
srom_1(3198) <= 1957900;
srom_1(3199) <= 2341625;
srom_1(3200) <= 2753706;
srom_1(3201) <= 3192211;
srom_1(3202) <= 3655084;
srom_1(3203) <= 4140154;
srom_1(3204) <= 4645146;
srom_1(3205) <= 5167693;
srom_1(3206) <= 5705344;
srom_1(3207) <= 6255577;
srom_1(3208) <= 6815814;
srom_1(3209) <= 7383425;
srom_1(3210) <= 7955750;
srom_1(3211) <= 8530105;
srom_1(3212) <= 9103796;
srom_1(3213) <= 9674134;
srom_1(3214) <= 10238443;
srom_1(3215) <= 10794078;
srom_1(3216) <= 11338432;
srom_1(3217) <= 11868954;
srom_1(3218) <= 12383156;
srom_1(3219) <= 12878625;
srom_1(3220) <= 13353040;
srom_1(3221) <= 13804174;
srom_1(3222) <= 14229913;
srom_1(3223) <= 14628260;
srom_1(3224) <= 14997347;
srom_1(3225) <= 15335444;
srom_1(3226) <= 15640964;
srom_1(3227) <= 15912476;
srom_1(3228) <= 16148705;
srom_1(3229) <= 16348545;
srom_1(3230) <= 16511058;
srom_1(3231) <= 16635482;
srom_1(3232) <= 16721234;
srom_1(3233) <= 16767911;
srom_1(3234) <= 16775294;
srom_1(3235) <= 16743350;
srom_1(3236) <= 16672227;
srom_1(3237) <= 16562259;
srom_1(3238) <= 16413963;
srom_1(3239) <= 16228033;
srom_1(3240) <= 16005341;
srom_1(3241) <= 15746931;
srom_1(3242) <= 15454016;
srom_1(3243) <= 15127969;
srom_1(3244) <= 14770318;
srom_1(3245) <= 14382742;
srom_1(3246) <= 13967057;
srom_1(3247) <= 13525212;
srom_1(3248) <= 13059280;
srom_1(3249) <= 12571446;
srom_1(3250) <= 12063998;
srom_1(3251) <= 11539314;
srom_1(3252) <= 10999855;
srom_1(3253) <= 10448151;
srom_1(3254) <= 9886789;
srom_1(3255) <= 9318402;
srom_1(3256) <= 8745655;
srom_1(3257) <= 8171233;
srom_1(3258) <= 7597831;
srom_1(3259) <= 7028137;
srom_1(3260) <= 6464822;
srom_1(3261) <= 5910529;
srom_1(3262) <= 5367857;
srom_1(3263) <= 4839349;
srom_1(3264) <= 4327486;
srom_1(3265) <= 3834666;
srom_1(3266) <= 3363202;
srom_1(3267) <= 2915303;
srom_1(3268) <= 2493071;
srom_1(3269) <= 2098484;
srom_1(3270) <= 1733395;
srom_1(3271) <= 1399513;
srom_1(3272) <= 1098406;
srom_1(3273) <= 831486;
srom_1(3274) <= 600003;
srom_1(3275) <= 405044;
srom_1(3276) <= 247522;
srom_1(3277) <= 128177;
srom_1(3278) <= 47567;
srom_1(3279) <= 6072;
srom_1(3280) <= 3885;
srom_1(3281) <= 41018;
srom_1(3282) <= 117294;
srom_1(3283) <= 232358;
srom_1(3284) <= 385670;
srom_1(3285) <= 576509;
srom_1(3286) <= 803983;
srom_1(3287) <= 1067023;
srom_1(3288) <= 1364397;
srom_1(3289) <= 1694710;
srom_1(3290) <= 2056412;
srom_1(3291) <= 2447809;
srom_1(3292) <= 2867064;
srom_1(3293) <= 3312211;
srom_1(3294) <= 3781163;
srom_1(3295) <= 4271722;
srom_1(3296) <= 4781585;
srom_1(3297) <= 5308364;
srom_1(3298) <= 5849586;
srom_1(3299) <= 6402715;
srom_1(3300) <= 6965157;
srom_1(3301) <= 7534273;
srom_1(3302) <= 8107396;
srom_1(3303) <= 8681837;
srom_1(3304) <= 9254904;
srom_1(3305) <= 9823908;
srom_1(3306) <= 10386181;
srom_1(3307) <= 10939087;
srom_1(3308) <= 11480033;
srom_1(3309) <= 12006482;
srom_1(3310) <= 12515966;
srom_1(3311) <= 13006095;
srom_1(3312) <= 13474571;
srom_1(3313) <= 13919198;
srom_1(3314) <= 14337889;
srom_1(3315) <= 14728683;
srom_1(3316) <= 15089745;
srom_1(3317) <= 15419384;
srom_1(3318) <= 15716052;
srom_1(3319) <= 15978360;
srom_1(3320) <= 16205077;
srom_1(3321) <= 16395140;
srom_1(3322) <= 16547657;
srom_1(3323) <= 16661914;
srom_1(3324) <= 16737375;
srom_1(3325) <= 16773685;
srom_1(3326) <= 16770675;
srom_1(3327) <= 16728358;
srom_1(3328) <= 16646933;
srom_1(3329) <= 16526782;
srom_1(3330) <= 16368469;
srom_1(3331) <= 16172735;
srom_1(3332) <= 15940499;
srom_1(3333) <= 15672849;
srom_1(3334) <= 15371041;
srom_1(3335) <= 15036490;
srom_1(3336) <= 14670765;
srom_1(3337) <= 14275580;
srom_1(3338) <= 13852790;
srom_1(3339) <= 13404376;
srom_1(3340) <= 12932441;
srom_1(3341) <= 12439199;
srom_1(3342) <= 11926962;
srom_1(3343) <= 11398133;
srom_1(3344) <= 10855191;
srom_1(3345) <= 10300682;
srom_1(3346) <= 9737207;
srom_1(3347) <= 9167408;
srom_1(3348) <= 8593957;
srom_1(3349) <= 8019542;
srom_1(3350) <= 7446859;
srom_1(3351) <= 6878592;
srom_1(3352) <= 6317405;
srom_1(3353) <= 5765931;
srom_1(3354) <= 5226756;
srom_1(3355) <= 4702408;
srom_1(3356) <= 4195346;
srom_1(3357) <= 3707947;
srom_1(3358) <= 3242498;
srom_1(3359) <= 2801180;
srom_1(3360) <= 2386064;
srom_1(3361) <= 1999095;
srom_1(3362) <= 1642090;
srom_1(3363) <= 1316721;
srom_1(3364) <= 1024515;
srom_1(3365) <= 766841;
srom_1(3366) <= 544908;
srom_1(3367) <= 359758;
srom_1(3368) <= 212257;
srom_1(3369) <= 103098;
srom_1(3370) <= 32792;
srom_1(3371) <= 1670;
srom_1(3372) <= 9877;
srom_1(3373) <= 57375;
srom_1(3374) <= 143941;
srom_1(3375) <= 269169;
srom_1(3376) <= 432472;
srom_1(3377) <= 633083;
srom_1(3378) <= 870063;
srom_1(3379) <= 1142301;
srom_1(3380) <= 1448518;
srom_1(3381) <= 1787280;
srom_1(3382) <= 2156998;
srom_1(3383) <= 2555938;
srom_1(3384) <= 2982229;
srom_1(3385) <= 3433873;
srom_1(3386) <= 3908751;
srom_1(3387) <= 4404637;
srom_1(3388) <= 4919205;
srom_1(3389) <= 5450043;
srom_1(3390) <= 5994660;
srom_1(3391) <= 6550503;
srom_1(3392) <= 7114966;
srom_1(3393) <= 7685401;
srom_1(3394) <= 8259134;
srom_1(3395) <= 8833474;
srom_1(3396) <= 9405727;
srom_1(3397) <= 9973212;
srom_1(3398) <= 10533265;
srom_1(3399) <= 11083261;
srom_1(3400) <= 11620622;
srom_1(3401) <= 12142826;
srom_1(3402) <= 12647425;
srom_1(3403) <= 13132054;
srom_1(3404) <= 13594438;
srom_1(3405) <= 14032411;
srom_1(3406) <= 14443918;
srom_1(3407) <= 14827029;
srom_1(3408) <= 15179949;
srom_1(3409) <= 15501022;
srom_1(3410) <= 15788742;
srom_1(3411) <= 16041760;
srom_1(3412) <= 16258890;
srom_1(3413) <= 16439114;
srom_1(3414) <= 16581586;
srom_1(3415) <= 16685638;
srom_1(3416) <= 16750783;
srom_1(3417) <= 16776714;
srom_1(3418) <= 16763311;
srom_1(3419) <= 16710636;
srom_1(3420) <= 16618936;
srom_1(3421) <= 16488641;
srom_1(3422) <= 16320363;
srom_1(3423) <= 16114889;
srom_1(3424) <= 15873185;
srom_1(3425) <= 15596383;
srom_1(3426) <= 15285781;
srom_1(3427) <= 14942835;
srom_1(3428) <= 14569155;
srom_1(3429) <= 14166492;
srom_1(3430) <= 13736735;
srom_1(3431) <= 13281898;
srom_1(3432) <= 12804115;
srom_1(3433) <= 12305626;
srom_1(3434) <= 11788769;
srom_1(3435) <= 11255967;
srom_1(3436) <= 10709720;
srom_1(3437) <= 10152588;
srom_1(3438) <= 9587183;
srom_1(3439) <= 9016159;
srom_1(3440) <= 8442191;
srom_1(3441) <= 7867973;
srom_1(3442) <= 7296195;
srom_1(3443) <= 6729541;
srom_1(3444) <= 6170666;
srom_1(3445) <= 5622192;
srom_1(3446) <= 5086691;
srom_1(3447) <= 4566673;
srom_1(3448) <= 4064578;
srom_1(3449) <= 3582760;
srom_1(3450) <= 3123478;
srom_1(3451) <= 2688886;
srom_1(3452) <= 2281022;
srom_1(3453) <= 1901799;
srom_1(3454) <= 1552994;
srom_1(3455) <= 1236244;
srom_1(3456) <= 953034;
srom_1(3457) <= 704691;
srom_1(3458) <= 492382;
srom_1(3459) <= 317100;
srom_1(3460) <= 179668;
srom_1(3461) <= 80731;
srom_1(3462) <= 20753;
srom_1(3463) <= 14;
srom_1(3464) <= 18612;
srom_1(3465) <= 76460;
srom_1(3466) <= 173287;
srom_1(3467) <= 308638;
srom_1(3468) <= 481878;
srom_1(3469) <= 692196;
srom_1(3470) <= 938606;
srom_1(3471) <= 1219950;
srom_1(3472) <= 1534911;
srom_1(3473) <= 1882012;
srom_1(3474) <= 2259624;
srom_1(3475) <= 2665977;
srom_1(3476) <= 3099165;
srom_1(3477) <= 3557157;
srom_1(3478) <= 4037806;
srom_1(3479) <= 4538857;
srom_1(3480) <= 5057961;
srom_1(3481) <= 5592684;
srom_1(3482) <= 6140517;
srom_1(3483) <= 6698892;
srom_1(3484) <= 7265192;
srom_1(3485) <= 7836759;
srom_1(3486) <= 8410914;
srom_1(3487) <= 8984964;
srom_1(3488) <= 9556218;
srom_1(3489) <= 10121997;
srom_1(3490) <= 10679647;
srom_1(3491) <= 11226554;
srom_1(3492) <= 11760152;
srom_1(3493) <= 12277940;
srom_1(3494) <= 12777490;
srom_1(3495) <= 13256459;
srom_1(3496) <= 13712601;
srom_1(3497) <= 14143776;
srom_1(3498) <= 14547964;
srom_1(3499) <= 14923269;
srom_1(3500) <= 15267930;
srom_1(3501) <= 15580331;
srom_1(3502) <= 15859008;
srom_1(3503) <= 16102654;
srom_1(3504) <= 16310126;
srom_1(3505) <= 16480452;
srom_1(3506) <= 16612832;
srom_1(3507) <= 16706645;
srom_1(3508) <= 16761453;
srom_1(3509) <= 16776997;
srom_1(3510) <= 16753205;
srom_1(3511) <= 16690189;
srom_1(3512) <= 16588244;
srom_1(3513) <= 16447848;
srom_1(3514) <= 16269660;
srom_1(3515) <= 16054514;
srom_1(3516) <= 15803420;
srom_1(3517) <= 15517556;
srom_1(3518) <= 15198262;
srom_1(3519) <= 14847035;
srom_1(3520) <= 14465522;
srom_1(3521) <= 14055512;
srom_1(3522) <= 13618928;
srom_1(3523) <= 13157818;
srom_1(3524) <= 12674343;
srom_1(3525) <= 12170770;
srom_1(3526) <= 11649462;
srom_1(3527) <= 11112863;
srom_1(3528) <= 10563488;
srom_1(3529) <= 10003915;
srom_1(3530) <= 9436767;
srom_1(3531) <= 8864704;
srom_1(3532) <= 8290409;
srom_1(3533) <= 7716573;
srom_1(3534) <= 7145890;
srom_1(3535) <= 6581033;
srom_1(3536) <= 6024653;
srom_1(3537) <= 5479359;
srom_1(3538) <= 4947707;
srom_1(3539) <= 4432190;
srom_1(3540) <= 3935227;
srom_1(3541) <= 3459147;
srom_1(3542) <= 3006182;
srom_1(3543) <= 2578458;
srom_1(3544) <= 2177980;
srom_1(3545) <= 1806625;
srom_1(3546) <= 1466136;
srom_1(3547) <= 1158108;
srom_1(3548) <= 883987;
srom_1(3549) <= 645057;
srom_1(3550) <= 442440;
srom_1(3551) <= 277085;
srom_1(3552) <= 149768;
srom_1(3553) <= 61085;
srom_1(3554) <= 11453;
srom_1(3555) <= 1104;
srom_1(3556) <= 30088;
srom_1(3557) <= 98267;
srom_1(3558) <= 205322;
srom_1(3559) <= 350752;
srom_1(3560) <= 533874;
srom_1(3561) <= 753829;
srom_1(3562) <= 1009587;
srom_1(3563) <= 1299947;
srom_1(3564) <= 1623549;
srom_1(3565) <= 1978874;
srom_1(3566) <= 2364256;
srom_1(3567) <= 2777889;
srom_1(3568) <= 3217833;
srom_1(3569) <= 3682024;
srom_1(3570) <= 4168285;
srom_1(3571) <= 4674338;
srom_1(3572) <= 5197807;
srom_1(3573) <= 5736240;
srom_1(3574) <= 6287110;
srom_1(3575) <= 6847835;
srom_1(3576) <= 7415785;
srom_1(3577) <= 7988298;
srom_1(3578) <= 8562687;
srom_1(3579) <= 9136260;
srom_1(3580) <= 9706327;
srom_1(3581) <= 10270215;
srom_1(3582) <= 10825279;
srom_1(3583) <= 11368917;
srom_1(3584) <= 11898579;
srom_1(3585) <= 12411781;
srom_1(3586) <= 12906118;
srom_1(3587) <= 13379270;
srom_1(3588) <= 13829020;
srom_1(3589) <= 14253258;
srom_1(3590) <= 14649994;
srom_1(3591) <= 15017368;
srom_1(3592) <= 15353658;
srom_1(3593) <= 15657286;
srom_1(3594) <= 15926829;
srom_1(3595) <= 16161023;
srom_1(3596) <= 16358769;
srom_1(3597) <= 16519140;
srom_1(3598) <= 16641385;
srom_1(3599) <= 16724929;
srom_1(3600) <= 16769382;
srom_1(3601) <= 16774534;
srom_1(3602) <= 16740361;
srom_1(3603) <= 16667025;
srom_1(3604) <= 16554868;
srom_1(3605) <= 16404416;
srom_1(3606) <= 16216376;
srom_1(3607) <= 15991629;
srom_1(3608) <= 15731228;
srom_1(3609) <= 15436396;
srom_1(3610) <= 15108514;
srom_1(3611) <= 14749119;
srom_1(3612) <= 14359899;
srom_1(3613) <= 13942677;
srom_1(3614) <= 13499409;
srom_1(3615) <= 13032176;
srom_1(3616) <= 12543167;
srom_1(3617) <= 12034676;
srom_1(3618) <= 11509088;
srom_1(3619) <= 10968866;
srom_1(3620) <= 10416545;
srom_1(3621) <= 9854714;
srom_1(3622) <= 9286008;
srom_1(3623) <= 8713094;
srom_1(3624) <= 8138658;
srom_1(3625) <= 7565394;
srom_1(3626) <= 6995991;
srom_1(3627) <= 6433118;
srom_1(3628) <= 5879414;
srom_1(3629) <= 5337478;
srom_1(3630) <= 4809849;
srom_1(3631) <= 4299002;
srom_1(3632) <= 3807333;
srom_1(3633) <= 3337147;
srom_1(3634) <= 2890649;
srom_1(3635) <= 2469933;
srom_1(3636) <= 2076971;
srom_1(3637) <= 1713607;
srom_1(3638) <= 1381544;
srom_1(3639) <= 1082340;
srom_1(3640) <= 817397;
srom_1(3641) <= 587959;
srom_1(3642) <= 395100;
srom_1(3643) <= 239726;
srom_1(3644) <= 122564;
srom_1(3645) <= 44165;
srom_1(3646) <= 4896;
srom_1(3647) <= 4941;
srom_1(3648) <= 44299;
srom_1(3649) <= 122787;
srom_1(3650) <= 240037;
srom_1(3651) <= 395497;
srom_1(3652) <= 588441;
srom_1(3653) <= 817962;
srom_1(3654) <= 1082984;
srom_1(3655) <= 1382265;
srom_1(3656) <= 1714400;
srom_1(3657) <= 2077834;
srom_1(3658) <= 2470861;
srom_1(3659) <= 2891638;
srom_1(3660) <= 3338193;
srom_1(3661) <= 3808430;
srom_1(3662) <= 4300146;
srom_1(3663) <= 4811034;
srom_1(3664) <= 5338698;
srom_1(3665) <= 5880665;
srom_1(3666) <= 6434391;
srom_1(3667) <= 6997282;
srom_1(3668) <= 7566698;
srom_1(3669) <= 8139967;
srom_1(3670) <= 8714403;
srom_1(3671) <= 9287311;
srom_1(3672) <= 9856004;
srom_1(3673) <= 10417816;
srom_1(3674) <= 10970113;
srom_1(3675) <= 11510304;
srom_1(3676) <= 12035856;
srom_1(3677) <= 12544305;
srom_1(3678) <= 13033267;
srom_1(3679) <= 13500448;
srom_1(3680) <= 13943658;
srom_1(3681) <= 14360819;
srom_1(3682) <= 14749973;
srom_1(3683) <= 15109298;
srom_1(3684) <= 15437106;
srom_1(3685) <= 15731862;
srom_1(3686) <= 15992182;
srom_1(3687) <= 16216847;
srom_1(3688) <= 16404803;
srom_1(3689) <= 16555167;
srom_1(3690) <= 16667236;
srom_1(3691) <= 16740484;
srom_1(3692) <= 16774567;
srom_1(3693) <= 16769325;
srom_1(3694) <= 16724783;
srom_1(3695) <= 16641150;
srom_1(3696) <= 16518818;
srom_1(3697) <= 16358360;
srom_1(3698) <= 16160530;
srom_1(3699) <= 15926254;
srom_1(3700) <= 15656632;
srom_1(3701) <= 15352928;
srom_1(3702) <= 15016565;
srom_1(3703) <= 14649122;
srom_1(3704) <= 14252321;
srom_1(3705) <= 13828023;
srom_1(3706) <= 13378217;
srom_1(3707) <= 12905014;
srom_1(3708) <= 12410632;
srom_1(3709) <= 11897389;
srom_1(3710) <= 11367692;
srom_1(3711) <= 10824025;
srom_1(3712) <= 10268938;
srom_1(3713) <= 9705033;
srom_1(3714) <= 9134955;
srom_1(3715) <= 8561377;
srom_1(3716) <= 7986989;
srom_1(3717) <= 7414484;
srom_1(3718) <= 6846548;
srom_1(3719) <= 6285842;
srom_1(3720) <= 5734997;
srom_1(3721) <= 5196596;
srom_1(3722) <= 4673163;
srom_1(3723) <= 4167153;
srom_1(3724) <= 3680939;
srom_1(3725) <= 3216801;
srom_1(3726) <= 2776915;
srom_1(3727) <= 2363345;
srom_1(3728) <= 1978029;
srom_1(3729) <= 1622774;
srom_1(3730) <= 1299247;
srom_1(3731) <= 1008964;
srom_1(3732) <= 753287;
srom_1(3733) <= 533414;
srom_1(3734) <= 350377;
srom_1(3735) <= 205034;
srom_1(3736) <= 98067;
srom_1(3737) <= 29977;
srom_1(3738) <= 1083;
srom_1(3739) <= 11522;
srom_1(3740) <= 61243;
srom_1(3741) <= 150014;
srom_1(3742) <= 277419;
srom_1(3743) <= 442860;
srom_1(3744) <= 645561;
srom_1(3745) <= 884572;
srom_1(3746) <= 1158773;
srom_1(3747) <= 1466876;
srom_1(3748) <= 1807438;
srom_1(3749) <= 2178861;
srom_1(3750) <= 2579403;
srom_1(3751) <= 3007187;
srom_1(3752) <= 3460207;
srom_1(3753) <= 3936337;
srom_1(3754) <= 4433345;
srom_1(3755) <= 4948902;
srom_1(3756) <= 5480588;
srom_1(3757) <= 6025910;
srom_1(3758) <= 6582313;
srom_1(3759) <= 7147185;
srom_1(3760) <= 7717879;
srom_1(3761) <= 8291718;
srom_1(3762) <= 8866012;
srom_1(3763) <= 9438067;
srom_1(3764) <= 10005201;
srom_1(3765) <= 10564754;
srom_1(3766) <= 11114102;
srom_1(3767) <= 11650669;
srom_1(3768) <= 12171940;
srom_1(3769) <= 12675469;
srom_1(3770) <= 13158895;
srom_1(3771) <= 13619952;
srom_1(3772) <= 14056478;
srom_1(3773) <= 14466425;
srom_1(3774) <= 14847870;
srom_1(3775) <= 15199027;
srom_1(3776) <= 15518246;
srom_1(3777) <= 15804033;
srom_1(3778) <= 16055046;
srom_1(3779) <= 16270108;
srom_1(3780) <= 16448211;
srom_1(3781) <= 16588521;
srom_1(3782) <= 16690377;
srom_1(3783) <= 16753304;
srom_1(3784) <= 16777006;
srom_1(3785) <= 16761372;
srom_1(3786) <= 16706476;
srom_1(3787) <= 16612573;
srom_1(3788) <= 16480106;
srom_1(3789) <= 16309695;
srom_1(3790) <= 16102140;
srom_1(3791) <= 15858412;
srom_1(3792) <= 15579657;
srom_1(3793) <= 15267180;
srom_1(3794) <= 14922447;
srom_1(3795) <= 14547075;
srom_1(3796) <= 14142823;
srom_1(3797) <= 13711588;
srom_1(3798) <= 13255392;
srom_1(3799) <= 12776374;
srom_1(3800) <= 12276780;
srom_1(3801) <= 11758953;
srom_1(3802) <= 11225321;
srom_1(3803) <= 10678387;
srom_1(3804) <= 10120715;
srom_1(3805) <= 9554921;
srom_1(3806) <= 8983658;
srom_1(3807) <= 8409604;
srom_1(3808) <= 7835452;
srom_1(3809) <= 7263893;
srom_1(3810) <= 6697609;
srom_1(3811) <= 6139255;
srom_1(3812) <= 5591448;
srom_1(3813) <= 5056759;
srom_1(3814) <= 4537693;
srom_1(3815) <= 4036686;
srom_1(3816) <= 3556087;
srom_1(3817) <= 3098148;
srom_1(3818) <= 2665019;
srom_1(3819) <= 2258729;
srom_1(3820) <= 1881185;
srom_1(3821) <= 1534156;
srom_1(3822) <= 1219270;
srom_1(3823) <= 938004;
srom_1(3824) <= 691675;
srom_1(3825) <= 481441;
srom_1(3826) <= 308286;
srom_1(3827) <= 173022;
srom_1(3828) <= 76284;
srom_1(3829) <= 18525;
srom_1(3830) <= 17;
srom_1(3831) <= 20845;
srom_1(3832) <= 80913;
srom_1(3833) <= 179938;
srom_1(3834) <= 317457;
srom_1(3835) <= 492824;
srom_1(3836) <= 705217;
srom_1(3837) <= 953640;
srom_1(3838) <= 1236928;
srom_1(3839) <= 1553753;
srom_1(3840) <= 1902629;
srom_1(3841) <= 2281920;
srom_1(3842) <= 2689847;
srom_1(3843) <= 3124498;
srom_1(3844) <= 3583834;
srom_1(3845) <= 4065701;
srom_1(3846) <= 4567840;
srom_1(3847) <= 5087895;
srom_1(3848) <= 5623429;
srom_1(3849) <= 6171930;
srom_1(3850) <= 6730825;
srom_1(3851) <= 7297494;
srom_1(3852) <= 7869280;
srom_1(3853) <= 8443501;
srom_1(3854) <= 9017465;
srom_1(3855) <= 9588480;
srom_1(3856) <= 10153868;
srom_1(3857) <= 10710978;
srom_1(3858) <= 11257198;
srom_1(3859) <= 11789966;
srom_1(3860) <= 12306784;
srom_1(3861) <= 12805229;
srom_1(3862) <= 13282962;
srom_1(3863) <= 13737744;
srom_1(3864) <= 14167442;
srom_1(3865) <= 14570041;
srom_1(3866) <= 14943653;
srom_1(3867) <= 15286526;
srom_1(3868) <= 15597053;
srom_1(3869) <= 15873776;
srom_1(3870) <= 16115399;
srom_1(3871) <= 16320789;
srom_1(3872) <= 16488982;
srom_1(3873) <= 16619189;
srom_1(3874) <= 16710801;
srom_1(3875) <= 16763386;
srom_1(3876) <= 16776700;
srom_1(3877) <= 16750679;
srom_1(3878) <= 16685445;
srom_1(3879) <= 16581304;
srom_1(3880) <= 16438745;
srom_1(3881) <= 16258437;
srom_1(3882) <= 16041224;
srom_1(3883) <= 15788125;
srom_1(3884) <= 15500327;
srom_1(3885) <= 15179180;
srom_1(3886) <= 14826190;
srom_1(3887) <= 14443011;
srom_1(3888) <= 14031442;
srom_1(3889) <= 13593411;
srom_1(3890) <= 13130973;
srom_1(3891) <= 12646297;
srom_1(3892) <= 12141654;
srom_1(3893) <= 11619413;
srom_1(3894) <= 11082021;
srom_1(3895) <= 10531999;
srom_1(3896) <= 9971925;
srom_1(3897) <= 9404427;
srom_1(3898) <= 8832165;
srom_1(3899) <= 8257824;
srom_1(3900) <= 7684095;
srom_1(3901) <= 7113671;
srom_1(3902) <= 6549225;
srom_1(3903) <= 5993404;
srom_1(3904) <= 5448816;
srom_1(3905) <= 4918013;
srom_1(3906) <= 4403485;
srom_1(3907) <= 3907644;
srom_1(3908) <= 3432816;
srom_1(3909) <= 2981228;
srom_1(3910) <= 2554997;
srom_1(3911) <= 2156121;
srom_1(3912) <= 1786472;
srom_1(3913) <= 1447782;
srom_1(3914) <= 1141641;
srom_1(3915) <= 869483;
srom_1(3916) <= 632584;
srom_1(3917) <= 432056;
srom_1(3918) <= 268840;
srom_1(3919) <= 143699;
srom_1(3920) <= 57222;
srom_1(3921) <= 9814;
srom_1(3922) <= 1696;
srom_1(3923) <= 32908;
srom_1(3924) <= 103303;
srom_1(3925) <= 212550;
srom_1(3926) <= 360137;
srom_1(3927) <= 545373;
srom_1(3928) <= 767388;
srom_1(3929) <= 1025142;
srom_1(3930) <= 1317426;
srom_1(3931) <= 1642868;
srom_1(3932) <= 1999944;
srom_1(3933) <= 2386979;
srom_1(3934) <= 2802157;
srom_1(3935) <= 3243532;
srom_1(3936) <= 3709034;
srom_1(3937) <= 4196480;
srom_1(3938) <= 4703585;
srom_1(3939) <= 5227970;
srom_1(3940) <= 5767176;
srom_1(3941) <= 6318675;
srom_1(3942) <= 6879880;
srom_1(3943) <= 7448161;
srom_1(3944) <= 8020851;
srom_1(3945) <= 8595266;
srom_1(3946) <= 9168712;
srom_1(3947) <= 9738500;
srom_1(3948) <= 10301958;
srom_1(3949) <= 10856443;
srom_1(3950) <= 11399356;
srom_1(3951) <= 11928150;
srom_1(3952) <= 12440346;
srom_1(3953) <= 12933543;
srom_1(3954) <= 13405426;
srom_1(3955) <= 13853784;
srom_1(3956) <= 14276514;
srom_1(3957) <= 14671633;
srom_1(3958) <= 15037289;
srom_1(3959) <= 15371767;
srom_1(3960) <= 15673499;
srom_1(3961) <= 15941069;
srom_1(3962) <= 16173223;
srom_1(3963) <= 16368873;
srom_1(3964) <= 16527100;
srom_1(3965) <= 16647163;
srom_1(3966) <= 16728499;
srom_1(3967) <= 16770726;
srom_1(3968) <= 16773647;
srom_1(3969) <= 16737247;
srom_1(3970) <= 16661698;
srom_1(3971) <= 16547353;
srom_1(3972) <= 16394749;
srom_1(3973) <= 16204602;
srom_1(3974) <= 15977802;
srom_1(3975) <= 15715415;
srom_1(3976) <= 15418669;
srom_1(3977) <= 15088957;
srom_1(3978) <= 14727825;
srom_1(3979) <= 14336966;
srom_1(3980) <= 13918213;
srom_1(3981) <= 13473530;
srom_1(3982) <= 13005002;
srom_1(3983) <= 12514826;
srom_1(3984) <= 12005300;
srom_1(3985) <= 11478815;
srom_1(3986) <= 10937839;
srom_1(3987) <= 10384909;
srom_1(3988) <= 9822617;
srom_1(3989) <= 9253601;
srom_1(3990) <= 8680528;
srom_1(3991) <= 8106087;
srom_1(3992) <= 7532970;
srom_1(3993) <= 6963866;
srom_1(3994) <= 6401442;
srom_1(3995) <= 5848338;
srom_1(3996) <= 5307145;
srom_1(3997) <= 4780403;
srom_1(3998) <= 4270580;
srom_1(3999) <= 3780069;
srom_1(4000) <= 3311168;
srom_1(4001) <= 2866078;
srom_1(4002) <= 2446884;
srom_1(4003) <= 2055553;
srom_1(4004) <= 1693920;
srom_1(4005) <= 1363681;
srom_1(4006) <= 1066384;
srom_1(4007) <= 803423;
srom_1(4008) <= 576032;
srom_1(4009) <= 385277;
srom_1(4010) <= 232052;
srom_1(4011) <= 117076;
srom_1(4012) <= 40888;
srom_1(4013) <= 3846;
srom_1(4014) <= 6122;
srom_1(4015) <= 47707;
srom_1(4016) <= 128405;
srom_1(4017) <= 247838;
srom_1(4018) <= 405446;
srom_1(4019) <= 600490;
srom_1(4020) <= 832054;
srom_1(4021) <= 1099055;
srom_1(4022) <= 1400238;
srom_1(4023) <= 1734192;
srom_1(4024) <= 2099351;
srom_1(4025) <= 2494003;
srom_1(4026) <= 2916296;
srom_1(4027) <= 3364251;
srom_1(4028) <= 3835767;
srom_1(4029) <= 4328632;
srom_1(4030) <= 4840536;
srom_1(4031) <= 5369079;
srom_1(4032) <= 5911781;
srom_1(4033) <= 6466097;
srom_1(4034) <= 7029429;
srom_1(4035) <= 7599135;
srom_1(4036) <= 8172543;
srom_1(4037) <= 8746964;
srom_1(4038) <= 9319704;
srom_1(4039) <= 9888078;
srom_1(4040) <= 10449421;
srom_1(4041) <= 11001100;
srom_1(4042) <= 11540528;
srom_1(4043) <= 12065175;
srom_1(4044) <= 12572582;
srom_1(4045) <= 13060369;
srom_1(4046) <= 13526248;
srom_1(4047) <= 13968035;
srom_1(4048) <= 14383658;
srom_1(4049) <= 14771168;
srom_1(4050) <= 15128749;
srom_1(4051) <= 15454722;
srom_1(4052) <= 15747560;
srom_1(4053) <= 16005889;
srom_1(4054) <= 16228499;
srom_1(4055) <= 16414344;
srom_1(4056) <= 16562554;
srom_1(4057) <= 16672433;
srom_1(4058) <= 16743467;
srom_1(4059) <= 16775322;
srom_1(4060) <= 16767849;
srom_1(4061) <= 16721082;
srom_1(4062) <= 16635242;
srom_1(4063) <= 16510731;
srom_1(4064) <= 16348132;
srom_1(4065) <= 16148208;
srom_1(4066) <= 15911896;
srom_1(4067) <= 15640306;
srom_1(4068) <= 15334709;
srom_1(4069) <= 14996540;
srom_1(4070) <= 14627384;
srom_1(4071) <= 14228973;
srom_1(4072) <= 13803174;
srom_1(4073) <= 13351984;
srom_1(4074) <= 12877519;
srom_1(4075) <= 12382004;
srom_1(4076) <= 11867762;
srom_1(4077) <= 11337206;
srom_1(4078) <= 10792823;
srom_1(4079) <= 10237165;
srom_1(4080) <= 9672839;
srom_1(4081) <= 9102491;
srom_1(4082) <= 8528795;
srom_1(4083) <= 7954442;
srom_1(4084) <= 7382124;
srom_1(4085) <= 6814527;
srom_1(4086) <= 6254311;
srom_1(4087) <= 5704103;
srom_1(4088) <= 5166484;
srom_1(4089) <= 4643974;
srom_1(4090) <= 4139024;
srom_1(4091) <= 3654002;
srom_1(4092) <= 3191183;
srom_1(4093) <= 2752735;
srom_1(4094) <= 2340717;
srom_1(4095) <= 1957059;
srom_1(4096) <= 1603560;
srom_1(4097) <= 1281879;
srom_1(4098) <= 993524;
srom_1(4099) <= 739847;
srom_1(4100) <= 522038;
srom_1(4101) <= 341118;
srom_1(4102) <= 197935;
srom_1(4103) <= 93161;
srom_1(4104) <= 27287;
srom_1(4105) <= 623;
srom_1(4106) <= 13292;
srom_1(4107) <= 65236;
srom_1(4108) <= 156212;
srom_1(4109) <= 285792;
srom_1(4110) <= 453368;
srom_1(4111) <= 658156;
srom_1(4112) <= 899195;
srom_1(4113) <= 1175354;
srom_1(4114) <= 1485338;
srom_1(4115) <= 1827694;
srom_1(4116) <= 2200817;
srom_1(4117) <= 2602956;
srom_1(4118) <= 3032226;
srom_1(4119) <= 3486614;
srom_1(4120) <= 3963989;
srom_1(4121) <= 4462113;
srom_1(4122) <= 4978650;
srom_1(4123) <= 5511176;
srom_1(4124) <= 6057197;
srom_1(4125) <= 6614150;
srom_1(4126) <= 7179423;
srom_1(4127) <= 7750368;
srom_1(4128) <= 8324305;
srom_1(4129) <= 8898543;
srom_1(4130) <= 9470391;
srom_1(4131) <= 10037165;
srom_1(4132) <= 10596209;
srom_1(4133) <= 11144901;
srom_1(4134) <= 11680667;
srom_1(4135) <= 12200996;
srom_1(4136) <= 12703448;
srom_1(4137) <= 13185665;
srom_1(4138) <= 13645387;
srom_1(4139) <= 14080459;
srom_1(4140) <= 14488840;
srom_1(4141) <= 14868614;
srom_1(4142) <= 15218001;
srom_1(4143) <= 15535364;
srom_1(4144) <= 15819212;
srom_1(4145) <= 16068216;
srom_1(4146) <= 16281207;
srom_1(4147) <= 16457188;
srom_1(4148) <= 16595332;
srom_1(4149) <= 16694992;
srom_1(4150) <= 16755700;
srom_1(4151) <= 16777172;
srom_1(4152) <= 16759307;
srom_1(4153) <= 16702190;
srom_1(4154) <= 16606087;
srom_1(4155) <= 16471449;
srom_1(4156) <= 16298908;
srom_1(4157) <= 16089273;
srom_1(4158) <= 15843527;
srom_1(4159) <= 15562823;
srom_1(4160) <= 15248476;
srom_1(4161) <= 14901960;
srom_1(4162) <= 14524901;
srom_1(4163) <= 14119068;
srom_1(4164) <= 13686362;
srom_1(4165) <= 13228813;
srom_1(4166) <= 12748566;
srom_1(4167) <= 12247874;
srom_1(4168) <= 11729085;
srom_1(4169) <= 11194631;
srom_1(4170) <= 10647019;
srom_1(4171) <= 10088817;
srom_1(4172) <= 9522641;
srom_1(4173) <= 8951148;
srom_1(4174) <= 8377016;
srom_1(4175) <= 7802939;
srom_1(4176) <= 7231608;
srom_1(4177) <= 6665703;
srom_1(4178) <= 6107878;
srom_1(4179) <= 5560747;
srom_1(4180) <= 5026877;
srom_1(4181) <= 4508771;
srom_1(4182) <= 4008860;
srom_1(4183) <= 3529486;
srom_1(4184) <= 3072899;
srom_1(4185) <= 2641238;
srom_1(4186) <= 2236529;
srom_1(4187) <= 1860670;
srom_1(4188) <= 1515422;
srom_1(4189) <= 1202405;
srom_1(4190) <= 923086;
srom_1(4191) <= 678776;
srom_1(4192) <= 470619;
srom_1(4193) <= 299593;
srom_1(4194) <= 166499;
srom_1(4195) <= 71962;
srom_1(4196) <= 16424;
srom_1(4197) <= 146;
srom_1(4198) <= 23204;
srom_1(4199) <= 85491;
srom_1(4200) <= 186714;
srom_1(4201) <= 326398;
srom_1(4202) <= 503889;
srom_1(4203) <= 718354;
srom_1(4204) <= 968787;
srom_1(4205) <= 1254014;
srom_1(4206) <= 1572698;
srom_1(4207) <= 1923345;
srom_1(4208) <= 2304308;
srom_1(4209) <= 2713804;
srom_1(4210) <= 3149910;
srom_1(4211) <= 3610583;
srom_1(4212) <= 4093661;
srom_1(4213) <= 4596880;
srom_1(4214) <= 5117879;
srom_1(4215) <= 5654216;
srom_1(4216) <= 6203376;
srom_1(4217) <= 6762783;
srom_1(4218) <= 7329813;
srom_1(4219) <= 7901809;
srom_1(4220) <= 8476088;
srom_1(4221) <= 9049956;
srom_1(4222) <= 9620724;
srom_1(4223) <= 10185713;
srom_1(4224) <= 10742275;
srom_1(4225) <= 11287800;
srom_1(4226) <= 11819729;
srom_1(4227) <= 12335569;
srom_1(4228) <= 12832901;
srom_1(4229) <= 13309391;
srom_1(4230) <= 13762806;
srom_1(4231) <= 14191020;
srom_1(4232) <= 14592024;
srom_1(4233) <= 14963938;
srom_1(4234) <= 15305018;
srom_1(4235) <= 15613665;
srom_1(4236) <= 15888431;
srom_1(4237) <= 16128028;
srom_1(4238) <= 16331332;
srom_1(4239) <= 16497390;
srom_1(4240) <= 16625423;
srom_1(4241) <= 16714830;
srom_1(4242) <= 16765193;
srom_1(4243) <= 16776276;
srom_1(4244) <= 16748026;
srom_1(4245) <= 16680575;
srom_1(4246) <= 16574241;
srom_1(4247) <= 16429521;
srom_1(4248) <= 16247095;
srom_1(4249) <= 16027818;
srom_1(4250) <= 15772718;
srom_1(4251) <= 15482991;
srom_1(4252) <= 15159996;
srom_1(4253) <= 14805248;
srom_1(4254) <= 14420410;
srom_1(4255) <= 14007286;
srom_1(4256) <= 13567815;
srom_1(4257) <= 13104057;
srom_1(4258) <= 12618186;
srom_1(4259) <= 12112482;
srom_1(4260) <= 11589315;
srom_1(4261) <= 11051138;
srom_1(4262) <= 10500476;
srom_1(4263) <= 9939911;
srom_1(4264) <= 9372071;
srom_1(4265) <= 8799620;
srom_1(4266) <= 8225241;
srom_1(4267) <= 7651628;
srom_1(4268) <= 7081471;
srom_1(4269) <= 6517444;
srom_1(4270) <= 5962191;
srom_1(4271) <= 5418317;
srom_1(4272) <= 4888371;
srom_1(4273) <= 4374839;
srom_1(4274) <= 3880129;
srom_1(4275) <= 3406561;
srom_1(4276) <= 2956355;
srom_1(4277) <= 2531623;
srom_1(4278) <= 2134356;
srom_1(4279) <= 1766418;
srom_1(4280) <= 1429534;
srom_1(4281) <= 1125282;
srom_1(4282) <= 855092;
srom_1(4283) <= 620228;
srom_1(4284) <= 421793;
srom_1(4285) <= 260717;
srom_1(4286) <= 137756;
srom_1(4287) <= 53485;
srom_1(4288) <= 8301;
srom_1(4289) <= 2415;
srom_1(4290) <= 35855;
srom_1(4291) <= 108464;
srom_1(4292) <= 219901;
srom_1(4293) <= 369644;
srom_1(4294) <= 556990;
srom_1(4295) <= 781062;
srom_1(4296) <= 1040808;
srom_1(4297) <= 1335011;
srom_1(4298) <= 1662290;
srom_1(4299) <= 2021111;
srom_1(4300) <= 2409792;
srom_1(4301) <= 2826509;
srom_1(4302) <= 3269309;
srom_1(4303) <= 3736115;
srom_1(4304) <= 4224739;
srom_1(4305) <= 4732888;
srom_1(4306) <= 5258180;
srom_1(4307) <= 5798151;
srom_1(4308) <= 6350270;
srom_1(4309) <= 6911948;
srom_1(4310) <= 7480550;
srom_1(4311) <= 8053410;
srom_1(4312) <= 8627843;
srom_1(4313) <= 9201153;
srom_1(4314) <= 9770653;
srom_1(4315) <= 10333672;
srom_1(4316) <= 10887570;
srom_1(4317) <= 11429750;
srom_1(4318) <= 11957668;
srom_1(4319) <= 12468850;
srom_1(4320) <= 12960899;
srom_1(4321) <= 13431506;
srom_1(4322) <= 13878465;
srom_1(4323) <= 14299681;
srom_1(4324) <= 14693177;
srom_1(4325) <= 15057110;
srom_1(4326) <= 15389771;
srom_1(4327) <= 15689601;
srom_1(4328) <= 15955195;
srom_1(4329) <= 16185306;
srom_1(4330) <= 16378856;
srom_1(4331) <= 16534937;
srom_1(4332) <= 16652817;
srom_1(4333) <= 16731943;
srom_1(4334) <= 16771944;
srom_1(4335) <= 16772633;
srom_1(4336) <= 16734007;
srom_1(4337) <= 16656246;
srom_1(4338) <= 16539715;
srom_1(4339) <= 16384961;
srom_1(4340) <= 16192709;
srom_1(4341) <= 15963861;
srom_1(4342) <= 15699490;
srom_1(4343) <= 15400836;
srom_1(4344) <= 15069299;
srom_1(4345) <= 14706434;
srom_1(4346) <= 14313943;
srom_1(4347) <= 13893666;
srom_1(4348) <= 13447573;
srom_1(4349) <= 12977757;
srom_1(4350) <= 12486422;
srom_1(4351) <= 11975870;
srom_1(4352) <= 11448496;
srom_1(4353) <= 10906773;
srom_1(4354) <= 10353242;
srom_1(4355) <= 9790498;
srom_1(4356) <= 9221180;
srom_1(4357) <= 8647958;
srom_1(4358) <= 8073519;
srom_1(4359) <= 7500559;
srom_1(4360) <= 6931762;
srom_1(4361) <= 6369797;
srom_1(4362) <= 5817299;
srom_1(4363) <= 5276859;
srom_1(4364) <= 4751011;
srom_1(4365) <= 4242221;
srom_1(4366) <= 3752874;
srom_1(4367) <= 3285266;
srom_1(4368) <= 2841590;
srom_1(4369) <= 2423925;
srom_1(4370) <= 2034231;
srom_1(4371) <= 1674334;
srom_1(4372) <= 1345924;
srom_1(4373) <= 1050538;
srom_1(4374) <= 789564;
srom_1(4375) <= 564224;
srom_1(4376) <= 375575;
srom_1(4377) <= 224502;
srom_1(4378) <= 111713;
srom_1(4379) <= 37738;
srom_1(4380) <= 2922;
srom_1(4381) <= 7430;
srom_1(4382) <= 51240;
srom_1(4383) <= 134147;
srom_1(4384) <= 255762;
srom_1(4385) <= 415515;
srom_1(4386) <= 612656;
srom_1(4387) <= 846261;
srom_1(4388) <= 1115235;
srom_1(4389) <= 1418317;
srom_1(4390) <= 1754084;
srom_1(4391) <= 2120963;
srom_1(4392) <= 2517233;
srom_1(4393) <= 2941036;
srom_1(4394) <= 3390384;
srom_1(4395) <= 3863171;
srom_1(4396) <= 4357180;
srom_1(4397) <= 4870092;
srom_1(4398) <= 5399505;
srom_1(4399) <= 5942934;
srom_1(4400) <= 6497832;
srom_1(4401) <= 7061597;
srom_1(4402) <= 7631584;
srom_1(4403) <= 8205121;
srom_1(4404) <= 8779519;
srom_1(4405) <= 9352083;
srom_1(4406) <= 9920130;
srom_1(4407) <= 10480994;
srom_1(4408) <= 11032047;
srom_1(4409) <= 11570704;
srom_1(4410) <= 12094438;
srom_1(4411) <= 12600795;
srom_1(4412) <= 13087400;
srom_1(4413) <= 13551970;
srom_1(4414) <= 13992327;
srom_1(4415) <= 14406407;
srom_1(4416) <= 14792267;
srom_1(4417) <= 15148098;
srom_1(4418) <= 15472231;
srom_1(4419) <= 15763147;
srom_1(4420) <= 16019482;
srom_1(4421) <= 16240032;
srom_1(4422) <= 16423764;
srom_1(4423) <= 16569817;
srom_1(4424) <= 16677505;
srom_1(4425) <= 16746324;
srom_1(4426) <= 16775951;
srom_1(4427) <= 16766246;
srom_1(4428) <= 16717256;
srom_1(4429) <= 16629210;
srom_1(4430) <= 16502521;
srom_1(4431) <= 16337783;
srom_1(4432) <= 16135768;
srom_1(4433) <= 15897425;
srom_1(4434) <= 15623870;
srom_1(4435) <= 15316386;
srom_1(4436) <= 14976416;
srom_1(4437) <= 14605553;
srom_1(4438) <= 14205536;
srom_1(4439) <= 13778243;
srom_1(4440) <= 13325675;
srom_1(4441) <= 12849955;
srom_1(4442) <= 12353315;
srom_1(4443) <= 11838083;
srom_1(4444) <= 11306676;
srom_1(4445) <= 10761584;
srom_1(4446) <= 10205365;
srom_1(4447) <= 9640626;
srom_1(4448) <= 9070016;
srom_1(4449) <= 8496211;
srom_1(4450) <= 7921901;
srom_1(4451) <= 7349780;
srom_1(4452) <= 6782530;
srom_1(4453) <= 6222811;
srom_1(4454) <= 5673249;
srom_1(4455) <= 5136420;
srom_1(4456) <= 4614842;
srom_1(4457) <= 4110960;
srom_1(4458) <= 3627137;
srom_1(4459) <= 3165643;
srom_1(4460) <= 2728641;
srom_1(4461) <= 2318180;
srom_1(4462) <= 1936186;
srom_1(4463) <= 1584449;
srom_1(4464) <= 1264619;
srom_1(4465) <= 978197;
srom_1(4466) <= 726524;
srom_1(4467) <= 510781;
srom_1(4468) <= 331980;
srom_1(4469) <= 190959;
srom_1(4470) <= 88380;
srom_1(4471) <= 24724;
srom_1(4472) <= 289;
srom_1(4473) <= 15189;
srom_1(4474) <= 69355;
srom_1(4475) <= 162533;
srom_1(4476) <= 294286;
srom_1(4477) <= 463996;
srom_1(4478) <= 670868;
srom_1(4479) <= 913930;
srom_1(4480) <= 1192044;
srom_1(4481) <= 1503904;
srom_1(4482) <= 1848050;
srom_1(4483) <= 2222867;
srom_1(4484) <= 2626596;
srom_1(4485) <= 3057346;
srom_1(4486) <= 3513096;
srom_1(4487) <= 3991709;
srom_1(4488) <= 4490940;
srom_1(4489) <= 5008449;
srom_1(4490) <= 5541809;
srom_1(4491) <= 6088518;
srom_1(4492) <= 6646013;
srom_1(4493) <= 7211680;
srom_1(4494) <= 7782866;
srom_1(4495) <= 8356892;
srom_1(4496) <= 8931067;
srom_1(4497) <= 9502698;
srom_1(4498) <= 10069105;
srom_1(4499) <= 10627632;
srom_1(4500) <= 11175659;
srom_1(4501) <= 11710616;
srom_1(4502) <= 12229995;
srom_1(4503) <= 12731361;
srom_1(4504) <= 13212362;
srom_1(4505) <= 13670743;
srom_1(4506) <= 14104354;
srom_1(4507) <= 14511162;
srom_1(4508) <= 14889260;
srom_1(4509) <= 15236873;
srom_1(4510) <= 15552373;
srom_1(4511) <= 15834279;
srom_1(4512) <= 16081270;
srom_1(4513) <= 16292187;
srom_1(4514) <= 16466042;
srom_1(4515) <= 16602019;
srom_1(4516) <= 16699480;
srom_1(4517) <= 16757969;
srom_1(4518) <= 16777211;
srom_1(4519) <= 16757116;
srom_1(4520) <= 16697778;
srom_1(4521) <= 16599476;
srom_1(4522) <= 16462670;
srom_1(4523) <= 16288002;
srom_1(4524) <= 16076291;
srom_1(4525) <= 15828530;
srom_1(4526) <= 15545880;
srom_1(4527) <= 15229668;
srom_1(4528) <= 14881375;
srom_1(4529) <= 14502636;
srom_1(4530) <= 14095225;
srom_1(4531) <= 13661055;
srom_1(4532) <= 13202160;
srom_1(4533) <= 12720693;
srom_1(4534) <= 12218911;
srom_1(4535) <= 11699168;
srom_1(4536) <= 11163900;
srom_1(4537) <= 10615618;
srom_1(4538) <= 10056892;
srom_1(4539) <= 9490344;
srom_1(4540) <= 8918629;
srom_1(4541) <= 8344428;
srom_1(4542) <= 7770435;
srom_1(4543) <= 7199341;
srom_1(4544) <= 6633823;
srom_1(4545) <= 6076535;
srom_1(4546) <= 5530088;
srom_1(4547) <= 4997046;
srom_1(4548) <= 4479908;
srom_1(4549) <= 3981099;
srom_1(4550) <= 3502959;
srom_1(4551) <= 3047729;
srom_1(4552) <= 2617544;
srom_1(4553) <= 2214422;
srom_1(4554) <= 1840253;
srom_1(4555) <= 1496791;
srom_1(4556) <= 1185647;
srom_1(4557) <= 908281;
srom_1(4558) <= 665992;
srom_1(4559) <= 459917;
srom_1(4560) <= 291023;
srom_1(4561) <= 160101;
srom_1(4562) <= 67765;
srom_1(4563) <= 14449;
srom_1(4564) <= 401;
srom_1(4565) <= 25689;
srom_1(4566) <= 90194;
srom_1(4567) <= 193613;
srom_1(4568) <= 335461;
srom_1(4569) <= 515072;
srom_1(4570) <= 731606;
srom_1(4571) <= 984046;
srom_1(4572) <= 1271208;
srom_1(4573) <= 1591746;
srom_1(4574) <= 1944157;
srom_1(4575) <= 2326789;
srom_1(4576) <= 2737846;
srom_1(4577) <= 3175402;
srom_1(4578) <= 3637404;
srom_1(4579) <= 4121686;
srom_1(4580) <= 4625977;
srom_1(4581) <= 5147913;
srom_1(4582) <= 5685045;
srom_1(4583) <= 6234855;
srom_1(4584) <= 6794765;
srom_1(4585) <= 7362149;
srom_1(4586) <= 7934346;
srom_1(4587) <= 8508673;
srom_1(4588) <= 9082438;
srom_1(4589) <= 9652949;
srom_1(4590) <= 10217531;
srom_1(4591) <= 10773536;
srom_1(4592) <= 11318358;
srom_1(4593) <= 11849441;
srom_1(4594) <= 12364295;
srom_1(4595) <= 12860505;
srom_1(4596) <= 13335746;
srom_1(4597) <= 13787787;
srom_1(4598) <= 14214510;
srom_1(4599) <= 14613914;
srom_1(4600) <= 14984124;
srom_1(4601) <= 15323406;
srom_1(4602) <= 15630169;
srom_1(4603) <= 15902973;
srom_1(4604) <= 16140540;
srom_1(4605) <= 16341755;
srom_1(4606) <= 16505675;
srom_1(4607) <= 16631532;
srom_1(4608) <= 16718734;
srom_1(4609) <= 16766874;
srom_1(4610) <= 16775725;
srom_1(4611) <= 16745246;
srom_1(4612) <= 16675580;
srom_1(4613) <= 16567054;
srom_1(4614) <= 16420176;
srom_1(4615) <= 16235635;
srom_1(4616) <= 16014297;
srom_1(4617) <= 15757199;
srom_1(4618) <= 15465547;
srom_1(4619) <= 15140709;
srom_1(4620) <= 14784209;
srom_1(4621) <= 14397717;
srom_1(4622) <= 13983046;
srom_1(4623) <= 13542141;
srom_1(4624) <= 13077070;
srom_1(4625) <= 12590012;
srom_1(4626) <= 12083253;
srom_1(4627) <= 11559168;
srom_1(4628) <= 11020215;
srom_1(4629) <= 10468922;
srom_1(4630) <= 9907874;
srom_1(4631) <= 9339701;
srom_1(4632) <= 8767068;
srom_1(4633) <= 8192661;
srom_1(4634) <= 7619172;
srom_1(4635) <= 7049291;
srom_1(4636) <= 6485691;
srom_1(4637) <= 5931015;
srom_1(4638) <= 5387863;
srom_1(4639) <= 4858782;
srom_1(4640) <= 4346254;
srom_1(4641) <= 3852682;
srom_1(4642) <= 3380380;
srom_1(4643) <= 2931564;
srom_1(4644) <= 2508338;
srom_1(4645) <= 2112686;
srom_1(4646) <= 1746464;
srom_1(4647) <= 1411390;
srom_1(4648) <= 1109034;
srom_1(4649) <= 840814;
srom_1(4650) <= 607989;
srom_1(4651) <= 411650;
srom_1(4652) <= 252717;
srom_1(4653) <= 131936;
srom_1(4654) <= 49874;
srom_1(4655) <= 6915;
srom_1(4656) <= 3260;
srom_1(4657) <= 38928;
srom_1(4658) <= 113750;
srom_1(4659) <= 227375;
srom_1(4660) <= 379271;
srom_1(4661) <= 568726;
srom_1(4662) <= 794851;
srom_1(4663) <= 1056586;
srom_1(4664) <= 1352703;
srom_1(4665) <= 1681813;
srom_1(4666) <= 2042375;
srom_1(4667) <= 2432695;
srom_1(4668) <= 2850946;
srom_1(4669) <= 3295164;
srom_1(4670) <= 3763267;
srom_1(4671) <= 4253060;
srom_1(4672) <= 4762246;
srom_1(4673) <= 5288437;
srom_1(4674) <= 5829166;
srom_1(4675) <= 6381897;
srom_1(4676) <= 6944038;
srom_1(4677) <= 7512953;
srom_1(4678) <= 8085975;
srom_1(4679) <= 8660415;
srom_1(4680) <= 9233581;
srom_1(4681) <= 9802785;
srom_1(4682) <= 10365357;
srom_1(4683) <= 10918659;
srom_1(4684) <= 11460098;
srom_1(4685) <= 11987132;
srom_1(4686) <= 12497292;
srom_1(4687) <= 12988186;
srom_1(4688) <= 13457510;
srom_1(4689) <= 13903064;
srom_1(4690) <= 14322759;
srom_1(4691) <= 14714627;
srom_1(4692) <= 15076830;
srom_1(4693) <= 15407669;
srom_1(4694) <= 15705594;
srom_1(4695) <= 15969207;
srom_1(4696) <= 16197272;
srom_1(4697) <= 16388719;
srom_1(4698) <= 16542651;
srom_1(4699) <= 16658346;
srom_1(4700) <= 16735261;
srom_1(4701) <= 16773036;
srom_1(4702) <= 16771493;
srom_1(4703) <= 16730641;
srom_1(4704) <= 16650669;
srom_1(4705) <= 16531954;
srom_1(4706) <= 16375052;
srom_1(4707) <= 16180699;
srom_1(4708) <= 15949806;
srom_1(4709) <= 15683456;
srom_1(4710) <= 15382898;
srom_1(4711) <= 15049541;
srom_1(4712) <= 14684949;
srom_1(4713) <= 14290831;
srom_1(4714) <= 13869035;
srom_1(4715) <= 13421540;
srom_1(4716) <= 12950444;
srom_1(4717) <= 12457956;
srom_1(4718) <= 11946385;
srom_1(4719) <= 11418130;
srom_1(4720) <= 10875670;
srom_1(4721) <= 10321546;
srom_1(4722) <= 9758358;
srom_1(4723) <= 9188747;
srom_1(4724) <= 8615384;
srom_1(4725) <= 8040957;
srom_1(4726) <= 7468161;
srom_1(4727) <= 6899680;
srom_1(4728) <= 6338182;
srom_1(4729) <= 5786300;
srom_1(4730) <= 5246620;
srom_1(4731) <= 4721674;
srom_1(4732) <= 4213923;
srom_1(4733) <= 3725749;
srom_1(4734) <= 3259441;
srom_1(4735) <= 2817186;
srom_1(4736) <= 2401056;
srom_1(4737) <= 2013004;
srom_1(4738) <= 1654850;
srom_1(4739) <= 1328273;
srom_1(4740) <= 1034803;
srom_1(4741) <= 775819;
srom_1(4742) <= 552533;
srom_1(4743) <= 365994;
srom_1(4744) <= 217075;
srom_1(4745) <= 106475;
srom_1(4746) <= 34713;
srom_1(4747) <= 2125;
srom_1(4748) <= 8865;
srom_1(4749) <= 54900;
srom_1(4750) <= 140014;
srom_1(4751) <= 263809;
srom_1(4752) <= 425704;
srom_1(4753) <= 624940;
srom_1(4754) <= 860582;
srom_1(4755) <= 1131526;
srom_1(4756) <= 1436501;
srom_1(4757) <= 1774076;
srom_1(4758) <= 2142669;
srom_1(4759) <= 2540552;
srom_1(4760) <= 2965858;
srom_1(4761) <= 3416594;
srom_1(4762) <= 3890644;
srom_1(4763) <= 4385788;
srom_1(4764) <= 4899702;
srom_1(4765) <= 5429976;
srom_1(4766) <= 5974125;
srom_1(4767) <= 6529596;
srom_1(4768) <= 7093784;
srom_1(4769) <= 7664044;
srom_1(4770) <= 8237703;
srom_1(4771) <= 8812068;
srom_1(4772) <= 9384448;
srom_1(4773) <= 9952158;
srom_1(4774) <= 10512536;
srom_1(4775) <= 11062955;
srom_1(4776) <= 11600832;
srom_1(4777) <= 12123646;
srom_1(4778) <= 12628945;
srom_1(4779) <= 13114360;
srom_1(4780) <= 13577614;
srom_1(4781) <= 14016535;
srom_1(4782) <= 14429065;
srom_1(4783) <= 14813269;
srom_1(4784) <= 15167345;
srom_1(4785) <= 15489634;
srom_1(4786) <= 15778623;
srom_1(4787) <= 16032959;
srom_1(4788) <= 16251447;
srom_1(4789) <= 16433064;
srom_1(4790) <= 16576957;
srom_1(4791) <= 16682452;
srom_1(4792) <= 16749055;
srom_1(4793) <= 16776453;
srom_1(4794) <= 16764517;
srom_1(4795) <= 16713304;
srom_1(4796) <= 16623053;
srom_1(4797) <= 16494188;
srom_1(4798) <= 16327314;
srom_1(4799) <= 16123212;
srom_1(4800) <= 15882840;
srom_1(4801) <= 15607324;
srom_1(4802) <= 15297958;
srom_1(4803) <= 14956191;
srom_1(4804) <= 14583627;
srom_1(4805) <= 14182012;
srom_1(4806) <= 13753230;
srom_1(4807) <= 13299291;
srom_1(4808) <= 12822325;
srom_1(4809) <= 12324567;
srom_1(4810) <= 11808352;
srom_1(4811) <= 11276101;
srom_1(4812) <= 10730309;
srom_1(4813) <= 10173537;
srom_1(4814) <= 9608394;
srom_1(4815) <= 9037531;
srom_1(4816) <= 8463625;
srom_1(4817) <= 7889367;
srom_1(4818) <= 7317451;
srom_1(4819) <= 6750557;
srom_1(4820) <= 6191345;
srom_1(4821) <= 5642436;
srom_1(4822) <= 5106406;
srom_1(4823) <= 4585766;
srom_1(4824) <= 4082960;
srom_1(4825) <= 3600344;
srom_1(4826) <= 3140182;
srom_1(4827) <= 2704631;
srom_1(4828) <= 2295735;
srom_1(4829) <= 1915410;
srom_1(4830) <= 1565440;
srom_1(4831) <= 1247467;
srom_1(4832) <= 962981;
srom_1(4833) <= 713316;
srom_1(4834) <= 499643;
srom_1(4835) <= 322964;
srom_1(4836) <= 184108;
srom_1(4837) <= 83725;
srom_1(4838) <= 22287;
srom_1(4839) <= 81;
srom_1(4840) <= 17213;
srom_1(4841) <= 73600;
srom_1(4842) <= 168979;
srom_1(4843) <= 302903;
srom_1(4844) <= 474744;
srom_1(4845) <= 683696;
srom_1(4846) <= 928778;
srom_1(4847) <= 1208842;
srom_1(4848) <= 1522575;
srom_1(4849) <= 1868505;
srom_1(4850) <= 2245009;
srom_1(4851) <= 2650323;
srom_1(4852) <= 3082546;
srom_1(4853) <= 3539651;
srom_1(4854) <= 4019495;
srom_1(4855) <= 4519826;
srom_1(4856) <= 5038300;
srom_1(4857) <= 5572484;
srom_1(4858) <= 6119874;
srom_1(4859) <= 6677903;
srom_1(4860) <= 7243954;
srom_1(4861) <= 7815373;
srom_1(4862) <= 8389480;
srom_1(4863) <= 8963583;
srom_1(4864) <= 9534989;
srom_1(4865) <= 10101020;
srom_1(4866) <= 10659020;
srom_1(4867) <= 11206374;
srom_1(4868) <= 11740514;
srom_1(4869) <= 12258937;
srom_1(4870) <= 12759209;
srom_1(4871) <= 13238987;
srom_1(4872) <= 13696019;
srom_1(4873) <= 14128164;
srom_1(4874) <= 14533393;
srom_1(4875) <= 14909807;
srom_1(4876) <= 15255642;
srom_1(4877) <= 15569274;
srom_1(4878) <= 15849234;
srom_1(4879) <= 16094208;
srom_1(4880) <= 16303048;
srom_1(4881) <= 16474775;
srom_1(4882) <= 16608582;
srom_1(4883) <= 16703844;
srom_1(4884) <= 16760112;
srom_1(4885) <= 16777124;
srom_1(4886) <= 16754799;
srom_1(4887) <= 16693242;
srom_1(4888) <= 16592741;
srom_1(4889) <= 16453769;
srom_1(4890) <= 16276976;
srom_1(4891) <= 16063192;
srom_1(4892) <= 15813420;
srom_1(4893) <= 15528830;
srom_1(4894) <= 15210756;
srom_1(4895) <= 14860692;
srom_1(4896) <= 14480277;
srom_1(4897) <= 14071297;
srom_1(4898) <= 13635669;
srom_1(4899) <= 13175435;
srom_1(4900) <= 12692754;
srom_1(4901) <= 12189890;
srom_1(4902) <= 11669200;
srom_1(4903) <= 11133126;
srom_1(4904) <= 10584182;
srom_1(4905) <= 10024943;
srom_1(4906) <= 9458030;
srom_1(4907) <= 8886102;
srom_1(4908) <= 8311842;
srom_1(4909) <= 7737941;
srom_1(4910) <= 7167091;
srom_1(4911) <= 6601970;
srom_1(4912) <= 6045227;
srom_1(4913) <= 5499472;
srom_1(4914) <= 4967266;
srom_1(4915) <= 4451104;
srom_1(4916) <= 3953405;
srom_1(4917) <= 3476506;
srom_1(4918) <= 3022640;
srom_1(4919) <= 2593938;
srom_1(4920) <= 2192408;
srom_1(4921) <= 1819935;
srom_1(4922) <= 1478265;
srom_1(4923) <= 1168999;
srom_1(4924) <= 893589;
srom_1(4925) <= 653325;
srom_1(4926) <= 449335;
srom_1(4927) <= 282575;
srom_1(4928) <= 153827;
srom_1(4929) <= 63694;
srom_1(4930) <= 12600;
srom_1(4931) <= 784;
srom_1(4932) <= 28301;
srom_1(4933) <= 95023;
srom_1(4934) <= 200636;
srom_1(4935) <= 344645;
srom_1(4936) <= 526375;
srom_1(4937) <= 744974;
srom_1(4938) <= 999416;
srom_1(4939) <= 1288509;
srom_1(4940) <= 1610897;
srom_1(4941) <= 1965068;
srom_1(4942) <= 2349360;
srom_1(4943) <= 2761973;
srom_1(4944) <= 3200972;
srom_1(4945) <= 3664296;
srom_1(4946) <= 4149775;
srom_1(4947) <= 4655131;
srom_1(4948) <= 5177995;
srom_1(4949) <= 5715914;
srom_1(4950) <= 6266366;
srom_1(4951) <= 6826771;
srom_1(4952) <= 7394499;
srom_1(4953) <= 7966889;
srom_1(4954) <= 8541257;
srom_1(4955) <= 9114909;
srom_1(4956) <= 9685155;
srom_1(4957) <= 10249320;
srom_1(4958) <= 10804761;
srom_1(4959) <= 11348871;
srom_1(4960) <= 11879100;
srom_1(4961) <= 12392960;
srom_1(4962) <= 12888043;
srom_1(4963) <= 13362026;
srom_1(4964) <= 13812687;
srom_1(4965) <= 14237913;
srom_1(4966) <= 14635709;
srom_1(4967) <= 15004211;
srom_1(4968) <= 15341690;
srom_1(4969) <= 15646563;
srom_1(4970) <= 15917401;
srom_1(4971) <= 16152934;
srom_1(4972) <= 16352058;
srom_1(4973) <= 16513838;
srom_1(4974) <= 16637516;
srom_1(4975) <= 16722513;
srom_1(4976) <= 16768428;
srom_1(4977) <= 16775048;
srom_1(4978) <= 16742341;
srom_1(4979) <= 16670460;
srom_1(4980) <= 16559743;
srom_1(4981) <= 16410709;
srom_1(4982) <= 16224056;
srom_1(4983) <= 16000660;
srom_1(4984) <= 15741569;
srom_1(4985) <= 15447997;
srom_1(4986) <= 15121321;
srom_1(4987) <= 14763073;
srom_1(4988) <= 14374933;
srom_1(4989) <= 13958722;
srom_1(4990) <= 13516389;
srom_1(4991) <= 13050011;
srom_1(4992) <= 12561775;
srom_1(4993) <= 12053968;
srom_1(4994) <= 11528974;
srom_1(4995) <= 10989253;
srom_1(4996) <= 10437337;
srom_1(4997) <= 9875814;
srom_1(4998) <= 9307316;
srom_1(4999) <= 8734511;
srom_1(5000) <= 8160083;
srom_1(5001) <= 7586727;
srom_1(5002) <= 7017132;
srom_1(5003) <= 6453968;
srom_1(5004) <= 5899875;
srom_1(5005) <= 5357454;
srom_1(5006) <= 4829246;
srom_1(5007) <= 4317730;
srom_1(5008) <= 3825303;
srom_1(5009) <= 3354276;
srom_1(5010) <= 2906855;
srom_1(5011) <= 2485141;
srom_1(5012) <= 2091110;
srom_1(5013) <= 1726611;
srom_1(5014) <= 1393351;
srom_1(5015) <= 1092895;
srom_1(5016) <= 826651;
srom_1(5017) <= 595867;
srom_1(5018) <= 401627;
srom_1(5019) <= 244840;
srom_1(5020) <= 126242;
srom_1(5021) <= 46389;
srom_1(5022) <= 5655;
srom_1(5023) <= 4232;
srom_1(5024) <= 42127;
srom_1(5025) <= 119160;
srom_1(5026) <= 234972;
srom_1(5027) <= 389020;
srom_1(5028) <= 580580;
srom_1(5029) <= 808754;
srom_1(5030) <= 1072474;
srom_1(5031) <= 1370501;
srom_1(5032) <= 1701438;
srom_1(5033) <= 2063734;
srom_1(5034) <= 2455689;
srom_1(5035) <= 2875465;
srom_1(5036) <= 3321095;
srom_1(5037) <= 3790488;
srom_1(5038) <= 4281443;
srom_1(5039) <= 4791659;
srom_1(5040) <= 5318741;
srom_1(5041) <= 5860219;
srom_1(5042) <= 6413554;
srom_1(5043) <= 6976150;
srom_1(5044) <= 7545370;
srom_1(5045) <= 8118543;
srom_1(5046) <= 8692984;
srom_1(5047) <= 9265997;
srom_1(5048) <= 9834896;
srom_1(5049) <= 10397012;
srom_1(5050) <= 10949711;
srom_1(5051) <= 11490399;
srom_1(5052) <= 12016542;
srom_1(5053) <= 12525673;
srom_1(5054) <= 13015403;
srom_1(5055) <= 13483437;
srom_1(5056) <= 13927579;
srom_1(5057) <= 14345747;
srom_1(5058) <= 14735981;
srom_1(5059) <= 15096449;
srom_1(5060) <= 15425461;
srom_1(5061) <= 15721476;
srom_1(5062) <= 15983104;
srom_1(5063) <= 16209119;
srom_1(5064) <= 16398461;
srom_1(5065) <= 16550242;
srom_1(5066) <= 16663750;
srom_1(5067) <= 16738453;
srom_1(5068) <= 16774001;
srom_1(5069) <= 16770227;
srom_1(5070) <= 16727149;
srom_1(5071) <= 16644968;
srom_1(5072) <= 16524070;
srom_1(5073) <= 16365023;
srom_1(5074) <= 16168571;
srom_1(5075) <= 15935636;
srom_1(5076) <= 15667311;
srom_1(5077) <= 15364853;
srom_1(5078) <= 15029682;
srom_1(5079) <= 14663368;
srom_1(5080) <= 14267629;
srom_1(5081) <= 13844322;
srom_1(5082) <= 13395431;
srom_1(5083) <= 12923062;
srom_1(5084) <= 12429428;
srom_1(5085) <= 11916846;
srom_1(5086) <= 11387719;
srom_1(5087) <= 10844528;
srom_1(5088) <= 10289820;
srom_1(5089) <= 9726197;
srom_1(5090) <= 9156302;
srom_1(5091) <= 8582806;
srom_1(5092) <= 8008400;
srom_1(5093) <= 7435777;
srom_1(5094) <= 6867621;
srom_1(5095) <= 6306599;
srom_1(5096) <= 5755339;
srom_1(5097) <= 5216428;
srom_1(5098) <= 4692392;
srom_1(5099) <= 4185689;
srom_1(5100) <= 3698695;
srom_1(5101) <= 3233694;
srom_1(5102) <= 2792865;
srom_1(5103) <= 2378278;
srom_1(5104) <= 1991874;
srom_1(5105) <= 1635467;
srom_1(5106) <= 1310728;
srom_1(5107) <= 1019179;
srom_1(5108) <= 762189;
srom_1(5109) <= 540961;
srom_1(5110) <= 356533;
srom_1(5111) <= 209771;
srom_1(5112) <= 101362;
srom_1(5113) <= 31814;
srom_1(5114) <= 1455;
srom_1(5115) <= 10426;
srom_1(5116) <= 58685;
srom_1(5117) <= 146006;
srom_1(5118) <= 271979;
srom_1(5119) <= 436014;
srom_1(5120) <= 637341;
srom_1(5121) <= 875017;
srom_1(5122) <= 1147926;
srom_1(5123) <= 1454790;
srom_1(5124) <= 1794168;
srom_1(5125) <= 2164470;
srom_1(5126) <= 2563959;
srom_1(5127) <= 2990763;
srom_1(5128) <= 3442878;
srom_1(5129) <= 3918185;
srom_1(5130) <= 4414456;
srom_1(5131) <= 4929363;
srom_1(5132) <= 5460492;
srom_1(5133) <= 6005352;
srom_1(5134) <= 6561387;
srom_1(5135) <= 7125991;
srom_1(5136) <= 7696516;
srom_1(5137) <= 8270286;
srom_1(5138) <= 8844611;
srom_1(5139) <= 9416798;
srom_1(5140) <= 9984163;
srom_1(5141) <= 10544046;
srom_1(5142) <= 11093822;
srom_1(5143) <= 11630911;
srom_1(5144) <= 12152797;
srom_1(5145) <= 12657031;
srom_1(5146) <= 13141249;
srom_1(5147) <= 13603180;
srom_1(5148) <= 14040658;
srom_1(5149) <= 14451632;
srom_1(5150) <= 14834174;
srom_1(5151) <= 15186490;
srom_1(5152) <= 15506929;
srom_1(5153) <= 15793988;
srom_1(5154) <= 16046320;
srom_1(5155) <= 16262743;
srom_1(5156) <= 16442241;
srom_1(5157) <= 16583973;
srom_1(5158) <= 16687274;
srom_1(5159) <= 16751660;
srom_1(5160) <= 16776828;
srom_1(5161) <= 16762662;
srom_1(5162) <= 16709226;
srom_1(5163) <= 16616772;
srom_1(5164) <= 16485734;
srom_1(5165) <= 16316725;
srom_1(5166) <= 16110539;
srom_1(5167) <= 15868141;
srom_1(5168) <= 15590670;
srom_1(5169) <= 15279426;
srom_1(5170) <= 14935868;
srom_1(5171) <= 14561608;
srom_1(5172) <= 14158401;
srom_1(5173) <= 13728137;
srom_1(5174) <= 13272834;
srom_1(5175) <= 12794627;
srom_1(5176) <= 12295759;
srom_1(5177) <= 11778570;
srom_1(5178) <= 11245483;
srom_1(5179) <= 10698999;
srom_1(5180) <= 10141682;
srom_1(5181) <= 9576143;
srom_1(5182) <= 9005036;
srom_1(5183) <= 8431038;
srom_1(5184) <= 7856841;
srom_1(5185) <= 7285138;
srom_1(5186) <= 6718609;
srom_1(5187) <= 6159911;
srom_1(5188) <= 5611665;
srom_1(5189) <= 5076441;
srom_1(5190) <= 4556748;
srom_1(5191) <= 4055024;
srom_1(5192) <= 3573622;
srom_1(5193) <= 3114800;
srom_1(5194) <= 2680707;
srom_1(5195) <= 2273382;
srom_1(5196) <= 1894732;
srom_1(5197) <= 1546535;
srom_1(5198) <= 1230422;
srom_1(5199) <= 947877;
srom_1(5200) <= 700223;
srom_1(5201) <= 488624;
srom_1(5202) <= 314069;
srom_1(5203) <= 177380;
srom_1(5204) <= 79195;
srom_1(5205) <= 19976;
srom_1(5206) <= 1;
srom_1(5207) <= 19362;
srom_1(5208) <= 77970;
srom_1(5209) <= 175549;
srom_1(5210) <= 311642;
srom_1(5211) <= 485611;
srom_1(5212) <= 696640;
srom_1(5213) <= 943739;
srom_1(5214) <= 1225749;
srom_1(5215) <= 1541349;
srom_1(5216) <= 1889057;
srom_1(5217) <= 2267245;
srom_1(5218) <= 2674137;
srom_1(5219) <= 3107827;
srom_1(5220) <= 3566280;
srom_1(5221) <= 4047346;
srom_1(5222) <= 4548770;
srom_1(5223) <= 5068201;
srom_1(5224) <= 5603202;
srom_1(5225) <= 6151265;
srom_1(5226) <= 6709819;
srom_1(5227) <= 7276246;
srom_1(5228) <= 7847889;
srom_1(5229) <= 8422068;
srom_1(5230) <= 8996089;
srom_1(5231) <= 9567262;
srom_1(5232) <= 10132908;
srom_1(5233) <= 10690375;
srom_1(5234) <= 11237047;
srom_1(5235) <= 11770362;
srom_1(5236) <= 12287819;
srom_1(5237) <= 12786992;
srom_1(5238) <= 13265538;
srom_1(5239) <= 13721215;
srom_1(5240) <= 14151886;
srom_1(5241) <= 14555531;
srom_1(5242) <= 14930256;
srom_1(5243) <= 15274306;
srom_1(5244) <= 15586067;
srom_1(5245) <= 15864076;
srom_1(5246) <= 16107030;
srom_1(5247) <= 16313789;
srom_1(5248) <= 16483385;
srom_1(5249) <= 16615022;
srom_1(5250) <= 16708082;
srom_1(5251) <= 16762129;
srom_1(5252) <= 16776910;
srom_1(5253) <= 16752355;
srom_1(5254) <= 16688580;
srom_1(5255) <= 16585883;
srom_1(5256) <= 16444746;
srom_1(5257) <= 16265832;
srom_1(5258) <= 16049978;
srom_1(5259) <= 15798198;
srom_1(5260) <= 15511671;
srom_1(5261) <= 15191742;
srom_1(5262) <= 14839911;
srom_1(5263) <= 14457827;
srom_1(5264) <= 14047283;
srom_1(5265) <= 13610203;
srom_1(5266) <= 13148638;
srom_1(5267) <= 12664751;
srom_1(5268) <= 12160811;
srom_1(5269) <= 11639183;
srom_1(5270) <= 11102311;
srom_1(5271) <= 10552714;
srom_1(5272) <= 9992969;
srom_1(5273) <= 9425700;
srom_1(5274) <= 8853568;
srom_1(5275) <= 8279256;
srom_1(5276) <= 7705456;
srom_1(5277) <= 7134860;
srom_1(5278) <= 6570143;
srom_1(5279) <= 6013954;
srom_1(5280) <= 5468900;
srom_1(5281) <= 4937538;
srom_1(5282) <= 4422358;
srom_1(5283) <= 3925778;
srom_1(5284) <= 3450126;
srom_1(5285) <= 2997632;
srom_1(5286) <= 2570418;
srom_1(5287) <= 2170488;
srom_1(5288) <= 1799716;
srom_1(5289) <= 1459842;
srom_1(5290) <= 1152460;
srom_1(5291) <= 879010;
srom_1(5292) <= 640775;
srom_1(5293) <= 438873;
srom_1(5294) <= 274249;
srom_1(5295) <= 147677;
srom_1(5296) <= 59749;
srom_1(5297) <= 10878;
srom_1(5298) <= 1293;
srom_1(5299) <= 31039;
srom_1(5300) <= 99976;
srom_1(5301) <= 207782;
srom_1(5302) <= 353950;
srom_1(5303) <= 537796;
srom_1(5304) <= 758457;
srom_1(5305) <= 1014898;
srom_1(5306) <= 1305917;
srom_1(5307) <= 1630150;
srom_1(5308) <= 1986075;
srom_1(5309) <= 2372023;
srom_1(5310) <= 2786186;
srom_1(5311) <= 3226620;
srom_1(5312) <= 3691260;
srom_1(5313) <= 4177928;
srom_1(5314) <= 4684342;
srom_1(5315) <= 5208125;
srom_1(5316) <= 5746824;
srom_1(5317) <= 6297910;
srom_1(5318) <= 6858801;
srom_1(5319) <= 7426865;
srom_1(5320) <= 7999439;
srom_1(5321) <= 8573838;
srom_1(5322) <= 9147369;
srom_1(5323) <= 9717341;
srom_1(5324) <= 10281082;
srom_1(5325) <= 10835949;
srom_1(5326) <= 11379340;
srom_1(5327) <= 11908706;
srom_1(5328) <= 12421565;
srom_1(5329) <= 12915512;
srom_1(5330) <= 13388231;
srom_1(5331) <= 13837505;
srom_1(5332) <= 14261227;
srom_1(5333) <= 14657411;
srom_1(5334) <= 15024198;
srom_1(5335) <= 15359868;
srom_1(5336) <= 15662848;
srom_1(5337) <= 15931716;
srom_1(5338) <= 16165212;
srom_1(5339) <= 16362241;
srom_1(5340) <= 16521879;
srom_1(5341) <= 16643377;
srom_1(5342) <= 16726165;
srom_1(5343) <= 16769856;
srom_1(5344) <= 16774244;
srom_1(5345) <= 16739310;
srom_1(5346) <= 16665216;
srom_1(5347) <= 16552310;
srom_1(5348) <= 16401121;
srom_1(5349) <= 16212359;
srom_1(5350) <= 15986909;
srom_1(5351) <= 15725828;
srom_1(5352) <= 15430340;
srom_1(5353) <= 15101831;
srom_1(5354) <= 14741842;
srom_1(5355) <= 14352060;
srom_1(5356) <= 13934313;
srom_1(5357) <= 13490560;
srom_1(5358) <= 13022883;
srom_1(5359) <= 12533474;
srom_1(5360) <= 12024628;
srom_1(5361) <= 11498732;
srom_1(5362) <= 10958251;
srom_1(5363) <= 10405720;
srom_1(5364) <= 9843731;
srom_1(5365) <= 9274918;
srom_1(5366) <= 8701948;
srom_1(5367) <= 8127509;
srom_1(5368) <= 7554295;
srom_1(5369) <= 6984993;
srom_1(5370) <= 6422273;
srom_1(5371) <= 5868774;
srom_1(5372) <= 5327091;
srom_1(5373) <= 4799764;
srom_1(5374) <= 4289267;
srom_1(5375) <= 3797994;
srom_1(5376) <= 3328247;
srom_1(5377) <= 2882230;
srom_1(5378) <= 2462034;
srom_1(5379) <= 2069630;
srom_1(5380) <= 1706858;
srom_1(5381) <= 1375418;
srom_1(5382) <= 1076866;
srom_1(5383) <= 812602;
srom_1(5384) <= 583863;
srom_1(5385) <= 391724;
srom_1(5386) <= 237085;
srom_1(5387) <= 120672;
srom_1(5388) <= 43029;
srom_1(5389) <= 4522;
srom_1(5390) <= 5331;
srom_1(5391) <= 45451;
srom_1(5392) <= 124696;
srom_1(5393) <= 242693;
srom_1(5394) <= 398889;
srom_1(5395) <= 592551;
srom_1(5396) <= 822772;
srom_1(5397) <= 1088472;
srom_1(5398) <= 1388404;
srom_1(5399) <= 1721163;
srom_1(5400) <= 2085188;
srom_1(5401) <= 2478772;
srom_1(5402) <= 2900068;
srom_1(5403) <= 3347103;
srom_1(5404) <= 3817779;
srom_1(5405) <= 4309889;
srom_1(5406) <= 4821126;
srom_1(5407) <= 5349091;
srom_1(5408) <= 5891310;
srom_1(5409) <= 6445240;
srom_1(5410) <= 7008283;
srom_1(5411) <= 7577799;
srom_1(5412) <= 8151116;
srom_1(5413) <= 8725548;
srom_1(5414) <= 9298399;
srom_1(5415) <= 9866984;
srom_1(5416) <= 10428637;
srom_1(5417) <= 10980723;
srom_1(5418) <= 11520654;
srom_1(5419) <= 12045897;
srom_1(5420) <= 12553991;
srom_1(5421) <= 13042551;
srom_1(5422) <= 13509287;
srom_1(5423) <= 13952011;
srom_1(5424) <= 14368646;
srom_1(5425) <= 14757239;
srom_1(5426) <= 15115966;
srom_1(5427) <= 15443147;
srom_1(5428) <= 15737247;
srom_1(5429) <= 15996887;
srom_1(5430) <= 16220848;
srom_1(5431) <= 16408082;
srom_1(5432) <= 16557709;
srom_1(5433) <= 16669029;
srom_1(5434) <= 16741519;
srom_1(5435) <= 16774840;
srom_1(5436) <= 16768834;
srom_1(5437) <= 16723531;
srom_1(5438) <= 16639142;
srom_1(5439) <= 16516064;
srom_1(5440) <= 16354873;
srom_1(5441) <= 16156326;
srom_1(5442) <= 15921353;
srom_1(5443) <= 15651057;
srom_1(5444) <= 15346704;
srom_1(5445) <= 15009723;
srom_1(5446) <= 14641692;
srom_1(5447) <= 14244339;
srom_1(5448) <= 13819527;
srom_1(5449) <= 13369247;
srom_1(5450) <= 12895611;
srom_1(5451) <= 12400840;
srom_1(5452) <= 11887255;
srom_1(5453) <= 11357263;
srom_1(5454) <= 10813350;
srom_1(5455) <= 10258066;
srom_1(5456) <= 9694016;
srom_1(5457) <= 9123845;
srom_1(5458) <= 8550226;
srom_1(5459) <= 7975849;
srom_1(5460) <= 7403407;
srom_1(5461) <= 6835585;
srom_1(5462) <= 6275046;
srom_1(5463) <= 5724418;
srom_1(5464) <= 5186284;
srom_1(5465) <= 4663166;
srom_1(5466) <= 4157518;
srom_1(5467) <= 3671712;
srom_1(5468) <= 3208024;
srom_1(5469) <= 2768630;
srom_1(5470) <= 2355590;
srom_1(5471) <= 1970840;
srom_1(5472) <= 1616186;
srom_1(5473) <= 1293290;
srom_1(5474) <= 1003667;
srom_1(5475) <= 748674;
srom_1(5476) <= 529507;
srom_1(5477) <= 347194;
srom_1(5478) <= 202590;
srom_1(5479) <= 96374;
srom_1(5480) <= 29042;
srom_1(5481) <= 911;
srom_1(5482) <= 12113;
srom_1(5483) <= 62596;
srom_1(5484) <= 152121;
srom_1(5485) <= 280271;
srom_1(5486) <= 446443;
srom_1(5487) <= 649859;
srom_1(5488) <= 889564;
srom_1(5489) <= 1164435;
srom_1(5490) <= 1473183;
srom_1(5491) <= 1814360;
srom_1(5492) <= 2186365;
srom_1(5493) <= 2587455;
srom_1(5494) <= 3015748;
srom_1(5495) <= 3469237;
srom_1(5496) <= 3945794;
srom_1(5497) <= 4443185;
srom_1(5498) <= 4959077;
srom_1(5499) <= 5491052;
srom_1(5500) <= 6036615;
srom_1(5501) <= 6593206;
srom_1(5502) <= 7158217;
srom_1(5503) <= 7728998;
srom_1(5504) <= 8302872;
srom_1(5505) <= 8877147;
srom_1(5506) <= 9449132;
srom_1(5507) <= 10016144;
srom_1(5508) <= 10575524;
srom_1(5509) <= 11124648;
srom_1(5510) <= 11660942;
srom_1(5511) <= 12181891;
srom_1(5512) <= 12685052;
srom_1(5513) <= 13168066;
srom_1(5514) <= 13628667;
srom_1(5515) <= 14064695;
srom_1(5516) <= 14474107;
srom_1(5517) <= 14854981;
srom_1(5518) <= 15205533;
srom_1(5519) <= 15524117;
srom_1(5520) <= 15809241;
srom_1(5521) <= 16059566;
srom_1(5522) <= 16273920;
srom_1(5523) <= 16451297;
srom_1(5524) <= 16590866;
srom_1(5525) <= 16691971;
srom_1(5526) <= 16754138;
srom_1(5527) <= 16777077;
srom_1(5528) <= 16760680;
srom_1(5529) <= 16705023;
srom_1(5530) <= 16610367;
srom_1(5531) <= 16477157;
srom_1(5532) <= 16306017;
srom_1(5533) <= 16097749;
srom_1(5534) <= 15853330;
srom_1(5535) <= 15573907;
srom_1(5536) <= 15260790;
srom_1(5537) <= 14915446;
srom_1(5538) <= 14539496;
srom_1(5539) <= 14134702;
srom_1(5540) <= 13702963;
srom_1(5541) <= 13246303;
srom_1(5542) <= 12766864;
srom_1(5543) <= 12266893;
srom_1(5544) <= 11748736;
srom_1(5545) <= 11214822;
srom_1(5546) <= 10667655;
srom_1(5547) <= 10109800;
srom_1(5548) <= 9543875;
srom_1(5549) <= 8972532;
srom_1(5550) <= 8398450;
srom_1(5551) <= 7824323;
srom_1(5552) <= 7252841;
srom_1(5553) <= 6686686;
srom_1(5554) <= 6128512;
srom_1(5555) <= 5580936;
srom_1(5556) <= 5046526;
srom_1(5557) <= 4527788;
srom_1(5558) <= 4027155;
srom_1(5559) <= 3546974;
srom_1(5560) <= 3089497;
srom_1(5561) <= 2656870;
srom_1(5562) <= 2251121;
srom_1(5563) <= 1874152;
srom_1(5564) <= 1527732;
srom_1(5565) <= 1213485;
srom_1(5566) <= 932885;
srom_1(5567) <= 687247;
srom_1(5568) <= 477724;
srom_1(5569) <= 305297;
srom_1(5570) <= 170776;
srom_1(5571) <= 74790;
srom_1(5572) <= 17792;
srom_1(5573) <= 47;
srom_1(5574) <= 21638;
srom_1(5575) <= 82466;
srom_1(5576) <= 182243;
srom_1(5577) <= 320503;
srom_1(5578) <= 496598;
srom_1(5579) <= 709700;
srom_1(5580) <= 958812;
srom_1(5581) <= 1242764;
srom_1(5582) <= 1560226;
srom_1(5583) <= 1909708;
srom_1(5584) <= 2289573;
srom_1(5585) <= 2698037;
srom_1(5586) <= 3133187;
srom_1(5587) <= 3592981;
srom_1(5588) <= 4075263;
srom_1(5589) <= 4577773;
srom_1(5590) <= 5098152;
srom_1(5591) <= 5633962;
srom_1(5592) <= 6182689;
srom_1(5593) <= 6741760;
srom_1(5594) <= 7308554;
srom_1(5595) <= 7880413;
srom_1(5596) <= 8454655;
srom_1(5597) <= 9028587;
srom_1(5598) <= 9599518;
srom_1(5599) <= 10164771;
srom_1(5600) <= 10721694;
srom_1(5601) <= 11267677;
srom_1(5602) <= 11800159;
srom_1(5603) <= 12316643;
srom_1(5604) <= 12814707;
srom_1(5605) <= 13292016;
srom_1(5606) <= 13746331;
srom_1(5607) <= 14175522;
srom_1(5608) <= 14577575;
srom_1(5609) <= 14950607;
srom_1(5610) <= 15292867;
srom_1(5611) <= 15602751;
srom_1(5612) <= 15878805;
srom_1(5613) <= 16119735;
srom_1(5614) <= 16324411;
srom_1(5615) <= 16491873;
srom_1(5616) <= 16621337;
srom_1(5617) <= 16712194;
srom_1(5618) <= 16764019;
srom_1(5619) <= 16776569;
srom_1(5620) <= 16749785;
srom_1(5621) <= 16683792;
srom_1(5622) <= 16578901;
srom_1(5623) <= 16435602;
srom_1(5624) <= 16254568;
srom_1(5625) <= 16036648;
srom_1(5626) <= 15782864;
srom_1(5627) <= 15494405;
srom_1(5628) <= 15172625;
srom_1(5629) <= 14819033;
srom_1(5630) <= 14435286;
srom_1(5631) <= 14023184;
srom_1(5632) <= 13584659;
srom_1(5633) <= 13121769;
srom_1(5634) <= 12636683;
srom_1(5635) <= 12131676;
srom_1(5636) <= 11609117;
srom_1(5637) <= 11071455;
srom_1(5638) <= 10521213;
srom_1(5639) <= 9960971;
srom_1(5640) <= 9393355;
srom_1(5641) <= 8821027;
srom_1(5642) <= 8246672;
srom_1(5643) <= 7672982;
srom_1(5644) <= 7102648;
srom_1(5645) <= 6538344;
srom_1(5646) <= 5982717;
srom_1(5647) <= 5438372;
srom_1(5648) <= 4907861;
srom_1(5649) <= 4393673;
srom_1(5650) <= 3898219;
srom_1(5651) <= 3423821;
srom_1(5652) <= 2972706;
srom_1(5653) <= 2546987;
srom_1(5654) <= 2148661;
srom_1(5655) <= 1779597;
srom_1(5656) <= 1441525;
srom_1(5657) <= 1136029;
srom_1(5658) <= 864544;
srom_1(5659) <= 628342;
srom_1(5660) <= 428530;
srom_1(5661) <= 266046;
srom_1(5662) <= 141651;
srom_1(5663) <= 55929;
srom_1(5664) <= 9282;
srom_1(5665) <= 1928;
srom_1(5666) <= 33903;
srom_1(5667) <= 105055;
srom_1(5668) <= 215052;
srom_1(5669) <= 363377;
srom_1(5670) <= 549336;
srom_1(5671) <= 772055;
srom_1(5672) <= 1030492;
srom_1(5673) <= 1323432;
srom_1(5674) <= 1649504;
srom_1(5675) <= 2007178;
srom_1(5676) <= 2394777;
srom_1(5677) <= 2810483;
srom_1(5678) <= 3252346;
srom_1(5679) <= 3718295;
srom_1(5680) <= 4206145;
srom_1(5681) <= 4713608;
srom_1(5682) <= 5238304;
srom_1(5683) <= 5777773;
srom_1(5684) <= 6329485;
srom_1(5685) <= 6890853;
srom_1(5686) <= 7459245;
srom_1(5687) <= 8031995;
srom_1(5688) <= 8606416;
srom_1(5689) <= 9179817;
srom_1(5690) <= 9749507;
srom_1(5691) <= 10312816;
srom_1(5692) <= 10867101;
srom_1(5693) <= 11409764;
srom_1(5694) <= 11938259;
srom_1(5695) <= 12450109;
srom_1(5696) <= 12942913;
srom_1(5697) <= 13414361;
srom_1(5698) <= 13862241;
srom_1(5699) <= 14284453;
srom_1(5700) <= 14679018;
srom_1(5701) <= 15044084;
srom_1(5702) <= 15377941;
srom_1(5703) <= 15679023;
srom_1(5704) <= 15945917;
srom_1(5705) <= 16177372;
srom_1(5706) <= 16372303;
srom_1(5707) <= 16529796;
srom_1(5708) <= 16649112;
srom_1(5709) <= 16729692;
srom_1(5710) <= 16771157;
srom_1(5711) <= 16773314;
srom_1(5712) <= 16736152;
srom_1(5713) <= 16659846;
srom_1(5714) <= 16544753;
srom_1(5715) <= 16391413;
srom_1(5716) <= 16200544;
srom_1(5717) <= 15973044;
srom_1(5718) <= 15709977;
srom_1(5719) <= 15412577;
srom_1(5720) <= 15082240;
srom_1(5721) <= 14720514;
srom_1(5722) <= 14329096;
srom_1(5723) <= 13909820;
srom_1(5724) <= 13464654;
srom_1(5725) <= 12995685;
srom_1(5726) <= 12505111;
srom_1(5727) <= 11995233;
srom_1(5728) <= 11468443;
srom_1(5729) <= 10927211;
srom_1(5730) <= 10374074;
srom_1(5731) <= 9811626;
srom_1(5732) <= 9242506;
srom_1(5733) <= 8669381;
srom_1(5734) <= 8094939;
srom_1(5735) <= 7521875;
srom_1(5736) <= 6952875;
srom_1(5737) <= 6390608;
srom_1(5738) <= 5837710;
srom_1(5739) <= 5296774;
srom_1(5740) <= 4770337;
srom_1(5741) <= 4260867;
srom_1(5742) <= 3770753;
srom_1(5743) <= 3302294;
srom_1(5744) <= 2857687;
srom_1(5745) <= 2439016;
srom_1(5746) <= 2048244;
srom_1(5747) <= 1687205;
srom_1(5748) <= 1357591;
srom_1(5749) <= 1060948;
srom_1(5750) <= 798667;
srom_1(5751) <= 571977;
srom_1(5752) <= 381943;
srom_1(5753) <= 229454;
srom_1(5754) <= 115227;
srom_1(5755) <= 39796;
srom_1(5756) <= 3515;
srom_1(5757) <= 6556;
srom_1(5758) <= 48902;
srom_1(5759) <= 130356;
srom_1(5760) <= 250536;
srom_1(5761) <= 408879;
srom_1(5762) <= 604641;
srom_1(5763) <= 836904;
srom_1(5764) <= 1104580;
srom_1(5765) <= 1406414;
srom_1(5766) <= 1740989;
srom_1(5767) <= 2106737;
srom_1(5768) <= 2501944;
srom_1(5769) <= 2924754;
srom_1(5770) <= 3373187;
srom_1(5771) <= 3845139;
srom_1(5772) <= 4338396;
srom_1(5773) <= 4850646;
srom_1(5774) <= 5379488;
srom_1(5775) <= 5922439;
srom_1(5776) <= 6476956;
srom_1(5777) <= 7040437;
srom_1(5778) <= 7610240;
srom_1(5779) <= 8183693;
srom_1(5780) <= 8758107;
srom_1(5781) <= 9330788;
srom_1(5782) <= 9899051;
srom_1(5783) <= 10460231;
srom_1(5784) <= 11011696;
srom_1(5785) <= 11550861;
srom_1(5786) <= 12075197;
srom_1(5787) <= 12582245;
srom_1(5788) <= 13069628;
srom_1(5789) <= 13535060;
srom_1(5790) <= 13976359;
srom_1(5791) <= 14391454;
srom_1(5792) <= 14778400;
srom_1(5793) <= 15135383;
srom_1(5794) <= 15460727;
srom_1(5795) <= 15752908;
srom_1(5796) <= 16010554;
srom_1(5797) <= 16232459;
srom_1(5798) <= 16417582;
srom_1(5799) <= 16565054;
srom_1(5800) <= 16674183;
srom_1(5801) <= 16744459;
srom_1(5802) <= 16775551;
srom_1(5803) <= 16767315;
srom_1(5804) <= 16719787;
srom_1(5805) <= 16633191;
srom_1(5806) <= 16507934;
srom_1(5807) <= 16344603;
srom_1(5808) <= 16143963;
srom_1(5809) <= 15906956;
srom_1(5810) <= 15634692;
srom_1(5811) <= 15328450;
srom_1(5812) <= 14989663;
srom_1(5813) <= 14619923;
srom_1(5814) <= 14220961;
srom_1(5815) <= 13794650;
srom_1(5816) <= 13342987;
srom_1(5817) <= 12868092;
srom_1(5818) <= 12372191;
srom_1(5819) <= 11857610;
srom_1(5820) <= 11326761;
srom_1(5821) <= 10782135;
srom_1(5822) <= 10226284;
srom_1(5823) <= 9661816;
srom_1(5824) <= 9091377;
srom_1(5825) <= 8517643;
srom_1(5826) <= 7943303;
srom_1(5827) <= 7371052;
srom_1(5828) <= 6803573;
srom_1(5829) <= 6243526;
srom_1(5830) <= 5693538;
srom_1(5831) <= 5156188;
srom_1(5832) <= 4633997;
srom_1(5833) <= 4129412;
srom_1(5834) <= 3644799;
srom_1(5835) <= 3182432;
srom_1(5836) <= 2744479;
srom_1(5837) <= 2332993;
srom_1(5838) <= 1949904;
srom_1(5839) <= 1597008;
srom_1(5840) <= 1275960;
srom_1(5841) <= 988266;
srom_1(5842) <= 735274;
srom_1(5843) <= 518172;
srom_1(5844) <= 337977;
srom_1(5845) <= 195534;
srom_1(5846) <= 91511;
srom_1(5847) <= 26396;
srom_1(5848) <= 494;
srom_1(5849) <= 13927;
srom_1(5850) <= 66632;
srom_1(5851) <= 158361;
srom_1(5852) <= 288685;
srom_1(5853) <= 456992;
srom_1(5854) <= 662494;
srom_1(5855) <= 904225;
srom_1(5856) <= 1181054;
srom_1(5857) <= 1491681;
srom_1(5858) <= 1834650;
srom_1(5859) <= 2208353;
srom_1(5860) <= 2611038;
srom_1(5861) <= 3040815;
srom_1(5862) <= 3495670;
srom_1(5863) <= 3973469;
srom_1(5864) <= 4471973;
srom_1(5865) <= 4988843;
srom_1(5866) <= 5521656;
srom_1(5867) <= 6067913;
srom_1(5868) <= 6625052;
srom_1(5869) <= 7190462;
srom_1(5870) <= 7761490;
srom_1(5871) <= 8335458;
srom_1(5872) <= 8909676;
srom_1(5873) <= 9481450;
srom_1(5874) <= 10048100;
srom_1(5875) <= 10606968;
srom_1(5876) <= 11155433;
srom_1(5877) <= 11690923;
srom_1(5878) <= 12210928;
srom_1(5879) <= 12713009;
srom_1(5880) <= 13194811;
srom_1(5881) <= 13654075;
srom_1(5882) <= 14088647;
srom_1(5883) <= 14496490;
srom_1(5884) <= 14875691;
srom_1(5885) <= 15224472;
srom_1(5886) <= 15541197;
srom_1(5887) <= 15824382;
srom_1(5888) <= 16072697;
srom_1(5889) <= 16284979;
srom_1(5890) <= 16460232;
srom_1(5891) <= 16597634;
srom_1(5892) <= 16696542;
srom_1(5893) <= 16756491;
srom_1(5894) <= 16777200;
srom_1(5895) <= 16758572;
srom_1(5896) <= 16700694;
srom_1(5897) <= 16603838;
srom_1(5898) <= 16468458;
srom_1(5899) <= 16295189;
srom_1(5900) <= 16084843;
srom_1(5901) <= 15838407;
srom_1(5902) <= 15557036;
srom_1(5903) <= 15242050;
srom_1(5904) <= 14894926;
srom_1(5905) <= 14517291;
srom_1(5906) <= 14110917;
srom_1(5907) <= 13677709;
srom_1(5908) <= 13219699;
srom_1(5909) <= 12739033;
srom_1(5910) <= 12237968;
srom_1(5911) <= 11718851;
srom_1(5912) <= 11184118;
srom_1(5913) <= 10636275;
srom_1(5914) <= 10077893;
srom_1(5915) <= 9511589;
srom_1(5916) <= 8940018;
srom_1(5917) <= 8365862;
srom_1(5918) <= 7791813;
srom_1(5919) <= 7220562;
srom_1(5920) <= 6654789;
srom_1(5921) <= 6097146;
srom_1(5922) <= 5550248;
srom_1(5923) <= 5016661;
srom_1(5924) <= 4498886;
srom_1(5925) <= 3999351;
srom_1(5926) <= 3520399;
srom_1(5927) <= 3064275;
srom_1(5928) <= 2633119;
srom_1(5929) <= 2228952;
srom_1(5930) <= 1853671;
srom_1(5931) <= 1509033;
srom_1(5932) <= 1196657;
srom_1(5933) <= 918006;
srom_1(5934) <= 674387;
srom_1(5935) <= 466943;
srom_1(5936) <= 296646;
srom_1(5937) <= 164295;
srom_1(5938) <= 70511;
srom_1(5939) <= 15734;
srom_1(5940) <= 219;
srom_1(5941) <= 24041;
srom_1(5942) <= 87086;
srom_1(5943) <= 189061;
srom_1(5944) <= 329486;
srom_1(5945) <= 507703;
srom_1(5946) <= 722876;
srom_1(5947) <= 973997;
srom_1(5948) <= 1259887;
srom_1(5949) <= 1579206;
srom_1(5950) <= 1930457;
srom_1(5951) <= 2311992;
srom_1(5952) <= 2722023;
srom_1(5953) <= 3158626;
srom_1(5954) <= 3619755;
srom_1(5955) <= 4103246;
srom_1(5956) <= 4606832;
srom_1(5957) <= 5128153;
srom_1(5958) <= 5664763;
srom_1(5959) <= 6214146;
srom_1(5960) <= 6773726;
srom_1(5961) <= 7340879;
srom_1(5962) <= 7912945;
srom_1(5963) <= 8487241;
srom_1(5964) <= 9061075;
srom_1(5965) <= 9631755;
srom_1(5966) <= 10196606;
srom_1(5967) <= 10752979;
srom_1(5968) <= 11298264;
srom_1(5969) <= 11829904;
srom_1(5970) <= 12345408;
srom_1(5971) <= 12842356;
srom_1(5972) <= 13318420;
srom_1(5973) <= 13771366;
srom_1(5974) <= 14199070;
srom_1(5975) <= 14599527;
srom_1(5976) <= 14970858;
srom_1(5977) <= 15311324;
srom_1(5978) <= 15619326;
srom_1(5979) <= 15893421;
srom_1(5980) <= 16132323;
srom_1(5981) <= 16334913;
srom_1(5982) <= 16500239;
srom_1(5983) <= 16627528;
srom_1(5984) <= 16716181;
srom_1(5985) <= 16765783;
srom_1(5986) <= 16776102;
srom_1(5987) <= 16747089;
srom_1(5988) <= 16678880;
srom_1(5989) <= 16571795;
srom_1(5990) <= 16426336;
srom_1(5991) <= 16243186;
srom_1(5992) <= 16023203;
srom_1(5993) <= 15767419;
srom_1(5994) <= 15477032;
srom_1(5995) <= 15153406;
srom_1(5996) <= 14798058;
srom_1(5997) <= 14412653;
srom_1(5998) <= 13998999;
srom_1(5999) <= 13559037;
srom_1(6000) <= 13094828;
srom_1(6001) <= 12608550;
srom_1(6002) <= 12102484;
srom_1(6003) <= 11579002;
srom_1(6004) <= 11040559;
srom_1(6005) <= 10489680;
srom_1(6006) <= 9928949;
srom_1(6007) <= 9360994;
srom_1(6008) <= 8788479;
srom_1(6009) <= 8214090;
srom_1(6010) <= 7640518;
srom_1(6011) <= 7070455;
srom_1(6012) <= 6506573;
srom_1(6013) <= 5951516;
srom_1(6014) <= 5407888;
srom_1(6015) <= 4878238;
srom_1(6016) <= 4365048;
srom_1(6017) <= 3870727;
srom_1(6018) <= 3397592;
srom_1(6019) <= 2947861;
srom_1(6020) <= 2523643;
srom_1(6021) <= 2126929;
srom_1(6022) <= 1759577;
srom_1(6023) <= 1423312;
srom_1(6024) <= 1119709;
srom_1(6025) <= 850192;
srom_1(6026) <= 616026;
srom_1(6027) <= 418308;
srom_1(6028) <= 257965;
srom_1(6029) <= 135750;
srom_1(6030) <= 52235;
srom_1(6031) <= 7812;
srom_1(6032) <= 2690;
srom_1(6033) <= 36892;
srom_1(6034) <= 110259;
srom_1(6035) <= 222445;
srom_1(6036) <= 372925;
srom_1(6037) <= 560994;
srom_1(6038) <= 785769;
srom_1(6039) <= 1046196;
srom_1(6040) <= 1341054;
srom_1(6041) <= 1668961;
srom_1(6042) <= 2028378;
srom_1(6043) <= 2417621;
srom_1(6044) <= 2834864;
srom_1(6045) <= 3278150;
srom_1(6046) <= 3745401;
srom_1(6047) <= 4234425;
srom_1(6048) <= 4742930;
srom_1(6049) <= 5268530;
srom_1(6050) <= 5808762;
srom_1(6051) <= 6361092;
srom_1(6052) <= 6922929;
srom_1(6053) <= 7491639;
srom_1(6054) <= 8064556;
srom_1(6055) <= 8638992;
srom_1(6056) <= 9212253;
srom_1(6057) <= 9781653;
srom_1(6058) <= 10344520;
srom_1(6059) <= 10898215;
srom_1(6060) <= 11440142;
srom_1(6061) <= 11967759;
srom_1(6062) <= 12478592;
srom_1(6063) <= 12970246;
srom_1(6064) <= 13440415;
srom_1(6065) <= 13886894;
srom_1(6066) <= 14307590;
srom_1(6067) <= 14700530;
srom_1(6068) <= 15063870;
srom_1(6069) <= 15395909;
srom_1(6070) <= 15695088;
srom_1(6071) <= 15960004;
srom_1(6072) <= 16189415;
srom_1(6073) <= 16382245;
srom_1(6074) <= 16537591;
srom_1(6075) <= 16654723;
srom_1(6076) <= 16733093;
srom_1(6077) <= 16772332;
srom_1(6078) <= 16772257;
srom_1(6079) <= 16732869;
srom_1(6080) <= 16654351;
srom_1(6081) <= 16537073;
srom_1(6082) <= 16381583;
srom_1(6083) <= 16188612;
srom_1(6084) <= 15959063;
srom_1(6085) <= 15694015;
srom_1(6086) <= 15394708;
srom_1(6087) <= 15062548;
srom_1(6088) <= 14699091;
srom_1(6089) <= 14306042;
srom_1(6090) <= 13885245;
srom_1(6091) <= 13438671;
srom_1(6092) <= 12968417;
srom_1(6093) <= 12476686;
srom_1(6094) <= 11965784;
srom_1(6095) <= 11438108;
srom_1(6096) <= 10896132;
srom_1(6097) <= 10342397;
srom_1(6098) <= 9779500;
srom_1(6099) <= 9210081;
srom_1(6100) <= 8636809;
srom_1(6101) <= 8062374;
srom_1(6102) <= 7489468;
srom_1(6103) <= 6920779;
srom_1(6104) <= 6358973;
srom_1(6105) <= 5806685;
srom_1(6106) <= 5266504;
srom_1(6107) <= 4740964;
srom_1(6108) <= 4232528;
srom_1(6109) <= 3743582;
srom_1(6110) <= 3276419;
srom_1(6111) <= 2833228;
srom_1(6112) <= 2416088;
srom_1(6113) <= 2026955;
srom_1(6114) <= 1667654;
srom_1(6115) <= 1339870;
srom_1(6116) <= 1045140;
srom_1(6117) <= 784846;
srom_1(6118) <= 560209;
srom_1(6119) <= 372282;
srom_1(6120) <= 221946;
srom_1(6121) <= 109906;
srom_1(6122) <= 36688;
srom_1(6123) <= 2635;
srom_1(6124) <= 7907;
srom_1(6125) <= 52479;
srom_1(6126) <= 136141;
srom_1(6127) <= 258503;
srom_1(6128) <= 418989;
srom_1(6129) <= 616847;
srom_1(6130) <= 851150;
srom_1(6131) <= 1120799;
srom_1(6132) <= 1424529;
srom_1(6133) <= 1760915;
srom_1(6134) <= 2128382;
srom_1(6135) <= 2525204;
srom_1(6136) <= 2949523;
srom_1(6137) <= 3399347;
srom_1(6138) <= 3872567;
srom_1(6139) <= 4366964;
srom_1(6140) <= 4880221;
srom_1(6141) <= 5409929;
srom_1(6142) <= 5953606;
srom_1(6143) <= 6508701;
srom_1(6144) <= 7072611;
srom_1(6145) <= 7642693;
srom_1(6146) <= 8216272;
srom_1(6147) <= 8790660;
srom_1(6148) <= 9363162;
srom_1(6149) <= 9931095;
srom_1(6150) <= 10491794;
srom_1(6151) <= 11042630;
srom_1(6152) <= 11581021;
srom_1(6153) <= 12104441;
srom_1(6154) <= 12610437;
srom_1(6155) <= 13096635;
srom_1(6156) <= 13560756;
srom_1(6157) <= 14000622;
srom_1(6158) <= 14414172;
srom_1(6159) <= 14799466;
srom_1(6160) <= 15154697;
srom_1(6161) <= 15478200;
srom_1(6162) <= 15768457;
srom_1(6163) <= 16024107;
srom_1(6164) <= 16243952;
srom_1(6165) <= 16426961;
srom_1(6166) <= 16572275;
srom_1(6167) <= 16679213;
srom_1(6168) <= 16747273;
srom_1(6169) <= 16776137;
srom_1(6170) <= 16765669;
srom_1(6171) <= 16715917;
srom_1(6172) <= 16627117;
srom_1(6173) <= 16499683;
srom_1(6174) <= 16334213;
srom_1(6175) <= 16131484;
srom_1(6176) <= 15892445;
srom_1(6177) <= 15618219;
srom_1(6178) <= 15310090;
srom_1(6179) <= 14969505;
srom_1(6180) <= 14598059;
srom_1(6181) <= 14197495;
srom_1(6182) <= 13769691;
srom_1(6183) <= 13316653;
srom_1(6184) <= 12840506;
srom_1(6185) <= 12343483;
srom_1(6186) <= 11827913;
srom_1(6187) <= 11296216;
srom_1(6188) <= 10750884;
srom_1(6189) <= 10194474;
srom_1(6190) <= 9629596;
srom_1(6191) <= 9058899;
srom_1(6192) <= 8485058;
srom_1(6193) <= 7910765;
srom_1(6194) <= 7338713;
srom_1(6195) <= 6771584;
srom_1(6196) <= 6212038;
srom_1(6197) <= 5662698;
srom_1(6198) <= 5126142;
srom_1(6199) <= 4604884;
srom_1(6200) <= 4101369;
srom_1(6201) <= 3617959;
srom_1(6202) <= 3156919;
srom_1(6203) <= 2720413;
srom_1(6204) <= 2310487;
srom_1(6205) <= 1929064;
srom_1(6206) <= 1577931;
srom_1(6207) <= 1258737;
srom_1(6208) <= 972976;
srom_1(6209) <= 721990;
srom_1(6210) <= 506955;
srom_1(6211) <= 328880;
srom_1(6212) <= 188600;
srom_1(6213) <= 86773;
srom_1(6214) <= 23876;
srom_1(6215) <= 204;
srom_1(6216) <= 15867;
srom_1(6217) <= 70794;
srom_1(6218) <= 164726;
srom_1(6219) <= 297222;
srom_1(6220) <= 467662;
srom_1(6221) <= 675245;
srom_1(6222) <= 918999;
srom_1(6223) <= 1197781;
srom_1(6224) <= 1510283;
srom_1(6225) <= 1855040;
srom_1(6226) <= 2230435;
srom_1(6227) <= 2634708;
srom_1(6228) <= 3065962;
srom_1(6229) <= 3522177;
srom_1(6230) <= 4001212;
srom_1(6231) <= 4500820;
srom_1(6232) <= 5018660;
srom_1(6233) <= 5552303;
srom_1(6234) <= 6099246;
srom_1(6235) <= 6656925;
srom_1(6236) <= 7222724;
srom_1(6237) <= 7793991;
srom_1(6238) <= 8368046;
srom_1(6239) <= 8942197;
srom_1(6240) <= 9513752;
srom_1(6241) <= 10080031;
srom_1(6242) <= 10638379;
srom_1(6243) <= 11186176;
srom_1(6244) <= 11720855;
srom_1(6245) <= 12239908;
srom_1(6246) <= 12740900;
srom_1(6247) <= 13221483;
srom_1(6248) <= 13679403;
srom_1(6249) <= 14112513;
srom_1(6250) <= 14518782;
srom_1(6251) <= 14896304;
srom_1(6252) <= 15243309;
srom_1(6253) <= 15558170;
srom_1(6254) <= 15839410;
srom_1(6255) <= 16085711;
srom_1(6256) <= 16295918;
srom_1(6257) <= 16469045;
srom_1(6258) <= 16604279;
srom_1(6259) <= 16700988;
srom_1(6260) <= 16758717;
srom_1(6261) <= 16777195;
srom_1(6262) <= 16756337;
srom_1(6263) <= 16696240;
srom_1(6264) <= 16597185;
srom_1(6265) <= 16459637;
srom_1(6266) <= 16284242;
srom_1(6267) <= 16071821;
srom_1(6268) <= 15823371;
srom_1(6269) <= 15540056;
srom_1(6270) <= 15223207;
srom_1(6271) <= 14874307;
srom_1(6272) <= 14494994;
srom_1(6273) <= 14087045;
srom_1(6274) <= 13652375;
srom_1(6275) <= 13193021;
srom_1(6276) <= 12711138;
srom_1(6277) <= 12208985;
srom_1(6278) <= 11688916;
srom_1(6279) <= 11153372;
srom_1(6280) <= 10604862;
srom_1(6281) <= 10045960;
srom_1(6282) <= 9479286;
srom_1(6283) <= 8907497;
srom_1(6284) <= 8333275;
srom_1(6285) <= 7759312;
srom_1(6286) <= 7188301;
srom_1(6287) <= 6622918;
srom_1(6288) <= 6065815;
srom_1(6289) <= 5519604;
srom_1(6290) <= 4986847;
srom_1(6291) <= 4470042;
srom_1(6292) <= 3971613;
srom_1(6293) <= 3493897;
srom_1(6294) <= 3039133;
srom_1(6295) <= 2609455;
srom_1(6296) <= 2206877;
srom_1(6297) <= 1833288;
srom_1(6298) <= 1490438;
srom_1(6299) <= 1179937;
srom_1(6300) <= 903240;
srom_1(6301) <= 661644;
srom_1(6302) <= 456282;
srom_1(6303) <= 288118;
srom_1(6304) <= 157939;
srom_1(6305) <= 66358;
srom_1(6306) <= 13802;
srom_1(6307) <= 518;
srom_1(6308) <= 26569;
srom_1(6309) <= 91833;
srom_1(6310) <= 196003;
srom_1(6311) <= 338590;
srom_1(6312) <= 518928;
srom_1(6313) <= 736168;
srom_1(6314) <= 989294;
srom_1(6315) <= 1277118;
srom_1(6316) <= 1598289;
srom_1(6317) <= 1951303;
srom_1(6318) <= 2334504;
srom_1(6319) <= 2746094;
srom_1(6320) <= 3184145;
srom_1(6321) <= 3646600;
srom_1(6322) <= 4131293;
srom_1(6323) <= 4635949;
srom_1(6324) <= 5158203;
srom_1(6325) <= 5695606;
srom_1(6326) <= 6245637;
srom_1(6327) <= 6805717;
srom_1(6328) <= 7373219;
srom_1(6329) <= 7945484;
srom_1(6330) <= 8519826;
srom_1(6331) <= 9093553;
srom_1(6332) <= 9663974;
srom_1(6333) <= 10228414;
srom_1(6334) <= 10784227;
srom_1(6335) <= 11328806;
srom_1(6336) <= 11859598;
srom_1(6337) <= 12374113;
srom_1(6338) <= 12869938;
srom_1(6339) <= 13344749;
srom_1(6340) <= 13796319;
srom_1(6341) <= 14222530;
srom_1(6342) <= 14621384;
srom_1(6343) <= 14991010;
srom_1(6344) <= 15329676;
srom_1(6345) <= 15635792;
srom_1(6346) <= 15907924;
srom_1(6347) <= 16144795;
srom_1(6348) <= 16345295;
srom_1(6349) <= 16508483;
srom_1(6350) <= 16633594;
srom_1(6351) <= 16720042;
srom_1(6352) <= 16767420;
srom_1(6353) <= 16775508;
srom_1(6354) <= 16744266;
srom_1(6355) <= 16673842;
srom_1(6356) <= 16564566;
srom_1(6357) <= 16416949;
srom_1(6358) <= 16231685;
srom_1(6359) <= 16009642;
srom_1(6360) <= 15751862;
srom_1(6361) <= 15459552;
srom_1(6362) <= 15134085;
srom_1(6363) <= 14776986;
srom_1(6364) <= 14389929;
srom_1(6365) <= 13974730;
srom_1(6366) <= 13533336;
srom_1(6367) <= 13067816;
srom_1(6368) <= 12580354;
srom_1(6369) <= 12073236;
srom_1(6370) <= 11548839;
srom_1(6371) <= 11009622;
srom_1(6372) <= 10458115;
srom_1(6373) <= 9896903;
srom_1(6374) <= 9328618;
srom_1(6375) <= 8755926;
srom_1(6376) <= 8181510;
srom_1(6377) <= 7608066;
srom_1(6378) <= 7038282;
srom_1(6379) <= 6474830;
srom_1(6380) <= 5920353;
srom_1(6381) <= 5377450;
srom_1(6382) <= 4848667;
srom_1(6383) <= 4336484;
srom_1(6384) <= 3843303;
srom_1(6385) <= 3371437;
srom_1(6386) <= 2923098;
srom_1(6387) <= 2500388;
srom_1(6388) <= 2105291;
srom_1(6389) <= 1739658;
srom_1(6390) <= 1405204;
srom_1(6391) <= 1103498;
srom_1(6392) <= 835954;
srom_1(6393) <= 603827;
srom_1(6394) <= 408206;
srom_1(6395) <= 250007;
srom_1(6396) <= 129973;
srom_1(6397) <= 48667;
srom_1(6398) <= 6470;
srom_1(6399) <= 3579;
srom_1(6400) <= 40008;
srom_1(6401) <= 115587;
srom_1(6402) <= 229962;
srom_1(6403) <= 382594;
srom_1(6404) <= 572770;
srom_1(6405) <= 799597;
srom_1(6406) <= 1062011;
srom_1(6407) <= 1358782;
srom_1(6408) <= 1688519;
srom_1(6409) <= 2049674;
srom_1(6410) <= 2440555;
srom_1(6411) <= 2859329;
srom_1(6412) <= 3304031;
srom_1(6413) <= 3772576;
srom_1(6414) <= 4262768;
srom_1(6415) <= 4772307;
srom_1(6416) <= 5298804;
srom_1(6417) <= 5839790;
srom_1(6418) <= 6392728;
srom_1(6419) <= 6955026;
srom_1(6420) <= 7524047;
srom_1(6421) <= 8097121;
srom_1(6422) <= 8671563;
srom_1(6423) <= 9244678;
srom_1(6424) <= 9813778;
srom_1(6425) <= 10376195;
srom_1(6426) <= 10929291;
srom_1(6427) <= 11470474;
srom_1(6428) <= 11997204;
srom_1(6429) <= 12507013;
srom_1(6430) <= 12997509;
srom_1(6431) <= 13466392;
srom_1(6432) <= 13911464;
srom_1(6433) <= 14330637;
srom_1(6434) <= 14721946;
srom_1(6435) <= 15083556;
srom_1(6436) <= 15413771;
srom_1(6437) <= 15711042;
srom_1(6438) <= 15973976;
srom_1(6439) <= 16201340;
srom_1(6440) <= 16392067;
srom_1(6441) <= 16545263;
srom_1(6442) <= 16660209;
srom_1(6443) <= 16736368;
srom_1(6444) <= 16773381;
srom_1(6445) <= 16771074;
srom_1(6446) <= 16729460;
srom_1(6447) <= 16648732;
srom_1(6448) <= 16529270;
srom_1(6449) <= 16371633;
srom_1(6450) <= 16176561;
srom_1(6451) <= 15944969;
srom_1(6452) <= 15677942;
srom_1(6453) <= 15376734;
srom_1(6454) <= 15042755;
srom_1(6455) <= 14677573;
srom_1(6456) <= 14282900;
srom_1(6457) <= 13860586;
srom_1(6458) <= 13412613;
srom_1(6459) <= 12941080;
srom_1(6460) <= 12448199;
srom_1(6461) <= 11936281;
srom_1(6462) <= 11407727;
srom_1(6463) <= 10865015;
srom_1(6464) <= 10310691;
srom_1(6465) <= 9747353;
srom_1(6466) <= 9177643;
srom_1(6467) <= 8604234;
srom_1(6468) <= 8029813;
srom_1(6469) <= 7457075;
srom_1(6470) <= 6888705;
srom_1(6471) <= 6327369;
srom_1(6472) <= 5775698;
srom_1(6473) <= 5236281;
srom_1(6474) <= 4711645;
srom_1(6475) <= 4204253;
srom_1(6476) <= 3716482;
srom_1(6477) <= 3250620;
srom_1(6478) <= 2808852;
srom_1(6479) <= 2393250;
srom_1(6480) <= 2005761;
srom_1(6481) <= 1648204;
srom_1(6482) <= 1322256;
srom_1(6483) <= 1029443;
srom_1(6484) <= 771141;
srom_1(6485) <= 548559;
srom_1(6486) <= 362742;
srom_1(6487) <= 214561;
srom_1(6488) <= 104711;
srom_1(6489) <= 33707;
srom_1(6490) <= 1882;
srom_1(6491) <= 9385;
srom_1(6492) <= 56181;
srom_1(6493) <= 142051;
srom_1(6494) <= 266592;
srom_1(6495) <= 429219;
srom_1(6496) <= 629171;
srom_1(6497) <= 865510;
srom_1(6498) <= 1137127;
srom_1(6499) <= 1442749;
srom_1(6500) <= 1780942;
srom_1(6501) <= 2150121;
srom_1(6502) <= 2548554;
srom_1(6503) <= 2974373;
srom_1(6504) <= 3425581;
srom_1(6505) <= 3900063;
srom_1(6506) <= 4395593;
srom_1(6507) <= 4909848;
srom_1(6508) <= 5440416;
srom_1(6509) <= 5984809;
srom_1(6510) <= 6540474;
srom_1(6511) <= 7104805;
srom_1(6512) <= 7675157;
srom_1(6513) <= 8248855;
srom_1(6514) <= 8823207;
srom_1(6515) <= 9395522;
srom_1(6516) <= 9963115;
srom_1(6517) <= 10523325;
srom_1(6518) <= 11073524;
srom_1(6519) <= 11611133;
srom_1(6520) <= 12133630;
srom_1(6521) <= 12638565;
srom_1(6522) <= 13123571;
srom_1(6523) <= 13586373;
srom_1(6524) <= 14024801;
srom_1(6525) <= 14436799;
srom_1(6526) <= 14820435;
srom_1(6527) <= 15173909;
srom_1(6528) <= 15495566;
srom_1(6529) <= 15783895;
srom_1(6530) <= 16037545;
srom_1(6531) <= 16255327;
srom_1(6532) <= 16436218;
srom_1(6533) <= 16579372;
srom_1(6534) <= 16684117;
srom_1(6535) <= 16749961;
srom_1(6536) <= 16776596;
srom_1(6537) <= 16763896;
srom_1(6538) <= 16711922;
srom_1(6539) <= 16620917;
srom_1(6540) <= 16491308;
srom_1(6541) <= 16323703;
srom_1(6542) <= 16118887;
srom_1(6543) <= 15877822;
srom_1(6544) <= 15601636;
srom_1(6545) <= 15291627;
srom_1(6546) <= 14949247;
srom_1(6547) <= 14576101;
srom_1(6548) <= 14173941;
srom_1(6549) <= 13744651;
srom_1(6550) <= 13290244;
srom_1(6551) <= 12812853;
srom_1(6552) <= 12314714;
srom_1(6553) <= 11798164;
srom_1(6554) <= 11265626;
srom_1(6555) <= 10719597;
srom_1(6556) <= 10162637;
srom_1(6557) <= 9597357;
srom_1(6558) <= 9026410;
srom_1(6559) <= 8452472;
srom_1(6560) <= 7878234;
srom_1(6561) <= 7306389;
srom_1(6562) <= 6739619;
srom_1(6563) <= 6180582;
srom_1(6564) <= 5631900;
srom_1(6565) <= 5096144;
srom_1(6566) <= 4575828;
srom_1(6567) <= 4073391;
srom_1(6568) <= 3591190;
srom_1(6569) <= 3131485;
srom_1(6570) <= 2696433;
srom_1(6571) <= 2288074;
srom_1(6572) <= 1908322;
srom_1(6573) <= 1558958;
srom_1(6574) <= 1241621;
srom_1(6575) <= 957798;
srom_1(6576) <= 708822;
srom_1(6577) <= 495858;
srom_1(6578) <= 319906;
srom_1(6579) <= 181791;
srom_1(6580) <= 82160;
srom_1(6581) <= 21482;
srom_1(6582) <= 40;
srom_1(6583) <= 17934;
srom_1(6584) <= 75082;
srom_1(6585) <= 171214;
srom_1(6586) <= 305881;
srom_1(6587) <= 478450;
srom_1(6588) <= 688113;
srom_1(6589) <= 933886;
srom_1(6590) <= 1214617;
srom_1(6591) <= 1528989;
srom_1(6592) <= 1875528;
srom_1(6593) <= 2252609;
srom_1(6594) <= 2658464;
srom_1(6595) <= 3091190;
srom_1(6596) <= 3548757;
srom_1(6597) <= 4029020;
srom_1(6598) <= 4529726;
srom_1(6599) <= 5048528;
srom_1(6600) <= 5582993;
srom_1(6601) <= 6130614;
srom_1(6602) <= 6688824;
srom_1(6603) <= 7255005;
srom_1(6604) <= 7826501;
srom_1(6605) <= 8400634;
srom_1(6606) <= 8974710;
srom_1(6607) <= 9546037;
srom_1(6608) <= 10111937;
srom_1(6609) <= 10669756;
srom_1(6610) <= 11216877;
srom_1(6611) <= 11750736;
srom_1(6612) <= 12268829;
srom_1(6613) <= 12768726;
srom_1(6614) <= 13248083;
srom_1(6615) <= 13704652;
srom_1(6616) <= 14136293;
srom_1(6617) <= 14540980;
srom_1(6618) <= 14916817;
srom_1(6619) <= 15262042;
srom_1(6620) <= 15575034;
srom_1(6621) <= 15854326;
srom_1(6622) <= 16098609;
srom_1(6623) <= 16306738;
srom_1(6624) <= 16477735;
srom_1(6625) <= 16610800;
srom_1(6626) <= 16705308;
srom_1(6627) <= 16760817;
srom_1(6628) <= 16777065;
srom_1(6629) <= 16753976;
srom_1(6630) <= 16691660;
srom_1(6631) <= 16590408;
srom_1(6632) <= 16450694;
srom_1(6633) <= 16273175;
srom_1(6634) <= 16058683;
srom_1(6635) <= 15808222;
srom_1(6636) <= 15522969;
srom_1(6637) <= 15204260;
srom_1(6638) <= 14853590;
srom_1(6639) <= 14472604;
srom_1(6640) <= 14063088;
srom_1(6641) <= 13626962;
srom_1(6642) <= 13166271;
srom_1(6643) <= 12683177;
srom_1(6644) <= 12179944;
srom_1(6645) <= 11658932;
srom_1(6646) <= 11122584;
srom_1(6647) <= 10573416;
srom_1(6648) <= 10014002;
srom_1(6649) <= 9446966;
srom_1(6650) <= 8874968;
srom_1(6651) <= 8300688;
srom_1(6652) <= 7726821;
srom_1(6653) <= 7156057;
srom_1(6654) <= 6591074;
srom_1(6655) <= 6034519;
srom_1(6656) <= 5489003;
srom_1(6657) <= 4957085;
srom_1(6658) <= 4441258;
srom_1(6659) <= 3943942;
srom_1(6660) <= 3467468;
srom_1(6661) <= 3014072;
srom_1(6662) <= 2585878;
srom_1(6663) <= 2184895;
srom_1(6664) <= 1813004;
srom_1(6665) <= 1471948;
srom_1(6666) <= 1163326;
srom_1(6667) <= 888586;
srom_1(6668) <= 649017;
srom_1(6669) <= 445741;
srom_1(6670) <= 279711;
srom_1(6671) <= 151708;
srom_1(6672) <= 62330;
srom_1(6673) <= 11996;
srom_1(6674) <= 944;
srom_1(6675) <= 29224;
srom_1(6676) <= 96704;
srom_1(6677) <= 203068;
srom_1(6678) <= 347816;
srom_1(6679) <= 530271;
srom_1(6680) <= 749576;
srom_1(6681) <= 1004703;
srom_1(6682) <= 1294455;
srom_1(6683) <= 1617475;
srom_1(6684) <= 1972247;
srom_1(6685) <= 2357107;
srom_1(6686) <= 2770251;
srom_1(6687) <= 3209741;
srom_1(6688) <= 3673517;
srom_1(6689) <= 4159404;
srom_1(6690) <= 4665123;
srom_1(6691) <= 5188302;
srom_1(6692) <= 5726489;
srom_1(6693) <= 6277159;
srom_1(6694) <= 6837731;
srom_1(6695) <= 7405575;
srom_1(6696) <= 7978029;
srom_1(6697) <= 8552409;
srom_1(6698) <= 9126020;
srom_1(6699) <= 9696173;
srom_1(6700) <= 10260195;
srom_1(6701) <= 10815440;
srom_1(6702) <= 11359305;
srom_1(6703) <= 11889239;
srom_1(6704) <= 12402757;
srom_1(6705) <= 12897452;
srom_1(6706) <= 13371004;
srom_1(6707) <= 13821191;
srom_1(6708) <= 14245903;
srom_1(6709) <= 14643148;
srom_1(6710) <= 15011063;
srom_1(6711) <= 15347923;
srom_1(6712) <= 15652149;
srom_1(6713) <= 15922313;
srom_1(6714) <= 16157150;
srom_1(6715) <= 16355557;
srom_1(6716) <= 16516604;
srom_1(6717) <= 16639536;
srom_1(6718) <= 16723777;
srom_1(6719) <= 16768931;
srom_1(6720) <= 16774787;
srom_1(6721) <= 16741318;
srom_1(6722) <= 16668679;
srom_1(6723) <= 16557213;
srom_1(6724) <= 16407441;
srom_1(6725) <= 16220066;
srom_1(6726) <= 15995967;
srom_1(6727) <= 15736194;
srom_1(6728) <= 15441966;
srom_1(6729) <= 15114662;
srom_1(6730) <= 14755817;
srom_1(6731) <= 14367115;
srom_1(6732) <= 13950377;
srom_1(6733) <= 13507558;
srom_1(6734) <= 13040734;
srom_1(6735) <= 12552095;
srom_1(6736) <= 12043932;
srom_1(6737) <= 11518628;
srom_1(6738) <= 10978646;
srom_1(6739) <= 10426519;
srom_1(6740) <= 9864835;
srom_1(6741) <= 9296229;
srom_1(6742) <= 8723366;
srom_1(6743) <= 8148934;
srom_1(6744) <= 7575625;
srom_1(6745) <= 7006129;
srom_1(6746) <= 6443116;
srom_1(6747) <= 5889226;
srom_1(6748) <= 5347056;
srom_1(6749) <= 4819150;
srom_1(6750) <= 4307981;
srom_1(6751) <= 3815948;
srom_1(6752) <= 3345358;
srom_1(6753) <= 2898418;
srom_1(6754) <= 2477222;
srom_1(6755) <= 2083748;
srom_1(6756) <= 1719838;
srom_1(6757) <= 1387201;
srom_1(6758) <= 1087397;
srom_1(6759) <= 821829;
srom_1(6760) <= 591746;
srom_1(6761) <= 398224;
srom_1(6762) <= 242172;
srom_1(6763) <= 124321;
srom_1(6764) <= 45225;
srom_1(6765) <= 5253;
srom_1(6766) <= 4594;
srom_1(6767) <= 43250;
srom_1(6768) <= 121041;
srom_1(6769) <= 237601;
srom_1(6770) <= 392384;
srom_1(6771) <= 584664;
srom_1(6772) <= 813539;
srom_1(6773) <= 1077937;
srom_1(6774) <= 1376616;
srom_1(6775) <= 1708178;
srom_1(6776) <= 2071066;
srom_1(6777) <= 2463579;
srom_1(6778) <= 2883877;
srom_1(6779) <= 3329988;
srom_1(6780) <= 3799821;
srom_1(6781) <= 4291172;
srom_1(6782) <= 4801738;
srom_1(6783) <= 5329124;
srom_1(6784) <= 5870856;
srom_1(6785) <= 6424395;
srom_1(6786) <= 6987145;
srom_1(6787) <= 7556467;
srom_1(6788) <= 8129692;
srom_1(6789) <= 8704130;
srom_1(6790) <= 9277089;
srom_1(6791) <= 9845881;
srom_1(6792) <= 10407840;
srom_1(6793) <= 10960329;
srom_1(6794) <= 11500760;
srom_1(6795) <= 12026596;
srom_1(6796) <= 12535372;
srom_1(6797) <= 13024703;
srom_1(6798) <= 13492293;
srom_1(6799) <= 13935951;
srom_1(6800) <= 14353595;
srom_1(6801) <= 14743267;
srom_1(6802) <= 15103140;
srom_1(6803) <= 15431527;
srom_1(6804) <= 15726886;
srom_1(6805) <= 15987834;
srom_1(6806) <= 16213147;
srom_1(6807) <= 16401767;
srom_1(6808) <= 16552812;
srom_1(6809) <= 16665571;
srom_1(6810) <= 16739517;
srom_1(6811) <= 16774302;
srom_1(6812) <= 16769764;
srom_1(6813) <= 16725924;
srom_1(6814) <= 16642988;
srom_1(6815) <= 16521344;
srom_1(6816) <= 16361562;
srom_1(6817) <= 16164393;
srom_1(6818) <= 15930760;
srom_1(6819) <= 15661760;
srom_1(6820) <= 15358653;
srom_1(6821) <= 15022862;
srom_1(6822) <= 14655960;
srom_1(6823) <= 14259668;
srom_1(6824) <= 13835845;
srom_1(6825) <= 13386478;
srom_1(6826) <= 12913674;
srom_1(6827) <= 12419651;
srom_1(6828) <= 11906724;
srom_1(6829) <= 11377300;
srom_1(6830) <= 10833861;
srom_1(6831) <= 10278955;
srom_1(6832) <= 9715185;
srom_1(6833) <= 9145194;
srom_1(6834) <= 8571655;
srom_1(6835) <= 7997258;
srom_1(6836) <= 7424696;
srom_1(6837) <= 6856654;
srom_1(6838) <= 6295796;
srom_1(6839) <= 5744752;
srom_1(6840) <= 5206105;
srom_1(6841) <= 4682383;
srom_1(6842) <= 4176040;
srom_1(6843) <= 3689452;
srom_1(6844) <= 3224899;
srom_1(6845) <= 2784561;
srom_1(6846) <= 2370502;
srom_1(6847) <= 1984664;
srom_1(6848) <= 1628857;
srom_1(6849) <= 1304748;
srom_1(6850) <= 1013857;
srom_1(6851) <= 757550;
srom_1(6852) <= 537027;
srom_1(6853) <= 353323;
srom_1(6854) <= 207299;
srom_1(6855) <= 99640;
srom_1(6856) <= 30851;
srom_1(6857) <= 1255;
srom_1(6858) <= 10989;
srom_1(6859) <= 60009;
srom_1(6860) <= 148085;
srom_1(6861) <= 274803;
srom_1(6862) <= 439570;
srom_1(6863) <= 641612;
srom_1(6864) <= 879983;
srom_1(6865) <= 1153564;
srom_1(6866) <= 1461073;
srom_1(6867) <= 1801068;
srom_1(6868) <= 2171954;
srom_1(6869) <= 2571991;
srom_1(6870) <= 2999305;
srom_1(6871) <= 3451891;
srom_1(6872) <= 3927627;
srom_1(6873) <= 4424282;
srom_1(6874) <= 4939528;
srom_1(6875) <= 5470947;
srom_1(6876) <= 6016048;
srom_1(6877) <= 6572275;
srom_1(6878) <= 7137019;
srom_1(6879) <= 7707632;
srom_1(6880) <= 8281439;
srom_1(6881) <= 8855748;
srom_1(6882) <= 9427867;
srom_1(6883) <= 9995112;
srom_1(6884) <= 10554824;
srom_1(6885) <= 11104377;
srom_1(6886) <= 11641195;
srom_1(6887) <= 12162761;
srom_1(6888) <= 12666629;
srom_1(6889) <= 13150435;
srom_1(6890) <= 13611912;
srom_1(6891) <= 14048895;
srom_1(6892) <= 14459334;
srom_1(6893) <= 14841306;
srom_1(6894) <= 15193019;
srom_1(6895) <= 15512824;
srom_1(6896) <= 15799221;
srom_1(6897) <= 16050867;
srom_1(6898) <= 16266582;
srom_1(6899) <= 16445355;
srom_1(6900) <= 16586346;
srom_1(6901) <= 16688896;
srom_1(6902) <= 16752522;
srom_1(6903) <= 16776928;
srom_1(6904) <= 16761998;
srom_1(6905) <= 16707802;
srom_1(6906) <= 16614594;
srom_1(6907) <= 16482812;
srom_1(6908) <= 16313073;
srom_1(6909) <= 16106174;
srom_1(6910) <= 15863085;
srom_1(6911) <= 15584945;
srom_1(6912) <= 15273059;
srom_1(6913) <= 14928890;
srom_1(6914) <= 14554050;
srom_1(6915) <= 14150299;
srom_1(6916) <= 13719530;
srom_1(6917) <= 13263762;
srom_1(6918) <= 12785132;
srom_1(6919) <= 12285886;
srom_1(6920) <= 11768364;
srom_1(6921) <= 11234993;
srom_1(6922) <= 10688275;
srom_1(6923) <= 10130773;
srom_1(6924) <= 9565101;
srom_1(6925) <= 8993912;
srom_1(6926) <= 8419884;
srom_1(6927) <= 7845710;
srom_1(6928) <= 7274082;
srom_1(6929) <= 6707680;
srom_1(6930) <= 6149160;
srom_1(6931) <= 5601143;
srom_1(6932) <= 5066196;
srom_1(6933) <= 4546829;
srom_1(6934) <= 4045478;
srom_1(6935) <= 3564493;
srom_1(6936) <= 3106131;
srom_1(6937) <= 2672539;
srom_1(6938) <= 2265752;
srom_1(6939) <= 1887677;
srom_1(6940) <= 1540088;
srom_1(6941) <= 1224613;
srom_1(6942) <= 942733;
srom_1(6943) <= 695769;
srom_1(6944) <= 484879;
srom_1(6945) <= 311053;
srom_1(6946) <= 175105;
srom_1(6947) <= 77673;
srom_1(6948) <= 19214;
srom_1(6949) <= 2;
srom_1(6950) <= 20127;
srom_1(6951) <= 79495;
srom_1(6952) <= 177827;
srom_1(6953) <= 314662;
srom_1(6954) <= 489358;
srom_1(6955) <= 701097;
srom_1(6956) <= 948885;
srom_1(6957) <= 1231561;
srom_1(6958) <= 1547798;
srom_1(6959) <= 1896115;
srom_1(6960) <= 2274876;
srom_1(6961) <= 2682308;
srom_1(6962) <= 3116498;
srom_1(6963) <= 3575410;
srom_1(6964) <= 4056894;
srom_1(6965) <= 4558690;
srom_1(6966) <= 5078447;
srom_1(6967) <= 5613725;
srom_1(6968) <= 6162016;
srom_1(6969) <= 6720749;
srom_1(6970) <= 7287302;
srom_1(6971) <= 7859020;
srom_1(6972) <= 8433221;
srom_1(6973) <= 9007213;
srom_1(6974) <= 9578304;
srom_1(6975) <= 10143817;
srom_1(6976) <= 10701098;
srom_1(6977) <= 11247536;
srom_1(6978) <= 11780567;
srom_1(6979) <= 12297691;
srom_1(6980) <= 12796485;
srom_1(6981) <= 13274609;
srom_1(6982) <= 13729821;
srom_1(6983) <= 14159985;
srom_1(6984) <= 14563086;
srom_1(6985) <= 14937233;
srom_1(6986) <= 15280671;
srom_1(6987) <= 15591789;
srom_1(6988) <= 15869130;
srom_1(6989) <= 16111391;
srom_1(6990) <= 16317438;
srom_1(6991) <= 16486304;
srom_1(6992) <= 16617197;
srom_1(6993) <= 16709503;
srom_1(6994) <= 16762790;
srom_1(6995) <= 16776807;
srom_1(6996) <= 16751489;
srom_1(6997) <= 16686955;
srom_1(6998) <= 16583507;
srom_1(6999) <= 16441630;
srom_1(7000) <= 16261990;
srom_1(7001) <= 16045429;
srom_1(7002) <= 15792962;
srom_1(7003) <= 15505774;
srom_1(7004) <= 15185211;
srom_1(7005) <= 14832776;
srom_1(7006) <= 14450122;
srom_1(7007) <= 14039044;
srom_1(7008) <= 13601469;
srom_1(7009) <= 13139449;
srom_1(7010) <= 12655151;
srom_1(7011) <= 12150846;
srom_1(7012) <= 11628898;
srom_1(7013) <= 11091755;
srom_1(7014) <= 10541936;
srom_1(7015) <= 9982020;
srom_1(7016) <= 9414631;
srom_1(7017) <= 8842431;
srom_1(7018) <= 8268103;
srom_1(7019) <= 7694340;
srom_1(7020) <= 7123833;
srom_1(7021) <= 6559256;
srom_1(7022) <= 6003258;
srom_1(7023) <= 5458446;
srom_1(7024) <= 4927375;
srom_1(7025) <= 4412534;
srom_1(7026) <= 3916338;
srom_1(7027) <= 3441115;
srom_1(7028) <= 2989091;
srom_1(7029) <= 2562388;
srom_1(7030) <= 2163007;
srom_1(7031) <= 1792819;
srom_1(7032) <= 1453561;
srom_1(7033) <= 1146824;
srom_1(7034) <= 874046;
srom_1(7035) <= 636506;
srom_1(7036) <= 435319;
srom_1(7037) <= 271428;
srom_1(7038) <= 145600;
srom_1(7039) <= 58427;
srom_1(7040) <= 10317;
srom_1(7041) <= 1496;
srom_1(7042) <= 32005;
srom_1(7043) <= 101700;
srom_1(7044) <= 210256;
srom_1(7045) <= 357163;
srom_1(7046) <= 541732;
srom_1(7047) <= 763098;
srom_1(7048) <= 1020223;
srom_1(7049) <= 1311900;
srom_1(7050) <= 1636763;
srom_1(7051) <= 1993287;
srom_1(7052) <= 2379801;
srom_1(7053) <= 2794492;
srom_1(7054) <= 3235416;
srom_1(7055) <= 3700506;
srom_1(7056) <= 4187579;
srom_1(7057) <= 4694352;
srom_1(7058) <= 5218449;
srom_1(7059) <= 5757412;
srom_1(7060) <= 6308714;
srom_1(7061) <= 6869769;
srom_1(7062) <= 7437946;
srom_1(7063) <= 8010581;
srom_1(7064) <= 8584989;
srom_1(7065) <= 9158476;
srom_1(7066) <= 9728353;
srom_1(7067) <= 10291947;
srom_1(7068) <= 10846616;
srom_1(7069) <= 11389758;
srom_1(7070) <= 11918827;
srom_1(7071) <= 12431342;
srom_1(7072) <= 12924898;
srom_1(7073) <= 13397183;
srom_1(7074) <= 13845981;
srom_1(7075) <= 14269187;
srom_1(7076) <= 14664817;
srom_1(7077) <= 15031015;
srom_1(7078) <= 15366066;
srom_1(7079) <= 15668396;
srom_1(7080) <= 15936589;
srom_1(7081) <= 16169387;
srom_1(7082) <= 16365698;
srom_1(7083) <= 16524602;
srom_1(7084) <= 16645354;
srom_1(7085) <= 16727386;
srom_1(7086) <= 16770316;
srom_1(7087) <= 16773940;
srom_1(7088) <= 16738243;
srom_1(7089) <= 16663392;
srom_1(7090) <= 16549737;
srom_1(7091) <= 16397812;
srom_1(7092) <= 16208329;
srom_1(7093) <= 15982176;
srom_1(7094) <= 15720415;
srom_1(7095) <= 15424273;
srom_1(7096) <= 15095137;
srom_1(7097) <= 14734553;
srom_1(7098) <= 14344210;
srom_1(7099) <= 13925939;
srom_1(7100) <= 13481702;
srom_1(7101) <= 13013582;
srom_1(7102) <= 12523773;
srom_1(7103) <= 12014574;
srom_1(7104) <= 11488370;
srom_1(7105) <= 10947631;
srom_1(7106) <= 10394892;
srom_1(7107) <= 9832745;
srom_1(7108) <= 9263826;
srom_1(7109) <= 8690802;
srom_1(7110) <= 8116361;
srom_1(7111) <= 7543197;
srom_1(7112) <= 6973998;
srom_1(7113) <= 6411432;
srom_1(7114) <= 5858137;
srom_1(7115) <= 5316709;
srom_1(7116) <= 4789686;
srom_1(7117) <= 4279540;
srom_1(7118) <= 3788662;
srom_1(7119) <= 3319355;
srom_1(7120) <= 2873820;
srom_1(7121) <= 2454145;
srom_1(7122) <= 2062300;
srom_1(7123) <= 1700120;
srom_1(7124) <= 1369305;
srom_1(7125) <= 1071406;
srom_1(7126) <= 807819;
srom_1(7127) <= 579782;
srom_1(7128) <= 388363;
srom_1(7129) <= 234460;
srom_1(7130) <= 118794;
srom_1(7131) <= 41908;
srom_1(7132) <= 4163;
srom_1(7133) <= 5736;
srom_1(7134) <= 46618;
srom_1(7135) <= 126619;
srom_1(7136) <= 245364;
srom_1(7137) <= 402295;
srom_1(7138) <= 596676;
srom_1(7139) <= 827596;
srom_1(7140) <= 1093973;
srom_1(7141) <= 1394556;
srom_1(7142) <= 1727938;
srom_1(7143) <= 2092553;
srom_1(7144) <= 2486693;
srom_1(7145) <= 2908508;
srom_1(7146) <= 3356022;
srom_1(7147) <= 3827135;
srom_1(7148) <= 4319639;
srom_1(7149) <= 4831224;
srom_1(7150) <= 5359490;
srom_1(7151) <= 5901961;
srom_1(7152) <= 6456092;
srom_1(7153) <= 7019286;
srom_1(7154) <= 7588901;
srom_1(7155) <= 8162266;
srom_1(7156) <= 8736692;
srom_1(7157) <= 9309486;
srom_1(7158) <= 9877962;
srom_1(7159) <= 10439454;
srom_1(7160) <= 10991329;
srom_1(7161) <= 11530998;
srom_1(7162) <= 12055932;
srom_1(7163) <= 12563668;
srom_1(7164) <= 13051826;
srom_1(7165) <= 13518117;
srom_1(7166) <= 13960354;
srom_1(7167) <= 14376463;
srom_1(7168) <= 14764492;
srom_1(7169) <= 15122623;
srom_1(7170) <= 15449176;
srom_1(7171) <= 15742620;
srom_1(7172) <= 16001578;
srom_1(7173) <= 16224836;
srom_1(7174) <= 16411347;
srom_1(7175) <= 16560237;
srom_1(7176) <= 16670807;
srom_1(7177) <= 16742540;
srom_1(7178) <= 16775097;
srom_1(7179) <= 16768328;
srom_1(7180) <= 16722263;
srom_1(7181) <= 16637119;
srom_1(7182) <= 16513295;
srom_1(7183) <= 16351371;
srom_1(7184) <= 16152108;
srom_1(7185) <= 15916438;
srom_1(7186) <= 15645468;
srom_1(7187) <= 15340468;
srom_1(7188) <= 15002868;
srom_1(7189) <= 14634252;
srom_1(7190) <= 14236348;
srom_1(7191) <= 13811021;
srom_1(7192) <= 13360268;
srom_1(7193) <= 12886200;
srom_1(7194) <= 12391041;
srom_1(7195) <= 11877114;
srom_1(7196) <= 11346828;
srom_1(7197) <= 10802670;
srom_1(7198) <= 10247191;
srom_1(7199) <= 9682997;
srom_1(7200) <= 9112733;
srom_1(7201) <= 8539074;
srom_1(7202) <= 7964709;
srom_1(7203) <= 7392331;
srom_1(7204) <= 6824626;
srom_1(7205) <= 6264254;
srom_1(7206) <= 5713845;
srom_1(7207) <= 5175978;
srom_1(7208) <= 4653176;
srom_1(7209) <= 4147891;
srom_1(7210) <= 3662492;
srom_1(7211) <= 3199256;
srom_1(7212) <= 2760354;
srom_1(7213) <= 2347845;
srom_1(7214) <= 1963664;
srom_1(7215) <= 1609611;
srom_1(7216) <= 1287347;
srom_1(7217) <= 998383;
srom_1(7218) <= 744075;
srom_1(7219) <= 525614;
srom_1(7220) <= 344026;
srom_1(7221) <= 200161;
srom_1(7222) <= 94695;
srom_1(7223) <= 28122;
srom_1(7224) <= 754;
srom_1(7225) <= 12720;
srom_1(7226) <= 63963;
srom_1(7227) <= 154243;
srom_1(7228) <= 283137;
srom_1(7229) <= 450040;
srom_1(7230) <= 654170;
srom_1(7231) <= 894570;
srom_1(7232) <= 1170111;
srom_1(7233) <= 1479503;
srom_1(7234) <= 1821293;
srom_1(7235) <= 2193880;
srom_1(7236) <= 2595517;
srom_1(7237) <= 3024319;
srom_1(7238) <= 3478276;
srom_1(7239) <= 3955259;
srom_1(7240) <= 4453031;
srom_1(7241) <= 4969259;
srom_1(7242) <= 5501522;
srom_1(7243) <= 6047323;
srom_1(7244) <= 6604103;
srom_1(7245) <= 7169251;
srom_1(7246) <= 7740118;
srom_1(7247) <= 8314025;
srom_1(7248) <= 8888282;
srom_1(7249) <= 9460196;
srom_1(7250) <= 10027084;
srom_1(7251) <= 10586290;
srom_1(7252) <= 11135189;
srom_1(7253) <= 11671209;
srom_1(7254) <= 12191836;
srom_1(7255) <= 12694628;
srom_1(7256) <= 13177228;
srom_1(7257) <= 13637372;
srom_1(7258) <= 14072903;
srom_1(7259) <= 14481778;
srom_1(7260) <= 14862081;
srom_1(7261) <= 15212027;
srom_1(7262) <= 15529975;
srom_1(7263) <= 15814436;
srom_1(7264) <= 16064074;
srom_1(7265) <= 16277719;
srom_1(7266) <= 16454369;
srom_1(7267) <= 16593196;
srom_1(7268) <= 16693549;
srom_1(7269) <= 16754958;
srom_1(7270) <= 16777133;
srom_1(7271) <= 16759972;
srom_1(7272) <= 16703555;
srom_1(7273) <= 16608146;
srom_1(7274) <= 16474193;
srom_1(7275) <= 16302324;
srom_1(7276) <= 16093345;
srom_1(7277) <= 15848235;
srom_1(7278) <= 15568145;
srom_1(7279) <= 15254387;
srom_1(7280) <= 14908434;
srom_1(7281) <= 14531906;
srom_1(7282) <= 14126571;
srom_1(7283) <= 13694328;
srom_1(7284) <= 13237205;
srom_1(7285) <= 12757346;
srom_1(7286) <= 12256999;
srom_1(7287) <= 11738513;
srom_1(7288) <= 11204318;
srom_1(7289) <= 10656918;
srom_1(7290) <= 10098882;
srom_1(7291) <= 9532826;
srom_1(7292) <= 8961404;
srom_1(7293) <= 8387297;
srom_1(7294) <= 7813195;
srom_1(7295) <= 7241791;
srom_1(7296) <= 6675766;
srom_1(7297) <= 6117772;
srom_1(7298) <= 5570428;
srom_1(7299) <= 5036298;
srom_1(7300) <= 4517889;
srom_1(7301) <= 4017631;
srom_1(7302) <= 3537870;
srom_1(7303) <= 3080856;
srom_1(7304) <= 2648731;
srom_1(7305) <= 2243523;
srom_1(7306) <= 1867131;
srom_1(7307) <= 1521321;
srom_1(7308) <= 1207713;
srom_1(7309) <= 927780;
srom_1(7310) <= 682833;
srom_1(7311) <= 474020;
srom_1(7312) <= 302322;
srom_1(7313) <= 168544;
srom_1(7314) <= 73312;
srom_1(7315) <= 17073;
srom_1(7316) <= 91;
srom_1(7317) <= 22446;
srom_1(7318) <= 84033;
srom_1(7319) <= 184563;
srom_1(7320) <= 323564;
srom_1(7321) <= 500385;
srom_1(7322) <= 714197;
srom_1(7323) <= 963997;
srom_1(7324) <= 1248613;
srom_1(7325) <= 1566711;
srom_1(7326) <= 1916799;
srom_1(7327) <= 2297236;
srom_1(7328) <= 2706237;
srom_1(7329) <= 3141885;
srom_1(7330) <= 3602137;
srom_1(7331) <= 4084834;
srom_1(7332) <= 4587712;
srom_1(7333) <= 5108415;
srom_1(7334) <= 5644499;
srom_1(7335) <= 6193452;
srom_1(7336) <= 6752698;
srom_1(7337) <= 7319616;
srom_1(7338) <= 7891547;
srom_1(7339) <= 8465808;
srom_1(7340) <= 9039708;
srom_1(7341) <= 9610554;
srom_1(7342) <= 10175670;
srom_1(7343) <= 10732406;
srom_1(7344) <= 11278151;
srom_1(7345) <= 11810346;
srom_1(7346) <= 12326495;
srom_1(7347) <= 12824178;
srom_1(7348) <= 13301061;
srom_1(7349) <= 13754908;
srom_1(7350) <= 14183591;
srom_1(7351) <= 14585099;
srom_1(7352) <= 14957550;
srom_1(7353) <= 15299196;
srom_1(7354) <= 15608436;
srom_1(7355) <= 15883820;
srom_1(7356) <= 16124057;
srom_1(7357) <= 16328019;
srom_1(7358) <= 16494750;
srom_1(7359) <= 16623470;
srom_1(7360) <= 16713573;
srom_1(7361) <= 16764637;
srom_1(7362) <= 16776423;
srom_1(7363) <= 16748876;
srom_1(7364) <= 16682125;
srom_1(7365) <= 16576482;
srom_1(7366) <= 16432444;
srom_1(7367) <= 16250686;
srom_1(7368) <= 16032059;
srom_1(7369) <= 15777590;
srom_1(7370) <= 15488471;
srom_1(7371) <= 15166059;
srom_1(7372) <= 14811865;
srom_1(7373) <= 14427550;
srom_1(7374) <= 14014916;
srom_1(7375) <= 13575898;
srom_1(7376) <= 13112556;
srom_1(7377) <= 12627061;
srom_1(7378) <= 12121691;
srom_1(7379) <= 11598815;
srom_1(7380) <= 11060885;
srom_1(7381) <= 10510424;
srom_1(7382) <= 9950013;
srom_1(7383) <= 9382280;
srom_1(7384) <= 8809888;
srom_1(7385) <= 8235520;
srom_1(7386) <= 7661869;
srom_1(7387) <= 7091627;
srom_1(7388) <= 6527467;
srom_1(7389) <= 5972034;
srom_1(7390) <= 5427933;
srom_1(7391) <= 4897716;
srom_1(7392) <= 4383869;
srom_1(7393) <= 3888802;
srom_1(7394) <= 3414835;
srom_1(7395) <= 2964193;
srom_1(7396) <= 2538987;
srom_1(7397) <= 2141212;
srom_1(7398) <= 1772734;
srom_1(7399) <= 1435279;
srom_1(7400) <= 1130431;
srom_1(7401) <= 859619;
srom_1(7402) <= 624113;
srom_1(7403) <= 425018;
srom_1(7404) <= 263266;
srom_1(7405) <= 139617;
srom_1(7406) <= 54651;
srom_1(7407) <= 8765;
srom_1(7408) <= 2175;
srom_1(7409) <= 34912;
srom_1(7410) <= 106822;
srom_1(7411) <= 217568;
srom_1(7412) <= 366632;
srom_1(7413) <= 553313;
srom_1(7414) <= 776736;
srom_1(7415) <= 1035854;
srom_1(7416) <= 1329452;
srom_1(7417) <= 1656152;
srom_1(7418) <= 2014424;
srom_1(7419) <= 2402585;
srom_1(7420) <= 2818818;
srom_1(7421) <= 3261169;
srom_1(7422) <= 3727565;
srom_1(7423) <= 4215817;
srom_1(7424) <= 4723638;
srom_1(7425) <= 5248644;
srom_1(7426) <= 5788375;
srom_1(7427) <= 6340300;
srom_1(7428) <= 6901829;
srom_1(7429) <= 7470331;
srom_1(7430) <= 8043138;
srom_1(7431) <= 8617566;
srom_1(7432) <= 9190920;
srom_1(7433) <= 9760512;
srom_1(7434) <= 10323670;
srom_1(7435) <= 10877755;
srom_1(7436) <= 11420166;
srom_1(7437) <= 11948362;
srom_1(7438) <= 12459865;
srom_1(7439) <= 12952276;
srom_1(7440) <= 13423287;
srom_1(7441) <= 13870688;
srom_1(7442) <= 14292382;
srom_1(7443) <= 14686391;
srom_1(7444) <= 15050868;
srom_1(7445) <= 15384103;
srom_1(7446) <= 15684533;
srom_1(7447) <= 15950751;
srom_1(7448) <= 16181507;
srom_1(7449) <= 16375720;
srom_1(7450) <= 16532478;
srom_1(7451) <= 16651047;
srom_1(7452) <= 16730870;
srom_1(7453) <= 16771574;
srom_1(7454) <= 16772967;
srom_1(7455) <= 16735043;
srom_1(7456) <= 16657979;
srom_1(7457) <= 16542138;
srom_1(7458) <= 16388062;
srom_1(7459) <= 16196474;
srom_1(7460) <= 15968272;
srom_1(7461) <= 15704526;
srom_1(7462) <= 15406473;
srom_1(7463) <= 15075512;
srom_1(7464) <= 14713193;
srom_1(7465) <= 14321216;
srom_1(7466) <= 13901418;
srom_1(7467) <= 13455770;
srom_1(7468) <= 12986360;
srom_1(7469) <= 12495389;
srom_1(7470) <= 11985160;
srom_1(7471) <= 11458066;
srom_1(7472) <= 10916578;
srom_1(7473) <= 10363235;
srom_1(7474) <= 9800633;
srom_1(7475) <= 9231409;
srom_1(7476) <= 8658233;
srom_1(7477) <= 8083793;
srom_1(7478) <= 7510782;
srom_1(7479) <= 6941887;
srom_1(7480) <= 6379777;
srom_1(7481) <= 5827087;
srom_1(7482) <= 5286408;
srom_1(7483) <= 4760277;
srom_1(7484) <= 4251160;
srom_1(7485) <= 3761446;
srom_1(7486) <= 3293429;
srom_1(7487) <= 2849306;
srom_1(7488) <= 2431158;
srom_1(7489) <= 2040947;
srom_1(7490) <= 1680502;
srom_1(7491) <= 1351514;
srom_1(7492) <= 1055525;
srom_1(7493) <= 793924;
srom_1(7494) <= 567936;
srom_1(7495) <= 378622;
srom_1(7496) <= 226870;
srom_1(7497) <= 113392;
srom_1(7498) <= 38718;
srom_1(7499) <= 3200;
srom_1(7500) <= 7004;
srom_1(7501) <= 50112;
srom_1(7502) <= 132322;
srom_1(7503) <= 253249;
srom_1(7504) <= 412325;
srom_1(7505) <= 608805;
srom_1(7506) <= 841767;
srom_1(7507) <= 1110119;
srom_1(7508) <= 1412602;
srom_1(7509) <= 1747798;
srom_1(7510) <= 2114135;
srom_1(7511) <= 2509895;
srom_1(7512) <= 2933222;
srom_1(7513) <= 3382132;
srom_1(7514) <= 3854519;
srom_1(7515) <= 4348167;
srom_1(7516) <= 4860763;
srom_1(7517) <= 5389902;
srom_1(7518) <= 5933102;
srom_1(7519) <= 6487818;
srom_1(7520) <= 7051447;
srom_1(7521) <= 7621346;
srom_1(7522) <= 8194843;
srom_1(7523) <= 8769249;
srom_1(7524) <= 9341870;
srom_1(7525) <= 9910021;
srom_1(7526) <= 10471037;
srom_1(7527) <= 11022288;
srom_1(7528) <= 11561189;
srom_1(7529) <= 12085213;
srom_1(7530) <= 12591902;
srom_1(7531) <= 13078880;
srom_1(7532) <= 13543864;
srom_1(7533) <= 13984673;
srom_1(7534) <= 14399240;
srom_1(7535) <= 14785621;
srom_1(7536) <= 15142005;
srom_1(7537) <= 15466719;
srom_1(7538) <= 15758242;
srom_1(7539) <= 16015206;
srom_1(7540) <= 16236406;
srom_1(7541) <= 16420806;
srom_1(7542) <= 16567539;
srom_1(7543) <= 16675919;
srom_1(7544) <= 16745437;
srom_1(7545) <= 16775766;
srom_1(7546) <= 16766765;
srom_1(7547) <= 16718477;
srom_1(7548) <= 16631126;
srom_1(7549) <= 16505124;
srom_1(7550) <= 16341060;
srom_1(7551) <= 16139705;
srom_1(7552) <= 15902002;
srom_1(7553) <= 15629066;
srom_1(7554) <= 15322178;
srom_1(7555) <= 14982775;
srom_1(7556) <= 14612450;
srom_1(7557) <= 14212939;
srom_1(7558) <= 13786116;
srom_1(7559) <= 13333982;
srom_1(7560) <= 12858658;
srom_1(7561) <= 12362372;
srom_1(7562) <= 11847452;
srom_1(7563) <= 11316312;
srom_1(7564) <= 10771443;
srom_1(7565) <= 10215400;
srom_1(7566) <= 9650790;
srom_1(7567) <= 9080262;
srom_1(7568) <= 8506490;
srom_1(7569) <= 7932166;
srom_1(7570) <= 7359982;
srom_1(7571) <= 6792621;
srom_1(7572) <= 6232745;
srom_1(7573) <= 5682978;
srom_1(7574) <= 5145899;
srom_1(7575) <= 4624026;
srom_1(7576) <= 4119806;
srom_1(7577) <= 3635605;
srom_1(7578) <= 3173691;
srom_1(7579) <= 2736233;
srom_1(7580) <= 2325280;
srom_1(7581) <= 1942760;
srom_1(7582) <= 1590467;
srom_1(7583) <= 1270053;
srom_1(7584) <= 983020;
srom_1(7585) <= 730714;
srom_1(7586) <= 514319;
srom_1(7587) <= 334850;
srom_1(7588) <= 193147;
srom_1(7589) <= 89875;
srom_1(7590) <= 25519;
srom_1(7591) <= 380;
srom_1(7592) <= 14577;
srom_1(7593) <= 68042;
srom_1(7594) <= 160526;
srom_1(7595) <= 291593;
srom_1(7596) <= 460631;
srom_1(7597) <= 666845;
srom_1(7598) <= 909269;
srom_1(7599) <= 1186767;
srom_1(7600) <= 1498036;
srom_1(7601) <= 1841618;
srom_1(7602) <= 2215901;
srom_1(7603) <= 2619129;
srom_1(7604) <= 3049413;
srom_1(7605) <= 3504734;
srom_1(7606) <= 3982957;
srom_1(7607) <= 4481840;
srom_1(7608) <= 4999043;
srom_1(7609) <= 5532141;
srom_1(7610) <= 6078633;
srom_1(7611) <= 6635958;
srom_1(7612) <= 7201502;
srom_1(7613) <= 7772613;
srom_1(7614) <= 8346612;
srom_1(7615) <= 8920808;
srom_1(7616) <= 9492508;
srom_1(7617) <= 10059032;
srom_1(7618) <= 10617723;
srom_1(7619) <= 11165960;
srom_1(7620) <= 11701174;
srom_1(7621) <= 12220853;
srom_1(7622) <= 12722562;
srom_1(7623) <= 13203948;
srom_1(7624) <= 13662753;
srom_1(7625) <= 14096825;
srom_1(7626) <= 14504130;
srom_1(7627) <= 14882757;
srom_1(7628) <= 15230931;
srom_1(7629) <= 15547019;
srom_1(7630) <= 15829538;
srom_1(7631) <= 16077164;
srom_1(7632) <= 16288736;
srom_1(7633) <= 16463262;
srom_1(7634) <= 16599923;
srom_1(7635) <= 16698078;
srom_1(7636) <= 16757267;
srom_1(7637) <= 16777213;
srom_1(7638) <= 16757821;
srom_1(7639) <= 16699183;
srom_1(7640) <= 16601575;
srom_1(7641) <= 16465453;
srom_1(7642) <= 16291455;
srom_1(7643) <= 16080399;
srom_1(7644) <= 15833273;
srom_1(7645) <= 15551237;
srom_1(7646) <= 15235612;
srom_1(7647) <= 14887880;
srom_1(7648) <= 14509670;
srom_1(7649) <= 14102756;
srom_1(7650) <= 13669047;
srom_1(7651) <= 13210576;
srom_1(7652) <= 12729493;
srom_1(7653) <= 12228054;
srom_1(7654) <= 11708611;
srom_1(7655) <= 11173599;
srom_1(7656) <= 10625527;
srom_1(7657) <= 10066966;
srom_1(7658) <= 9500534;
srom_1(7659) <= 8928888;
srom_1(7660) <= 8354709;
srom_1(7661) <= 7780688;
srom_1(7662) <= 7209518;
srom_1(7663) <= 6643878;
srom_1(7664) <= 6086418;
srom_1(7665) <= 5539755;
srom_1(7666) <= 5006451;
srom_1(7667) <= 4489007;
srom_1(7668) <= 3989850;
srom_1(7669) <= 3511319;
srom_1(7670) <= 3055661;
srom_1(7671) <= 2625010;
srom_1(7672) <= 2221386;
srom_1(7673) <= 1846683;
srom_1(7674) <= 1502657;
srom_1(7675) <= 1190922;
srom_1(7676) <= 912939;
srom_1(7677) <= 670012;
srom_1(7678) <= 463281;
srom_1(7679) <= 293713;
srom_1(7680) <= 162106;
srom_1(7681) <= 69076;
srom_1(7682) <= 15058;
srom_1(7683) <= 307;
srom_1(7684) <= 24892;
srom_1(7685) <= 88697;
srom_1(7686) <= 191423;
srom_1(7687) <= 332588;
srom_1(7688) <= 511531;
srom_1(7689) <= 727413;
srom_1(7690) <= 979220;
srom_1(7691) <= 1265772;
srom_1(7692) <= 1585726;
srom_1(7693) <= 1937581;
srom_1(7694) <= 2319687;
srom_1(7695) <= 2730252;
srom_1(7696) <= 3167351;
srom_1(7697) <= 3628935;
srom_1(7698) <= 4112838;
srom_1(7699) <= 4616792;
srom_1(7700) <= 5138433;
srom_1(7701) <= 5675315;
srom_1(7702) <= 6224921;
srom_1(7703) <= 6784673;
srom_1(7704) <= 7351946;
srom_1(7705) <= 7924081;
srom_1(7706) <= 8498394;
srom_1(7707) <= 9072192;
srom_1(7708) <= 9642785;
srom_1(7709) <= 10207496;
srom_1(7710) <= 10763678;
srom_1(7711) <= 11308722;
srom_1(7712) <= 11840073;
srom_1(7713) <= 12355239;
srom_1(7714) <= 12851804;
srom_1(7715) <= 13327440;
srom_1(7716) <= 13779915;
srom_1(7717) <= 14207109;
srom_1(7718) <= 14607018;
srom_1(7719) <= 14977767;
srom_1(7720) <= 15317617;
srom_1(7721) <= 15624974;
srom_1(7722) <= 15898398;
srom_1(7723) <= 16136605;
srom_1(7724) <= 16338480;
srom_1(7725) <= 16503075;
srom_1(7726) <= 16629618;
srom_1(7727) <= 16717516;
srom_1(7728) <= 16766357;
srom_1(7729) <= 16775913;
srom_1(7730) <= 16746137;
srom_1(7731) <= 16677170;
srom_1(7732) <= 16569334;
srom_1(7733) <= 16423137;
srom_1(7734) <= 16239263;
srom_1(7735) <= 16018575;
srom_1(7736) <= 15762107;
srom_1(7737) <= 15471062;
srom_1(7738) <= 15146805;
srom_1(7739) <= 14790856;
srom_1(7740) <= 14404885;
srom_1(7741) <= 13990702;
srom_1(7742) <= 13550249;
srom_1(7743) <= 13085591;
srom_1(7744) <= 12598907;
srom_1(7745) <= 12092480;
srom_1(7746) <= 11568683;
srom_1(7747) <= 11029975;
srom_1(7748) <= 10478880;
srom_1(7749) <= 9917983;
srom_1(7750) <= 9349914;
srom_1(7751) <= 8777338;
srom_1(7752) <= 8202938;
srom_1(7753) <= 7629410;
srom_1(7754) <= 7059441;
srom_1(7755) <= 6495705;
srom_1(7756) <= 5940846;
srom_1(7757) <= 5397465;
srom_1(7758) <= 4868111;
srom_1(7759) <= 4355265;
srom_1(7760) <= 3861333;
srom_1(7761) <= 3388631;
srom_1(7762) <= 2939376;
srom_1(7763) <= 2515674;
srom_1(7764) <= 2119512;
srom_1(7765) <= 1752748;
srom_1(7766) <= 1417102;
srom_1(7767) <= 1114148;
srom_1(7768) <= 845306;
srom_1(7769) <= 611837;
srom_1(7770) <= 414837;
srom_1(7771) <= 255228;
srom_1(7772) <= 133759;
srom_1(7773) <= 51000;
srom_1(7774) <= 7339;
srom_1(7775) <= 2980;
srom_1(7776) <= 37945;
srom_1(7777) <= 112069;
srom_1(7778) <= 225004;
srom_1(7779) <= 376221;
srom_1(7780) <= 565011;
srom_1(7781) <= 790489;
srom_1(7782) <= 1051596;
srom_1(7783) <= 1347110;
srom_1(7784) <= 1675643;
srom_1(7785) <= 2035656;
srom_1(7786) <= 2425460;
srom_1(7787) <= 2843228;
srom_1(7788) <= 3286999;
srom_1(7789) <= 3754694;
srom_1(7790) <= 4244119;
srom_1(7791) <= 4752978;
srom_1(7792) <= 5278887;
srom_1(7793) <= 5819378;
srom_1(7794) <= 6371916;
srom_1(7795) <= 6933912;
srom_1(7796) <= 7502730;
srom_1(7797) <= 8075701;
srom_1(7798) <= 8650140;
srom_1(7799) <= 9223353;
srom_1(7800) <= 9792651;
srom_1(7801) <= 10355365;
srom_1(7802) <= 10908856;
srom_1(7803) <= 11450529;
srom_1(7804) <= 11977843;
srom_1(7805) <= 12488327;
srom_1(7806) <= 12979585;
srom_1(7807) <= 13449315;
srom_1(7808) <= 13895313;
srom_1(7809) <= 14315488;
srom_1(7810) <= 14707870;
srom_1(7811) <= 15070619;
srom_1(7812) <= 15402034;
srom_1(7813) <= 15700561;
srom_1(7814) <= 15964799;
srom_1(7815) <= 16193510;
srom_1(7816) <= 16385620;
srom_1(7817) <= 16540231;
srom_1(7818) <= 16656615;
srom_1(7819) <= 16734228;
srom_1(7820) <= 16772705;
srom_1(7821) <= 16771867;
srom_1(7822) <= 16731716;
srom_1(7823) <= 16652442;
srom_1(7824) <= 16534416;
srom_1(7825) <= 16378191;
srom_1(7826) <= 16184500;
srom_1(7827) <= 15954252;
srom_1(7828) <= 15688526;
srom_1(7829) <= 15388568;
srom_1(7830) <= 15055785;
srom_1(7831) <= 14691737;
srom_1(7832) <= 14298132;
srom_1(7833) <= 13876814;
srom_1(7834) <= 13429761;
srom_1(7835) <= 12959068;
srom_1(7836) <= 12466942;
srom_1(7837) <= 11955692;
srom_1(7838) <= 11427715;
srom_1(7839) <= 10885486;
srom_1(7840) <= 10331548;
srom_1(7841) <= 9768499;
srom_1(7842) <= 9198980;
srom_1(7843) <= 8625660;
srom_1(7844) <= 8051229;
srom_1(7845) <= 7478380;
srom_1(7846) <= 6909799;
srom_1(7847) <= 6348153;
srom_1(7848) <= 5796075;
srom_1(7849) <= 5256154;
srom_1(7850) <= 4730923;
srom_1(7851) <= 4222843;
srom_1(7852) <= 3734299;
srom_1(7853) <= 3267580;
srom_1(7854) <= 2824875;
srom_1(7855) <= 2408261;
srom_1(7856) <= 2019690;
srom_1(7857) <= 1660986;
srom_1(7858) <= 1333829;
srom_1(7859) <= 1039755;
srom_1(7860) <= 780142;
srom_1(7861) <= 556208;
srom_1(7862) <= 369003;
srom_1(7863) <= 219404;
srom_1(7864) <= 108114;
srom_1(7865) <= 35654;
srom_1(7866) <= 2363;
srom_1(7867) <= 8399;
srom_1(7868) <= 53732;
srom_1(7869) <= 138150;
srom_1(7870) <= 261257;
srom_1(7871) <= 422477;
srom_1(7872) <= 621052;
srom_1(7873) <= 856052;
srom_1(7874) <= 1126375;
srom_1(7875) <= 1430753;
srom_1(7876) <= 1767759;
srom_1(7877) <= 2135812;
srom_1(7878) <= 2533186;
srom_1(7879) <= 2958019;
srom_1(7880) <= 3408317;
srom_1(7881) <= 3881970;
srom_1(7882) <= 4376756;
srom_1(7883) <= 4890355;
srom_1(7884) <= 5420359;
srom_1(7885) <= 5964281;
srom_1(7886) <= 6519572;
srom_1(7887) <= 7083628;
srom_1(7888) <= 7653803;
srom_1(7889) <= 8227424;
srom_1(7890) <= 8801801;
srom_1(7891) <= 9374240;
srom_1(7892) <= 9942057;
srom_1(7893) <= 10502589;
srom_1(7894) <= 11053209;
srom_1(7895) <= 11591333;
srom_1(7896) <= 12114438;
srom_1(7897) <= 12620072;
srom_1(7898) <= 13105862;
srom_1(7899) <= 13569532;
srom_1(7900) <= 14008907;
srom_1(7901) <= 14421927;
srom_1(7902) <= 14806654;
srom_1(7903) <= 15161284;
srom_1(7904) <= 15484156;
srom_1(7905) <= 15773753;
srom_1(7906) <= 16028720;
srom_1(7907) <= 16247859;
srom_1(7908) <= 16430143;
srom_1(7909) <= 16574718;
srom_1(7910) <= 16680905;
srom_1(7911) <= 16748207;
srom_1(7912) <= 16776308;
srom_1(7913) <= 16765076;
srom_1(7914) <= 16714564;
srom_1(7915) <= 16625009;
srom_1(7916) <= 16496830;
srom_1(7917) <= 16330629;
srom_1(7918) <= 16127186;
srom_1(7919) <= 15887453;
srom_1(7920) <= 15612556;
srom_1(7921) <= 15303783;
srom_1(7922) <= 14962582;
srom_1(7923) <= 14590554;
srom_1(7924) <= 14189443;
srom_1(7925) <= 13761130;
srom_1(7926) <= 13307623;
srom_1(7927) <= 12831049;
srom_1(7928) <= 12333643;
srom_1(7929) <= 11817737;
srom_1(7930) <= 11285751;
srom_1(7931) <= 10740179;
srom_1(7932) <= 10183580;
srom_1(7933) <= 9618564;
srom_1(7934) <= 9047780;
srom_1(7935) <= 8473905;
srom_1(7936) <= 7899630;
srom_1(7937) <= 7327648;
srom_1(7938) <= 6760641;
srom_1(7939) <= 6201268;
srom_1(7940) <= 5652152;
srom_1(7941) <= 5115869;
srom_1(7942) <= 4594932;
srom_1(7943) <= 4091786;
srom_1(7944) <= 3608788;
srom_1(7945) <= 3148205;
srom_1(7946) <= 2712196;
srom_1(7947) <= 2302806;
srom_1(7948) <= 1921954;
srom_1(7949) <= 1571426;
srom_1(7950) <= 1252866;
srom_1(7951) <= 967769;
srom_1(7952) <= 717470;
srom_1(7953) <= 503144;
srom_1(7954) <= 325795;
srom_1(7955) <= 186256;
srom_1(7956) <= 85180;
srom_1(7957) <= 23042;
srom_1(7958) <= 133;
srom_1(7959) <= 16561;
srom_1(7960) <= 72247;
srom_1(7961) <= 166933;
srom_1(7962) <= 300172;
srom_1(7963) <= 471341;
srom_1(7964) <= 679636;
srom_1(7965) <= 924082;
srom_1(7966) <= 1203531;
srom_1(7967) <= 1516674;
srom_1(7968) <= 1862041;
srom_1(7969) <= 2238014;
srom_1(7970) <= 2642829;
srom_1(7971) <= 3074588;
srom_1(7972) <= 3531266;
srom_1(7973) <= 4010722;
srom_1(7974) <= 4510707;
srom_1(7975) <= 5028877;
srom_1(7976) <= 5562802;
srom_1(7977) <= 6109979;
srom_1(7978) <= 6667840;
srom_1(7979) <= 7233771;
srom_1(7980) <= 7805117;
srom_1(7981) <= 8379199;
srom_1(7982) <= 8953326;
srom_1(7983) <= 9524804;
srom_1(7984) <= 10090954;
srom_1(7985) <= 10649122;
srom_1(7986) <= 11196689;
srom_1(7987) <= 11731088;
srom_1(7988) <= 12249813;
srom_1(7989) <= 12750431;
srom_1(7990) <= 13230596;
srom_1(7991) <= 13688054;
srom_1(7992) <= 14120662;
srom_1(7993) <= 14526390;
srom_1(7994) <= 14903336;
srom_1(7995) <= 15249732;
srom_1(7996) <= 15563954;
srom_1(7997) <= 15844528;
srom_1(7998) <= 16090139;
srom_1(7999) <= 16299635;
srom_1(8000) <= 16472033;
srom_1(8001) <= 16606525;
srom_1(8002) <= 16702481;
srom_1(8003) <= 16759450;
srom_1(8004) <= 16777165;
srom_1(8005) <= 16755543;
srom_1(8006) <= 16694686;
srom_1(8007) <= 16594879;
srom_1(8008) <= 16456590;
srom_1(8009) <= 16280467;
srom_1(8010) <= 16067337;
srom_1(8011) <= 15818199;
srom_1(8012) <= 15534220;
srom_1(8013) <= 15216733;
srom_1(8014) <= 14867227;
srom_1(8015) <= 14487341;
srom_1(8016) <= 14078855;
srom_1(8017) <= 13643686;
srom_1(8018) <= 13183874;
srom_1(8019) <= 12701575;
srom_1(8020) <= 12199051;
srom_1(8021) <= 11678659;
srom_1(8022) <= 11142839;
srom_1(8023) <= 10594103;
srom_1(8024) <= 10035025;
srom_1(8025) <= 9468226;
srom_1(8026) <= 8896364;
srom_1(8027) <= 8322122;
srom_1(8028) <= 7748191;
srom_1(8029) <= 7177263;
srom_1(8030) <= 6612016;
srom_1(8031) <= 6055099;
srom_1(8032) <= 5509126;
srom_1(8033) <= 4976655;
srom_1(8034) <= 4460184;
srom_1(8035) <= 3962135;
srom_1(8036) <= 3484843;
srom_1(8037) <= 3030546;
srom_1(8038) <= 2601375;
srom_1(8039) <= 2199343;
srom_1(8040) <= 1826334;
srom_1(8041) <= 1484098;
srom_1(8042) <= 1174239;
srom_1(8043) <= 898212;
srom_1(8044) <= 657309;
srom_1(8045) <= 452661;
srom_1(8046) <= 285227;
srom_1(8047) <= 155793;
srom_1(8048) <= 64965;
srom_1(8049) <= 13170;
srom_1(8050) <= 650;
srom_1(8051) <= 27464;
srom_1(8052) <= 93486;
srom_1(8053) <= 198407;
srom_1(8054) <= 341734;
srom_1(8055) <= 522797;
srom_1(8056) <= 740744;
srom_1(8057) <= 994555;
srom_1(8058) <= 1283040;
srom_1(8059) <= 1604844;
srom_1(8060) <= 1958461;
srom_1(8061) <= 2342230;
srom_1(8062) <= 2754353;
srom_1(8063) <= 3192897;
srom_1(8064) <= 3655805;
srom_1(8065) <= 4140907;
srom_1(8066) <= 4645928;
srom_1(8067) <= 5168500;
srom_1(8068) <= 5706171;
srom_1(8069) <= 6256422;
srom_1(8070) <= 6816671;
srom_1(8071) <= 7384292;
srom_1(8072) <= 7956622;
srom_1(8073) <= 8530978;
srom_1(8074) <= 9104666;
srom_1(8075) <= 9674997;
srom_1(8076) <= 10239295;
srom_1(8077) <= 10794914;
srom_1(8078) <= 11339250;
srom_1(8079) <= 11869749;
srom_1(8080) <= 12383924;
srom_1(8081) <= 12879363;
srom_1(8082) <= 13353744;
srom_1(8083) <= 13804841;
srom_1(8084) <= 14230540;
srom_1(8085) <= 14628844;
srom_1(8086) <= 14997885;
srom_1(8087) <= 15335933;
srom_1(8088) <= 15641403;
srom_1(8089) <= 15912862;
srom_1(8090) <= 16149037;
srom_1(8091) <= 16348821;
srom_1(8092) <= 16511276;
srom_1(8093) <= 16635642;
srom_1(8094) <= 16721334;
srom_1(8095) <= 16767952;
srom_1(8096) <= 16775275;
srom_1(8097) <= 16743271;
srom_1(8098) <= 16672089;
srom_1(8099) <= 16562063;
srom_1(8100) <= 16413709;
srom_1(8101) <= 16227722;
srom_1(8102) <= 16004975;
srom_1(8103) <= 15746512;
srom_1(8104) <= 15453545;
srom_1(8105) <= 15127449;
srom_1(8106) <= 14769751;
srom_1(8107) <= 14382131;
srom_1(8108) <= 13966404;
srom_1(8109) <= 13524522;
srom_1(8110) <= 13058555;
srom_1(8111) <= 12570689;
srom_1(8112) <= 12063212;
srom_1(8113) <= 11538504;
srom_1(8114) <= 10999025;
srom_1(8115) <= 10447304;
srom_1(8116) <= 9885930;
srom_1(8117) <= 9317534;
srom_1(8118) <= 8744782;
srom_1(8119) <= 8170360;
srom_1(8120) <= 7596961;
srom_1(8121) <= 7027275;
srom_1(8122) <= 6463972;
srom_1(8123) <= 5909695;
srom_1(8124) <= 5367042;
srom_1(8125) <= 4838558;
srom_1(8126) <= 4326722;
srom_1(8127) <= 3833933;
srom_1(8128) <= 3362503;
srom_1(8129) <= 2914641;
srom_1(8130) <= 2492449;
srom_1(8131) <= 2097907;
srom_1(8132) <= 1732863;
srom_1(8133) <= 1399030;
srom_1(8134) <= 1097974;
srom_1(8135) <= 831107;
srom_1(8136) <= 599679;
srom_1(8137) <= 404776;
srom_1(8138) <= 247312;
srom_1(8139) <= 128025;
srom_1(8140) <= 47475;
srom_1(8141) <= 6039;
srom_1(8142) <= 3912;
srom_1(8143) <= 41104;
srom_1(8144) <= 117440;
srom_1(8145) <= 232562;
srom_1(8146) <= 385931;
srom_1(8147) <= 576828;
srom_1(8148) <= 804356;
srom_1(8149) <= 1067449;
srom_1(8150) <= 1364874;
srom_1(8151) <= 1695236;
srom_1(8152) <= 2056985;
srom_1(8153) <= 2448425;
srom_1(8154) <= 2867721;
srom_1(8155) <= 3312906;
srom_1(8156) <= 3781893;
srom_1(8157) <= 4272483;
srom_1(8158) <= 4782374;
srom_1(8159) <= 5309176;
srom_1(8160) <= 5850419;
srom_1(8161) <= 6403564;
srom_1(8162) <= 6966017;
srom_1(8163) <= 7535142;
srom_1(8164) <= 8108269;
srom_1(8165) <= 8682710;
srom_1(8166) <= 9255772;
srom_1(8167) <= 9824768;
srom_1(8168) <= 10387029;
srom_1(8169) <= 10939919;
srom_1(8170) <= 11480845;
srom_1(8171) <= 12007270;
srom_1(8172) <= 12516726;
srom_1(8173) <= 13006824;
srom_1(8174) <= 13475266;
srom_1(8175) <= 13919854;
srom_1(8176) <= 14338505;
srom_1(8177) <= 14729254;
srom_1(8178) <= 15090270;
srom_1(8179) <= 15419860;
srom_1(8180) <= 15716478;
srom_1(8181) <= 15978732;
srom_1(8182) <= 16205394;
srom_1(8183) <= 16395401;
srom_1(8184) <= 16547860;
srom_1(8185) <= 16662059;
srom_1(8186) <= 16737460;
srom_1(8187) <= 16773710;
srom_1(8188) <= 16770640;
srom_1(8189) <= 16728264;
srom_1(8190) <= 16646780;
srom_1(8191) <= 16526571;
srom_1(8192) <= 16368200;
srom_1(8193) <= 16172410;
srom_1(8194) <= 15940119;
srom_1(8195) <= 15672416;
srom_1(8196) <= 15370557;
srom_1(8197) <= 15035958;
srom_1(8198) <= 14670186;
srom_1(8199) <= 14274958;
srom_1(8200) <= 13852127;
srom_1(8201) <= 13403676;
srom_1(8202) <= 12931707;
srom_1(8203) <= 12438434;
srom_1(8204) <= 11926171;
srom_1(8205) <= 11397318;
srom_1(8206) <= 10854356;
srom_1(8207) <= 10299832;
srom_1(8208) <= 9736345;
srom_1(8209) <= 9166538;
srom_1(8210) <= 8593084;
srom_1(8211) <= 8018670;
srom_1(8212) <= 7445991;
srom_1(8213) <= 6877733;
srom_1(8214) <= 6316559;
srom_1(8215) <= 5765102;
srom_1(8216) <= 5225947;
srom_1(8217) <= 4701624;
srom_1(8218) <= 4194589;
srom_1(8219) <= 3707222;
srom_1(8220) <= 3241808;
srom_1(8221) <= 2800529;
srom_1(8222) <= 2385454;
srom_1(8223) <= 1998530;
srom_1(8224) <= 1641571;
srom_1(8225) <= 1316251;
srom_1(8226) <= 1024096;
srom_1(8227) <= 766476;
srom_1(8228) <= 544599;
srom_1(8229) <= 359505;
srom_1(8230) <= 212062;
srom_1(8231) <= 102961;
srom_1(8232) <= 32715;
srom_1(8233) <= 1653;
srom_1(8234) <= 9920;
srom_1(8235) <= 57477;
srom_1(8236) <= 144102;
srom_1(8237) <= 269388;
srom_1(8238) <= 432748;
srom_1(8239) <= 633416;
srom_1(8240) <= 870451;
srom_1(8241) <= 1142741;
srom_1(8242) <= 1449009;
srom_1(8243) <= 1787819;
srom_1(8244) <= 2157583;
srom_1(8245) <= 2556566;
srom_1(8246) <= 2982897;
srom_1(8247) <= 3434578;
srom_1(8248) <= 3909490;
srom_1(8249) <= 4405406;
srom_1(8250) <= 4920000;
srom_1(8251) <= 5450861;
srom_1(8252) <= 5995497;
srom_1(8253) <= 6551355;
srom_1(8254) <= 7115829;
srom_1(8255) <= 7686271;
srom_1(8256) <= 8260007;
srom_1(8257) <= 8834346;
srom_1(8258) <= 9406594;
srom_1(8259) <= 9974069;
srom_1(8260) <= 10534109;
srom_1(8261) <= 11084088;
srom_1(8262) <= 11621428;
srom_1(8263) <= 12143607;
srom_1(8264) <= 12648178;
srom_1(8265) <= 13132774;
srom_1(8266) <= 13595123;
srom_1(8267) <= 14033057;
srom_1(8268) <= 14444522;
srom_1(8269) <= 14827589;
srom_1(8270) <= 15180462;
srom_1(8271) <= 15501485;
srom_1(8272) <= 15789153;
srom_1(8273) <= 16042118;
srom_1(8274) <= 16259192;
srom_1(8275) <= 16439359;
srom_1(8276) <= 16581773;
srom_1(8277) <= 16685767;
srom_1(8278) <= 16750852;
srom_1(8279) <= 16776724;
srom_1(8280) <= 16763261;
srom_1(8281) <= 16710526;
srom_1(8282) <= 16618767;
srom_1(8283) <= 16488414;
srom_1(8284) <= 16320078;
srom_1(8285) <= 16114549;
srom_1(8286) <= 15872790;
srom_1(8287) <= 15595936;
srom_1(8288) <= 15285283;
srom_1(8289) <= 14942290;
srom_1(8290) <= 14568564;
srom_1(8291) <= 14165859;
srom_1(8292) <= 13736062;
srom_1(8293) <= 13281189;
srom_1(8294) <= 12803372;
srom_1(8295) <= 12304854;
srom_1(8296) <= 11787971;
srom_1(8297) <= 11255147;
srom_1(8298) <= 10708880;
srom_1(8299) <= 10151734;
srom_1(8300) <= 9586319;
srom_1(8301) <= 9015288;
srom_1(8302) <= 8441318;
srom_1(8303) <= 7867101;
srom_1(8304) <= 7295330;
srom_1(8305) <= 6728685;
srom_1(8306) <= 6169824;
srom_1(8307) <= 5621368;
srom_1(8308) <= 5085888;
srom_1(8309) <= 4565896;
srom_1(8310) <= 4063830;
srom_1(8311) <= 3582044;
srom_1(8312) <= 3122798;
srom_1(8313) <= 2688245;
srom_1(8314) <= 2280423;
srom_1(8315) <= 1901245;
srom_1(8316) <= 1552488;
srom_1(8317) <= 1235788;
srom_1(8318) <= 952629;
srom_1(8319) <= 704341;
srom_1(8320) <= 492087;
srom_1(8321) <= 316862;
srom_1(8322) <= 179489;
srom_1(8323) <= 80611;
srom_1(8324) <= 20692;
srom_1(8325) <= 12;
srom_1(8326) <= 18670;
srom_1(8327) <= 76578;
srom_1(8328) <= 173463;
srom_1(8329) <= 308872;
srom_1(8330) <= 482170;
srom_1(8331) <= 692544;
srom_1(8332) <= 939007;
srom_1(8333) <= 1220404;
srom_1(8334) <= 1535415;
srom_1(8335) <= 1882563;
srom_1(8336) <= 2260220;
srom_1(8337) <= 2666615;
srom_1(8338) <= 3099843;
srom_1(8339) <= 3557871;
srom_1(8340) <= 4038553;
srom_1(8341) <= 4539633;
srom_1(8342) <= 5058763;
srom_1(8343) <= 5593507;
srom_1(8344) <= 6141358;
srom_1(8345) <= 6699748;
srom_1(8346) <= 7266057;
srom_1(8347) <= 7837630;
srom_1(8348) <= 8411787;
srom_1(8349) <= 8985835;
srom_1(8350) <= 9557083;
srom_1(8351) <= 10122851;
srom_1(8352) <= 10680487;
srom_1(8353) <= 11227375;
srom_1(8354) <= 11760952;
srom_1(8355) <= 12278714;
srom_1(8356) <= 12778234;
srom_1(8357) <= 13257170;
srom_1(8358) <= 13713276;
srom_1(8359) <= 14144412;
srom_1(8360) <= 14548557;
srom_1(8361) <= 14923816;
srom_1(8362) <= 15268429;
srom_1(8363) <= 15580781;
srom_1(8364) <= 15859406;
srom_1(8365) <= 16102997;
srom_1(8366) <= 16310414;
srom_1(8367) <= 16480682;
srom_1(8368) <= 16613004;
srom_1(8369) <= 16706758;
srom_1(8370) <= 16761506;
srom_1(8371) <= 16776991;
srom_1(8372) <= 16753139;
srom_1(8373) <= 16690064;
srom_1(8374) <= 16588060;
srom_1(8375) <= 16447606;
srom_1(8376) <= 16269360;
srom_1(8377) <= 16054159;
srom_1(8378) <= 15803012;
srom_1(8379) <= 15517096;
srom_1(8380) <= 15197752;
srom_1(8381) <= 14846477;
srom_1(8382) <= 14464920;
srom_1(8383) <= 14054868;
srom_1(8384) <= 13618245;
srom_1(8385) <= 13157099;
srom_1(8386) <= 12673592;
srom_1(8387) <= 12169991;
srom_1(8388) <= 11648658;
srom_1(8389) <= 11112037;
srom_1(8390) <= 10562645;
srom_1(8391) <= 10003058;
srom_1(8392) <= 9435901;
srom_1(8393) <= 8863832;
srom_1(8394) <= 8289535;
srom_1(8395) <= 7715703;
srom_1(8396) <= 7145026;
srom_1(8397) <= 6580181;
srom_1(8398) <= 6023815;
srom_1(8399) <= 5478540;
srom_1(8400) <= 4946910;
srom_1(8401) <= 4431420;
srom_1(8402) <= 3934487;
srom_1(8403) <= 3458440;
srom_1(8404) <= 3005513;
srom_1(8405) <= 2577828;
srom_1(8406) <= 2177393;
srom_1(8407) <= 1806084;
srom_1(8408) <= 1465643;
srom_1(8409) <= 1157666;
srom_1(8410) <= 883597;
srom_1(8411) <= 644722;
srom_1(8412) <= 442160;
srom_1(8413) <= 276862;
srom_1(8414) <= 149603;
srom_1(8415) <= 60980;
srom_1(8416) <= 11407;
srom_1(8417) <= 1119;
srom_1(8418) <= 30161;
srom_1(8419) <= 98400;
srom_1(8420) <= 205514;
srom_1(8421) <= 351002;
srom_1(8422) <= 534180;
srom_1(8423) <= 754191;
srom_1(8424) <= 1010002;
srom_1(8425) <= 1300414;
srom_1(8426) <= 1624065;
srom_1(8427) <= 1979437;
srom_1(8428) <= 2364864;
srom_1(8429) <= 2778538;
srom_1(8430) <= 3218520;
srom_1(8431) <= 3682746;
srom_1(8432) <= 4169040;
srom_1(8433) <= 4675121;
srom_1(8434) <= 5198615;
srom_1(8435) <= 5737068;
srom_1(8436) <= 6287956;
srom_1(8437) <= 6848694;
srom_1(8438) <= 7416653;
srom_1(8439) <= 7989170;
srom_1(8440) <= 8563560;
srom_1(8441) <= 9137130;
srom_1(8442) <= 9707189;
srom_1(8443) <= 10271066;
srom_1(8444) <= 10826114;
srom_1(8445) <= 11369733;
srom_1(8446) <= 11899372;
srom_1(8447) <= 12412548;
srom_1(8448) <= 12906854;
srom_1(8449) <= 13379972;
srom_1(8450) <= 13829685;
srom_1(8451) <= 14253882;
srom_1(8452) <= 14650575;
srom_1(8453) <= 15017903;
srom_1(8454) <= 15354145;
srom_1(8455) <= 15657722;
srom_1(8456) <= 15927212;
srom_1(8457) <= 16161351;
srom_1(8458) <= 16359041;
srom_1(8459) <= 16519355;
srom_1(8460) <= 16641541;
srom_1(8461) <= 16725027;
srom_1(8462) <= 16769419;
srom_1(8463) <= 16774512;
srom_1(8464) <= 16740280;
srom_1(8465) <= 16666884;
srom_1(8466) <= 16554668;
srom_1(8467) <= 16404159;
srom_1(8468) <= 16216062;
srom_1(8469) <= 15991260;
srom_1(8470) <= 15730806;
srom_1(8471) <= 15435922;
srom_1(8472) <= 15107991;
srom_1(8473) <= 14748550;
srom_1(8474) <= 14359285;
srom_1(8475) <= 13942022;
srom_1(8476) <= 13498717;
srom_1(8477) <= 13031449;
srom_1(8478) <= 12542409;
srom_1(8479) <= 12033890;
srom_1(8480) <= 11508277;
srom_1(8481) <= 10968035;
srom_1(8482) <= 10415698;
srom_1(8483) <= 9853854;
srom_1(8484) <= 9285140;
srom_1(8485) <= 8712221;
srom_1(8486) <= 8137785;
srom_1(8487) <= 7564525;
srom_1(8488) <= 6995129;
srom_1(8489) <= 6432268;
srom_1(8490) <= 5878581;
srom_1(8491) <= 5336664;
srom_1(8492) <= 4809059;
srom_1(8493) <= 4298240;
srom_1(8494) <= 3806601;
srom_1(8495) <= 3336450;
srom_1(8496) <= 2889989;
srom_1(8497) <= 2469314;
srom_1(8498) <= 2076396;
srom_1(8499) <= 1713078;
srom_1(8500) <= 1381064;
srom_1(8501) <= 1081911;
srom_1(8502) <= 817021;
srom_1(8503) <= 587638;
srom_1(8504) <= 394835;
srom_1(8505) <= 239518;
srom_1(8506) <= 122415;
srom_1(8507) <= 44075;
srom_1(8508) <= 4866;
srom_1(8509) <= 4971;
srom_1(8510) <= 44389;
srom_1(8511) <= 122936;
srom_1(8512) <= 240244;
srom_1(8513) <= 395762;
srom_1(8514) <= 588762;
srom_1(8515) <= 818338;
srom_1(8516) <= 1083413;
srom_1(8517) <= 1382745;
srom_1(8518) <= 1714930;
srom_1(8519) <= 2078409;
srom_1(8520) <= 2471480;
srom_1(8521) <= 2892298;
srom_1(8522) <= 3338890;
srom_1(8523) <= 3809162;
srom_1(8524) <= 4300909;
srom_1(8525) <= 4811824;
srom_1(8526) <= 5339512;
srom_1(8527) <= 5881498;
srom_1(8528) <= 6435241;
srom_1(8529) <= 6998144;
srom_1(8530) <= 7567567;
srom_1(8531) <= 8140840;
srom_1(8532) <= 8715276;
srom_1(8533) <= 9288179;
srom_1(8534) <= 9856864;
srom_1(8535) <= 10418664;
srom_1(8536) <= 10970944;
srom_1(8537) <= 11511114;
srom_1(8538) <= 12036643;
srom_1(8539) <= 12545064;
srom_1(8540) <= 13033994;
srom_1(8541) <= 13501141;
srom_1(8542) <= 13944313;
srom_1(8543) <= 14361432;
srom_1(8544) <= 14750543;
srom_1(8545) <= 15109820;
srom_1(8546) <= 15437579;
srom_1(8547) <= 15732284;
srom_1(8548) <= 15992551;
srom_1(8549) <= 16217161;
srom_1(8550) <= 16405060;
srom_1(8551) <= 16555367;
srom_1(8552) <= 16667377;
srom_1(8553) <= 16740566;
srom_1(8554) <= 16774589;
srom_1(8555) <= 16769287;
srom_1(8556) <= 16724686;
srom_1(8557) <= 16640993;
srom_1(8558) <= 16518603;
srom_1(8559) <= 16358088;
srom_1(8560) <= 16160201;
srom_1(8561) <= 15925871;
srom_1(8562) <= 15656196;
srom_1(8563) <= 15352441;
srom_1(8564) <= 15016030;
srom_1(8565) <= 14648541;
srom_1(8566) <= 14251696;
srom_1(8567) <= 13827358;
srom_1(8568) <= 13377515;
srom_1(8569) <= 12904278;
srom_1(8570) <= 12409865;
srom_1(8571) <= 11896596;
srom_1(8572) <= 11366876;
srom_1(8573) <= 10823190;
srom_1(8574) <= 10268087;
srom_1(8575) <= 9704171;
srom_1(8576) <= 9134085;
srom_1(8577) <= 8560504;
srom_1(8578) <= 7986117;
srom_1(8579) <= 7413617;
srom_1(8580) <= 6845689;
srom_1(8581) <= 6284997;
srom_1(8582) <= 5734169;
srom_1(8583) <= 5195788;
srom_1(8584) <= 4672380;
srom_1(8585) <= 4166399;
srom_1(8586) <= 3680216;
srom_1(8587) <= 3216114;
srom_1(8588) <= 2776266;
srom_1(8589) <= 2362737;
srom_1(8590) <= 1977465;
srom_1(8591) <= 1622258;
srom_1(8592) <= 1298780;
srom_1(8593) <= 1008549;
srom_1(8594) <= 752925;
srom_1(8595) <= 533108;
srom_1(8596) <= 350127;
srom_1(8597) <= 204842;
srom_1(8598) <= 97934;
srom_1(8599) <= 29903;
srom_1(8600) <= 1069;
srom_1(8601) <= 11567;
srom_1(8602) <= 61348;
srom_1(8603) <= 150179;
srom_1(8604) <= 277642;
srom_1(8605) <= 443140;
srom_1(8606) <= 645897;
srom_1(8607) <= 884963;
srom_1(8608) <= 1159216;
srom_1(8609) <= 1467369;
srom_1(8610) <= 1807979;
srom_1(8611) <= 2179448;
srom_1(8612) <= 2580033;
srom_1(8613) <= 3007857;
srom_1(8614) <= 3460913;
srom_1(8615) <= 3937077;
srom_1(8616) <= 4434116;
srom_1(8617) <= 4949698;
srom_1(8618) <= 5481407;
srom_1(8619) <= 6026748;
srom_1(8620) <= 6583165;
srom_1(8621) <= 7148049;
srom_1(8622) <= 7718750;
srom_1(8623) <= 8292592;
srom_1(8624) <= 8866884;
srom_1(8625) <= 9438934;
srom_1(8626) <= 10006058;
srom_1(8627) <= 10565597;
srom_1(8628) <= 11114928;
srom_1(8629) <= 11651474;
srom_1(8630) <= 12172719;
srom_1(8631) <= 12676219;
srom_1(8632) <= 13159614;
srom_1(8633) <= 13620635;
srom_1(8634) <= 14057122;
srom_1(8635) <= 14467027;
srom_1(8636) <= 14848428;
srom_1(8637) <= 15199536;
srom_1(8638) <= 15518707;
srom_1(8639) <= 15804441;
srom_1(8640) <= 16055400;
srom_1(8641) <= 16270407;
srom_1(8642) <= 16448454;
srom_1(8643) <= 16588705;
srom_1(8644) <= 16690503;
srom_1(8645) <= 16753370;
srom_1(8646) <= 16777013;
srom_1(8647) <= 16761319;
srom_1(8648) <= 16706362;
srom_1(8649) <= 16612401;
srom_1(8650) <= 16479876;
srom_1(8651) <= 16309408;
srom_1(8652) <= 16101796;
srom_1(8653) <= 15858015;
srom_1(8654) <= 15579207;
srom_1(8655) <= 15266680;
srom_1(8656) <= 14921899;
srom_1(8657) <= 14546482;
srom_1(8658) <= 14142188;
srom_1(8659) <= 13710913;
srom_1(8660) <= 13254681;
srom_1(8661) <= 12775629;
srom_1(8662) <= 12276006;
srom_1(8663) <= 11758153;
srom_1(8664) <= 11224499;
srom_1(8665) <= 10677547;
srom_1(8666) <= 10119861;
srom_1(8667) <= 9554056;
srom_1(8668) <= 8982787;
srom_1(8669) <= 8408731;
srom_1(8670) <= 7834580;
srom_1(8671) <= 7263028;
srom_1(8672) <= 6696754;
srom_1(8673) <= 6138414;
srom_1(8674) <= 5590625;
srom_1(8675) <= 5055957;
srom_1(8676) <= 4536918;
srom_1(8677) <= 4035940;
srom_1(8678) <= 3555373;
srom_1(8679) <= 3097471;
srom_1(8680) <= 2664381;
srom_1(8681) <= 2258133;
srom_1(8682) <= 1880634;
srom_1(8683) <= 1533653;
srom_1(8684) <= 1218817;
srom_1(8685) <= 937602;
srom_1(8686) <= 691328;
srom_1(8687) <= 481149;
srom_1(8688) <= 308051;
srom_1(8689) <= 172846;
srom_1(8690) <= 76166;
srom_1(8691) <= 18467;
srom_1(8692) <= 18;
srom_1(8693) <= 20907;
srom_1(8694) <= 81034;
srom_1(8695) <= 180118;
srom_1(8696) <= 317695;
srom_1(8697) <= 493119;
srom_1(8698) <= 705568;
srom_1(8699) <= 954045;
srom_1(8700) <= 1237385;
srom_1(8701) <= 1554260;
srom_1(8702) <= 1903183;
srom_1(8703) <= 2282519;
srom_1(8704) <= 2690488;
srom_1(8705) <= 3125178;
srom_1(8706) <= 3584550;
srom_1(8707) <= 4066449;
srom_1(8708) <= 4568617;
srom_1(8709) <= 5088698;
srom_1(8710) <= 5624254;
srom_1(8711) <= 6172772;
srom_1(8712) <= 6731681;
srom_1(8713) <= 7298360;
srom_1(8714) <= 7870152;
srom_1(8715) <= 8444375;
srom_1(8716) <= 9018336;
srom_1(8717) <= 9589344;
srom_1(8718) <= 10154722;
srom_1(8719) <= 10711818;
srom_1(8720) <= 11258019;
srom_1(8721) <= 11790765;
srom_1(8722) <= 12307557;
srom_1(8723) <= 12805971;
srom_1(8724) <= 13283671;
srom_1(8725) <= 13738416;
srom_1(8726) <= 14168075;
srom_1(8727) <= 14570631;
srom_1(8728) <= 14944198;
srom_1(8729) <= 15287023;
srom_1(8730) <= 15597499;
srom_1(8731) <= 15874171;
srom_1(8732) <= 16115739;
srom_1(8733) <= 16321073;
srom_1(8734) <= 16489209;
srom_1(8735) <= 16619358;
srom_1(8736) <= 16710910;
srom_1(8737) <= 16763436;
srom_1(8738) <= 16776690;
srom_1(8739) <= 16750609;
srom_1(8740) <= 16685316;
srom_1(8741) <= 16581117;
srom_1(8742) <= 16438500;
srom_1(8743) <= 16258134;
srom_1(8744) <= 16040866;
srom_1(8745) <= 15787713;
srom_1(8746) <= 15499864;
srom_1(8747) <= 15178667;
srom_1(8748) <= 14825630;
srom_1(8749) <= 14442407;
srom_1(8750) <= 14030795;
srom_1(8751) <= 13592726;
srom_1(8752) <= 13130253;
srom_1(8753) <= 12645544;
srom_1(8754) <= 12140873;
srom_1(8755) <= 11618607;
srom_1(8756) <= 11081194;
srom_1(8757) <= 10531154;
srom_1(8758) <= 9971068;
srom_1(8759) <= 9403560;
srom_1(8760) <= 8831293;
srom_1(8761) <= 8256951;
srom_1(8762) <= 7683225;
srom_1(8763) <= 7112808;
srom_1(8764) <= 6548373;
srom_1(8765) <= 5992567;
srom_1(8766) <= 5447998;
srom_1(8767) <= 4917218;
srom_1(8768) <= 4402716;
srom_1(8769) <= 3906906;
srom_1(8770) <= 3432112;
srom_1(8771) <= 2980560;
srom_1(8772) <= 2554369;
srom_1(8773) <= 2155537;
srom_1(8774) <= 1785933;
srom_1(8775) <= 1447292;
srom_1(8776) <= 1141201;
srom_1(8777) <= 869095;
srom_1(8778) <= 632252;
srom_1(8779) <= 431780;
srom_1(8780) <= 268620;
srom_1(8781) <= 143538;
srom_1(8782) <= 57120;
srom_1(8783) <= 9772;
srom_1(8784) <= 1714;
srom_1(8785) <= 32986;
srom_1(8786) <= 103439;
srom_1(8787) <= 212745;
srom_1(8788) <= 360390;
srom_1(8789) <= 545683;
srom_1(8790) <= 767753;
srom_1(8791) <= 1025560;
srom_1(8792) <= 1317895;
srom_1(8793) <= 1643388;
srom_1(8794) <= 2000510;
srom_1(8795) <= 2387589;
srom_1(8796) <= 2802809;
srom_1(8797) <= 3244222;
srom_1(8798) <= 3709759;
srom_1(8799) <= 4197237;
srom_1(8800) <= 4704369;
srom_1(8801) <= 5228779;
srom_1(8802) <= 5768005;
srom_1(8803) <= 6319521;
srom_1(8804) <= 6880739;
srom_1(8805) <= 7449029;
srom_1(8806) <= 8021724;
srom_1(8807) <= 8596139;
srom_1(8808) <= 9169582;
srom_1(8809) <= 9739362;
srom_1(8810) <= 10302808;
srom_1(8811) <= 10857278;
srom_1(8812) <= 11400171;
srom_1(8813) <= 11928942;
srom_1(8814) <= 12441111;
srom_1(8815) <= 12934277;
srom_1(8816) <= 13406126;
srom_1(8817) <= 13854446;
srom_1(8818) <= 14277136;
srom_1(8819) <= 14672212;
srom_1(8820) <= 15037822;
srom_1(8821) <= 15372251;
srom_1(8822) <= 15673932;
srom_1(8823) <= 15941449;
srom_1(8824) <= 16173549;
srom_1(8825) <= 16369142;
srom_1(8826) <= 16527312;
srom_1(8827) <= 16647316;
srom_1(8828) <= 16728593;
srom_1(8829) <= 16770761;
srom_1(8830) <= 16773621;
srom_1(8831) <= 16737162;
srom_1(8832) <= 16661553;
srom_1(8833) <= 16547150;
srom_1(8834) <= 16394488;
srom_1(8835) <= 16204284;
srom_1(8836) <= 15977430;
srom_1(8837) <= 15714989;
srom_1(8838) <= 15418192;
srom_1(8839) <= 15088431;
srom_1(8840) <= 14727253;
srom_1(8841) <= 14336350;
srom_1(8842) <= 13917556;
srom_1(8843) <= 13472835;
srom_1(8844) <= 13004272;
srom_1(8845) <= 12514065;
srom_1(8846) <= 12004512;
srom_1(8847) <= 11478003;
srom_1(8848) <= 10937007;
srom_1(8849) <= 10384060;
srom_1(8850) <= 9821756;
srom_1(8851) <= 9252732;
srom_1(8852) <= 8679655;
srom_1(8853) <= 8105214;
srom_1(8854) <= 7532101;
srom_1(8855) <= 6963005;
srom_1(8856) <= 6400594;
srom_1(8857) <= 5847505;
srom_1(8858) <= 5306333;
srom_1(8859) <= 4779614;
srom_1(8860) <= 4269820;
srom_1(8861) <= 3779339;
srom_1(8862) <= 3310473;
srom_1(8863) <= 2865420;
srom_1(8864) <= 2446268;
srom_1(8865) <= 2054981;
srom_1(8866) <= 1693394;
srom_1(8867) <= 1363204;
srom_1(8868) <= 1065958;
srom_1(8869) <= 803050;
srom_1(8870) <= 575714;
srom_1(8871) <= 385015;
srom_1(8872) <= 231848;
srom_1(8873) <= 116931;
srom_1(8874) <= 40802;
srom_1(8875) <= 3819;
srom_1(8876) <= 6156;
srom_1(8877) <= 47800;
srom_1(8878) <= 128557;
srom_1(8879) <= 248049;
srom_1(8880) <= 405714;
srom_1(8881) <= 600814;
srom_1(8882) <= 832434;
srom_1(8883) <= 1099487;
srom_1(8884) <= 1400721;
srom_1(8885) <= 1734724;
srom_1(8886) <= 2099929;
srom_1(8887) <= 2494624;
srom_1(8888) <= 2916958;
srom_1(8889) <= 3364950;
srom_1(8890) <= 3836500;
srom_1(8891) <= 4329396;
srom_1(8892) <= 4841328;
srom_1(8893) <= 5369894;
srom_1(8894) <= 5912615;
srom_1(8895) <= 6466947;
srom_1(8896) <= 7030291;
srom_1(8897) <= 7600004;
srom_1(8898) <= 8173416;
srom_1(8899) <= 8747836;
srom_1(8900) <= 9320572;
srom_1(8901) <= 9888937;
srom_1(8902) <= 10450267;
srom_1(8903) <= 11001930;
srom_1(8904) <= 11541337;
srom_1(8905) <= 12065960;
srom_1(8906) <= 12573339;
srom_1(8907) <= 13061094;
srom_1(8908) <= 13526938;
srom_1(8909) <= 13968687;
srom_1(8910) <= 14384269;
srom_1(8911) <= 14771735;
srom_1(8912) <= 15129268;
srom_1(8913) <= 15455193;
srom_1(8914) <= 15747979;
srom_1(8915) <= 16006255;
srom_1(8916) <= 16228809;
srom_1(8917) <= 16414598;
srom_1(8918) <= 16562750;
srom_1(8919) <= 16672571;
srom_1(8920) <= 16743545;
srom_1(8921) <= 16775341;
srom_1(8922) <= 16767807;
srom_1(8923) <= 16720981;
srom_1(8924) <= 16635082;
srom_1(8925) <= 16510512;
srom_1(8926) <= 16347856;
srom_1(8927) <= 16147876;
srom_1(8928) <= 15911510;
srom_1(8929) <= 15639867;
srom_1(8930) <= 15334220;
srom_1(8931) <= 14996002;
srom_1(8932) <= 14626801;
srom_1(8933) <= 14228346;
srom_1(8934) <= 13802506;
srom_1(8935) <= 13351280;
srom_1(8936) <= 12876781;
srom_1(8937) <= 12381236;
srom_1(8938) <= 11866968;
srom_1(8939) <= 11336388;
srom_1(8940) <= 10791986;
srom_1(8941) <= 10236313;
srom_1(8942) <= 9671976;
srom_1(8943) <= 9101621;
srom_1(8944) <= 8527922;
srom_1(8945) <= 7953570;
srom_1(8946) <= 7381257;
srom_1(8947) <= 6813669;
srom_1(8948) <= 6253466;
srom_1(8949) <= 5703275;
srom_1(8950) <= 5165677;
srom_1(8951) <= 4643193;
srom_1(8952) <= 4138271;
srom_1(8953) <= 3653282;
srom_1(8954) <= 3190497;
srom_1(8955) <= 2752089;
srom_1(8956) <= 2340112;
srom_1(8957) <= 1956498;
srom_1(8958) <= 1603047;
srom_1(8959) <= 1281415;
srom_1(8960) <= 993112;
srom_1(8961) <= 739489;
srom_1(8962) <= 521735;
srom_1(8963) <= 340871;
srom_1(8964) <= 197746;
srom_1(8965) <= 93031;
srom_1(8966) <= 27217;
srom_1(8967) <= 612;
srom_1(8968) <= 13341;
srom_1(8969) <= 65345;
srom_1(8970) <= 156379;
srom_1(8971) <= 286018;
srom_1(8972) <= 453652;
srom_1(8973) <= 658495;
srom_1(8974) <= 899588;
srom_1(8975) <= 1175800;
srom_1(8976) <= 1485834;
srom_1(8977) <= 1828239;
srom_1(8978) <= 2201407;
srom_1(8979) <= 2603589;
srom_1(8980) <= 3032898;
srom_1(8981) <= 3487323;
srom_1(8982) <= 3964731;
srom_1(8983) <= 4462885;
srom_1(8984) <= 4979448;
srom_1(8985) <= 5511997;
srom_1(8986) <= 6058036;
srom_1(8987) <= 6615003;
srom_1(8988) <= 7180288;
srom_1(8989) <= 7751238;
srom_1(8990) <= 8325178;
srom_1(8991) <= 8899415;
srom_1(8992) <= 9471257;
srom_1(8993) <= 10038022;
srom_1(8994) <= 10597052;
srom_1(8995) <= 11145726;
srom_1(8996) <= 11681471;
srom_1(8997) <= 12201774;
srom_1(8998) <= 12704196;
srom_1(8999) <= 13186381;
srom_1(9000) <= 13646068;
srom_1(9001) <= 14081101;
srom_1(9002) <= 14489439;
srom_1(9003) <= 14869169;
srom_1(9004) <= 15218509;
srom_1(9005) <= 15535821;
srom_1(9006) <= 15819617;
srom_1(9007) <= 16068567;
srom_1(9008) <= 16281503;
srom_1(9009) <= 16457427;
srom_1(9010) <= 16595512;
srom_1(9011) <= 16695113;
srom_1(9012) <= 16755762;
srom_1(9013) <= 16777175;
srom_1(9014) <= 16759250;
srom_1(9015) <= 16702073;
srom_1(9016) <= 16605911;
srom_1(9017) <= 16471215;
srom_1(9018) <= 16298618;
srom_1(9019) <= 16088927;
srom_1(9020) <= 15843127;
srom_1(9021) <= 15562370;
srom_1(9022) <= 15247973;
srom_1(9023) <= 14901410;
srom_1(9024) <= 14524306;
srom_1(9025) <= 14118430;
srom_1(9026) <= 13685684;
srom_1(9027) <= 13228099;
srom_1(9028) <= 12747820;
srom_1(9029) <= 12247099;
srom_1(9030) <= 11728284;
srom_1(9031) <= 11193808;
srom_1(9032) <= 10646178;
srom_1(9033) <= 10087961;
srom_1(9034) <= 9521776;
srom_1(9035) <= 8950276;
srom_1(9036) <= 8376143;
srom_1(9037) <= 7802068;
srom_1(9038) <= 7230743;
srom_1(9039) <= 6664849;
srom_1(9040) <= 6107037;
srom_1(9041) <= 5559925;
srom_1(9042) <= 5026077;
srom_1(9043) <= 4507997;
srom_1(9044) <= 4008115;
srom_1(9045) <= 3528774;
srom_1(9046) <= 3072223;
srom_1(9047) <= 2640602;
srom_1(9048) <= 2235936;
srom_1(9049) <= 1860121;
srom_1(9050) <= 1514921;
srom_1(9051) <= 1201954;
srom_1(9052) <= 922688;
srom_1(9053) <= 678432;
srom_1(9054) <= 470331;
srom_1(9055) <= 299362;
srom_1(9056) <= 166326;
srom_1(9057) <= 71848;
srom_1(9058) <= 16369;
srom_1(9059) <= 151;
srom_1(9060) <= 23269;
srom_1(9061) <= 85615;
srom_1(9062) <= 186897;
srom_1(9063) <= 326639;
srom_1(9064) <= 504187;
srom_1(9065) <= 718707;
srom_1(9066) <= 969194;
srom_1(9067) <= 1254474;
srom_1(9068) <= 1573208;
srom_1(9069) <= 1923901;
srom_1(9070) <= 2304910;
srom_1(9071) <= 2714447;
srom_1(9072) <= 3150592;
srom_1(9073) <= 3611301;
srom_1(9074) <= 4094411;
srom_1(9075) <= 4597659;
srom_1(9076) <= 5118683;
srom_1(9077) <= 5655042;
srom_1(9078) <= 6204219;
srom_1(9079) <= 6763639;
srom_1(9080) <= 7330680;
srom_1(9081) <= 7902681;
srom_1(9082) <= 8476961;
srom_1(9083) <= 9050827;
srom_1(9084) <= 9621587;
srom_1(9085) <= 10186566;
srom_1(9086) <= 10743113;
srom_1(9087) <= 11288619;
srom_1(9088) <= 11820526;
srom_1(9089) <= 12336340;
srom_1(9090) <= 12833641;
srom_1(9091) <= 13310098;
srom_1(9092) <= 13763477;
srom_1(9093) <= 14191650;
srom_1(9094) <= 14592612;
srom_1(9095) <= 14964480;
srom_1(9096) <= 15305513;
srom_1(9097) <= 15614109;
srom_1(9098) <= 15888822;
srom_1(9099) <= 16128365;
srom_1(9100) <= 16331613;
srom_1(9101) <= 16497613;
srom_1(9102) <= 16625588;
srom_1(9103) <= 16714936;
srom_1(9104) <= 16765240;
srom_1(9105) <= 16776263;
srom_1(9106) <= 16747953;
srom_1(9107) <= 16680443;
srom_1(9108) <= 16574050;
srom_1(9109) <= 16429272;
srom_1(9110) <= 16246790;
srom_1(9111) <= 16027457;
srom_1(9112) <= 15772303;
srom_1(9113) <= 15482525;
srom_1(9114) <= 15159480;
srom_1(9115) <= 14804685;
srom_1(9116) <= 14419803;
srom_1(9117) <= 14006638;
srom_1(9118) <= 13567128;
srom_1(9119) <= 13103335;
srom_1(9120) <= 12617432;
srom_1(9121) <= 12111699;
srom_1(9122) <= 11588507;
srom_1(9123) <= 11050310;
srom_1(9124) <= 10499631;
srom_1(9125) <= 9939053;
srom_1(9126) <= 9371204;
srom_1(9127) <= 8798748;
srom_1(9128) <= 8224368;
srom_1(9129) <= 7650758;
srom_1(9130) <= 7080609;
srom_1(9131) <= 6516593;
srom_1(9132) <= 5961355;
srom_1(9133) <= 5417500;
srom_1(9134) <= 4887577;
srom_1(9135) <= 4374072;
srom_1(9136) <= 3879392;
srom_1(9137) <= 3405858;
srom_1(9138) <= 2955690;
srom_1(9139) <= 2530998;
srom_1(9140) <= 2133774;
srom_1(9141) <= 1765882;
srom_1(9142) <= 1429046;
srom_1(9143) <= 1124846;
srom_1(9144) <= 854707;
srom_1(9145) <= 619898;
srom_1(9146) <= 421520;
srom_1(9147) <= 260501;
srom_1(9148) <= 137598;
srom_1(9149) <= 53387;
srom_1(9150) <= 8262;
srom_1(9151) <= 2436;
srom_1(9152) <= 35936;
srom_1(9153) <= 108604;
srom_1(9154) <= 220099;
srom_1(9155) <= 369900;
srom_1(9156) <= 557303;
srom_1(9157) <= 781430;
srom_1(9158) <= 1041230;
srom_1(9159) <= 1335484;
srom_1(9160) <= 1662812;
srom_1(9161) <= 2021680;
srom_1(9162) <= 2410405;
srom_1(9163) <= 2827163;
srom_1(9164) <= 3270001;
srom_1(9165) <= 3736842;
srom_1(9166) <= 4225497;
srom_1(9167) <= 4733674;
srom_1(9168) <= 5258990;
srom_1(9169) <= 5798982;
srom_1(9170) <= 6351118;
srom_1(9171) <= 6912808;
srom_1(9172) <= 7481418;
srom_1(9173) <= 8054283;
srom_1(9174) <= 8628716;
srom_1(9175) <= 9202022;
srom_1(9176) <= 9771514;
srom_1(9177) <= 10334522;
srom_1(9178) <= 10888404;
srom_1(9179) <= 11430564;
srom_1(9180) <= 11958459;
srom_1(9181) <= 12469613;
srom_1(9182) <= 12961631;
srom_1(9183) <= 13432204;
srom_1(9184) <= 13879126;
srom_1(9185) <= 14300301;
srom_1(9186) <= 14693753;
srom_1(9187) <= 15057639;
srom_1(9188) <= 15390252;
srom_1(9189) <= 15690031;
srom_1(9190) <= 15955572;
srom_1(9191) <= 16185628;
srom_1(9192) <= 16379122;
srom_1(9193) <= 16535145;
srom_1(9194) <= 16652967;
srom_1(9195) <= 16732034;
srom_1(9196) <= 16771975;
srom_1(9197) <= 16772605;
srom_1(9198) <= 16733918;
srom_1(9199) <= 16656098;
srom_1(9200) <= 16539509;
srom_1(9201) <= 16384697;
srom_1(9202) <= 16192389;
srom_1(9203) <= 15963486;
srom_1(9204) <= 15699062;
srom_1(9205) <= 15400357;
srom_1(9206) <= 15068771;
srom_1(9207) <= 14705860;
srom_1(9208) <= 14313325;
srom_1(9209) <= 13893007;
srom_1(9210) <= 13446876;
srom_1(9211) <= 12977026;
srom_1(9212) <= 12485660;
srom_1(9213) <= 11975080;
srom_1(9214) <= 11447683;
srom_1(9215) <= 10905940;
srom_1(9216) <= 10352393;
srom_1(9217) <= 9789637;
srom_1(9218) <= 9220311;
srom_1(9219) <= 8647085;
srom_1(9220) <= 8072647;
srom_1(9221) <= 7499690;
srom_1(9222) <= 6930902;
srom_1(9223) <= 6368950;
srom_1(9224) <= 5816468;
srom_1(9225) <= 5276048;
srom_1(9226) <= 4750224;
srom_1(9227) <= 4241461;
srom_1(9228) <= 3752146;
srom_1(9229) <= 3284573;
srom_1(9230) <= 2840935;
srom_1(9231) <= 2423311;
srom_1(9232) <= 2033661;
srom_1(9233) <= 1673811;
srom_1(9234) <= 1345449;
srom_1(9235) <= 1050115;
srom_1(9236) <= 789194;
srom_1(9237) <= 563909;
srom_1(9238) <= 375316;
srom_1(9239) <= 224301;
srom_1(9240) <= 111571;
srom_1(9241) <= 37655;
srom_1(9242) <= 2899;
srom_1(9243) <= 7467;
srom_1(9244) <= 51337;
srom_1(9245) <= 134303;
srom_1(9246) <= 255976;
srom_1(9247) <= 415786;
srom_1(9248) <= 612984;
srom_1(9249) <= 846644;
srom_1(9250) <= 1115671;
srom_1(9251) <= 1418803;
srom_1(9252) <= 1754619;
srom_1(9253) <= 2121543;
srom_1(9254) <= 2517857;
srom_1(9255) <= 2941700;
srom_1(9256) <= 3391086;
srom_1(9257) <= 3863907;
srom_1(9258) <= 4357945;
srom_1(9259) <= 4870885;
srom_1(9260) <= 5400321;
srom_1(9261) <= 5943770;
srom_1(9262) <= 6498683;
srom_1(9263) <= 7062459;
srom_1(9264) <= 7632454;
srom_1(9265) <= 8205994;
srom_1(9266) <= 8780391;
srom_1(9267) <= 9352951;
srom_1(9268) <= 9920988;
srom_1(9269) <= 10481840;
srom_1(9270) <= 11032876;
srom_1(9271) <= 11571512;
srom_1(9272) <= 12095222;
srom_1(9273) <= 12601550;
srom_1(9274) <= 13088123;
srom_1(9275) <= 13552658;
srom_1(9276) <= 13992977;
srom_1(9277) <= 14407015;
srom_1(9278) <= 14792831;
srom_1(9279) <= 15148615;
srom_1(9280) <= 15472699;
srom_1(9281) <= 15763564;
srom_1(9282) <= 16019844;
srom_1(9283) <= 16240339;
srom_1(9284) <= 16424015;
srom_1(9285) <= 16570010;
srom_1(9286) <= 16677640;
srom_1(9287) <= 16746399;
srom_1(9288) <= 16775966;
srom_1(9289) <= 16766201;
srom_1(9290) <= 16717152;
srom_1(9291) <= 16629046;
srom_1(9292) <= 16502299;
srom_1(9293) <= 16337504;
srom_1(9294) <= 16135433;
srom_1(9295) <= 15897035;
srom_1(9296) <= 15623428;
srom_1(9297) <= 15315893;
srom_1(9298) <= 14975875;
srom_1(9299) <= 14604966;
srom_1(9300) <= 14204907;
srom_1(9301) <= 13777573;
srom_1(9302) <= 13324969;
srom_1(9303) <= 12849216;
srom_1(9304) <= 12352546;
srom_1(9305) <= 11837287;
srom_1(9306) <= 11305857;
srom_1(9307) <= 10760746;
srom_1(9308) <= 10204512;
srom_1(9309) <= 9639762;
srom_1(9310) <= 9069146;
srom_1(9311) <= 8495338;
srom_1(9312) <= 7921029;
srom_1(9313) <= 7348913;
srom_1(9314) <= 6781673;
srom_1(9315) <= 6221968;
srom_1(9316) <= 5672423;
srom_1(9317) <= 5135615;
srom_1(9318) <= 4614062;
srom_1(9319) <= 4110208;
srom_1(9320) <= 3626418;
srom_1(9321) <= 3164959;
srom_1(9322) <= 2727996;
srom_1(9323) <= 2317577;
srom_1(9324) <= 1935628;
srom_1(9325) <= 1583938;
srom_1(9326) <= 1264158;
srom_1(9327) <= 977787;
srom_1(9328) <= 726168;
srom_1(9329) <= 510481;
srom_1(9330) <= 331737;
srom_1(9331) <= 190774;
srom_1(9332) <= 88254;
srom_1(9333) <= 24657;
srom_1(9334) <= 282;
srom_1(9335) <= 15242;
srom_1(9336) <= 69468;
srom_1(9337) <= 162705;
srom_1(9338) <= 294516;
srom_1(9339) <= 464283;
srom_1(9340) <= 671210;
srom_1(9341) <= 914326;
srom_1(9342) <= 1192492;
srom_1(9343) <= 1504403;
srom_1(9344) <= 1848597;
srom_1(9345) <= 2223459;
srom_1(9346) <= 2627231;
srom_1(9347) <= 3058020;
srom_1(9348) <= 3513807;
srom_1(9349) <= 3992453;
srom_1(9350) <= 4491714;
srom_1(9351) <= 5009249;
srom_1(9352) <= 5542630;
srom_1(9353) <= 6089358;
srom_1(9354) <= 6646868;
srom_1(9355) <= 7212545;
srom_1(9356) <= 7783737;
srom_1(9357) <= 8357765;
srom_1(9358) <= 8931939;
srom_1(9359) <= 9503564;
srom_1(9360) <= 10069961;
srom_1(9361) <= 10628473;
srom_1(9362) <= 11176482;
srom_1(9363) <= 11711418;
srom_1(9364) <= 12230772;
srom_1(9365) <= 12732108;
srom_1(9366) <= 13213077;
srom_1(9367) <= 13671422;
srom_1(9368) <= 14104994;
srom_1(9369) <= 14511759;
srom_1(9370) <= 14889812;
srom_1(9371) <= 15237377;
srom_1(9372) <= 15552827;
srom_1(9373) <= 15834681;
srom_1(9374) <= 16081618;
srom_1(9375) <= 16292480;
srom_1(9376) <= 16466278;
srom_1(9377) <= 16602196;
srom_1(9378) <= 16699599;
srom_1(9379) <= 16758028;
srom_1(9380) <= 16777210;
srom_1(9381) <= 16757056;
srom_1(9382) <= 16697658;
srom_1(9383) <= 16599297;
srom_1(9384) <= 16462433;
srom_1(9385) <= 16287708;
srom_1(9386) <= 16075941;
srom_1(9387) <= 15828126;
srom_1(9388) <= 15545425;
srom_1(9389) <= 15229162;
srom_1(9390) <= 14880822;
srom_1(9391) <= 14502038;
srom_1(9392) <= 14094585;
srom_1(9393) <= 13660376;
srom_1(9394) <= 13201445;
srom_1(9395) <= 12719945;
srom_1(9396) <= 12218134;
srom_1(9397) <= 11698365;
srom_1(9398) <= 11163076;
srom_1(9399) <= 10614776;
srom_1(9400) <= 10056036;
srom_1(9401) <= 9489478;
srom_1(9402) <= 8917757;
srom_1(9403) <= 8343555;
srom_1(9404) <= 7769564;
srom_1(9405) <= 7198476;
srom_1(9406) <= 6632969;
srom_1(9407) <= 6075695;
srom_1(9408) <= 5529267;
srom_1(9409) <= 4996247;
srom_1(9410) <= 4479135;
srom_1(9411) <= 3980356;
srom_1(9412) <= 3502249;
srom_1(9413) <= 3047056;
srom_1(9414) <= 2616911;
srom_1(9415) <= 2213831;
srom_1(9416) <= 1839707;
srom_1(9417) <= 1496293;
srom_1(9418) <= 1185200;
srom_1(9419) <= 907886;
srom_1(9420) <= 665651;
srom_1(9421) <= 459632;
srom_1(9422) <= 290795;
srom_1(9423) <= 159931;
srom_1(9424) <= 67654;
srom_1(9425) <= 14397;
srom_1(9426) <= 410;
srom_1(9427) <= 25758;
srom_1(9428) <= 90322;
srom_1(9429) <= 193799;
srom_1(9430) <= 335705;
srom_1(9431) <= 515374;
srom_1(9432) <= 731963;
srom_1(9433) <= 984456;
srom_1(9434) <= 1271670;
srom_1(9435) <= 1592258;
srom_1(9436) <= 1944717;
srom_1(9437) <= 2327392;
srom_1(9438) <= 2738491;
srom_1(9439) <= 3176086;
srom_1(9440) <= 3638123;
srom_1(9441) <= 4122438;
srom_1(9442) <= 4626758;
srom_1(9443) <= 5148718;
srom_1(9444) <= 5685871;
srom_1(9445) <= 6235699;
srom_1(9446) <= 6795622;
srom_1(9447) <= 7363015;
srom_1(9448) <= 7935218;
srom_1(9449) <= 8509547;
srom_1(9450) <= 9083308;
srom_1(9451) <= 9653812;
srom_1(9452) <= 10218383;
srom_1(9453) <= 10774373;
srom_1(9454) <= 11319176;
srom_1(9455) <= 11850236;
srom_1(9456) <= 12365064;
srom_1(9457) <= 12861244;
srom_1(9458) <= 13336451;
srom_1(9459) <= 13788456;
srom_1(9460) <= 14215139;
srom_1(9461) <= 14614499;
srom_1(9462) <= 14984664;
srom_1(9463) <= 15323898;
srom_1(9464) <= 15630609;
srom_1(9465) <= 15903361;
srom_1(9466) <= 16140873;
srom_1(9467) <= 16342033;
srom_1(9468) <= 16505896;
srom_1(9469) <= 16631694;
srom_1(9470) <= 16718837;
srom_1(9471) <= 16766917;
srom_1(9472) <= 16775709;
srom_1(9473) <= 16745170;
srom_1(9474) <= 16675445;
srom_1(9475) <= 16566860;
srom_1(9476) <= 16419924;
srom_1(9477) <= 16235326;
srom_1(9478) <= 16013933;
srom_1(9479) <= 15756781;
srom_1(9480) <= 15465078;
srom_1(9481) <= 15140191;
srom_1(9482) <= 14783644;
srom_1(9483) <= 14397107;
srom_1(9484) <= 13982395;
srom_1(9485) <= 13541452;
srom_1(9486) <= 13076345;
srom_1(9487) <= 12589256;
srom_1(9488) <= 12082469;
srom_1(9489) <= 11558359;
srom_1(9490) <= 11019386;
srom_1(9491) <= 10468076;
srom_1(9492) <= 9907015;
srom_1(9493) <= 9338833;
srom_1(9494) <= 8766196;
srom_1(9495) <= 8191788;
srom_1(9496) <= 7618302;
srom_1(9497) <= 7048429;
srom_1(9498) <= 6484841;
srom_1(9499) <= 5930180;
srom_1(9500) <= 5387047;
srom_1(9501) <= 4857990;
srom_1(9502) <= 4345489;
srom_1(9503) <= 3851947;
srom_1(9504) <= 3379680;
srom_1(9505) <= 2930901;
srom_1(9506) <= 2507715;
srom_1(9507) <= 2112107;
srom_1(9508) <= 1745931;
srom_1(9509) <= 1410905;
srom_1(9510) <= 1108600;
srom_1(9511) <= 840433;
srom_1(9512) <= 607663;
srom_1(9513) <= 411379;
srom_1(9514) <= 252504;
srom_1(9515) <= 131782;
srom_1(9516) <= 49779;
srom_1(9517) <= 6880;
srom_1(9518) <= 3285;
srom_1(9519) <= 39012;
srom_1(9520) <= 113893;
srom_1(9521) <= 227577;
srom_1(9522) <= 379531;
srom_1(9523) <= 569042;
srom_1(9524) <= 795222;
srom_1(9525) <= 1057010;
srom_1(9526) <= 1353178;
srom_1(9527) <= 1682338;
srom_1(9528) <= 2042946;
srom_1(9529) <= 2433311;
srom_1(9530) <= 2851602;
srom_1(9531) <= 3295858;
srom_1(9532) <= 3763996;
srom_1(9533) <= 4253820;
srom_1(9534) <= 4763033;
srom_1(9535) <= 5289248;
srom_1(9536) <= 5829997;
srom_1(9537) <= 6382745;
srom_1(9538) <= 6944898;
srom_1(9539) <= 7513822;
srom_1(9540) <= 8086847;
srom_1(9541) <= 8661288;
srom_1(9542) <= 9234450;
srom_1(9543) <= 9803646;
srom_1(9544) <= 10366206;
srom_1(9545) <= 10919492;
srom_1(9546) <= 11460910;
srom_1(9547) <= 11987921;
srom_1(9548) <= 12498054;
srom_1(9549) <= 12988916;
srom_1(9550) <= 13458205;
srom_1(9551) <= 13903722;
srom_1(9552) <= 14323376;
srom_1(9553) <= 14715200;
srom_1(9554) <= 15077357;
srom_1(9555) <= 15408147;
srom_1(9556) <= 15706021;
srom_1(9557) <= 15969581;
srom_1(9558) <= 16197591;
srom_1(9559) <= 16388981;
srom_1(9560) <= 16542856;
srom_1(9561) <= 16658492;
srom_1(9562) <= 16735348;
srom_1(9563) <= 16773063;
srom_1(9564) <= 16771461;
srom_1(9565) <= 16730549;
srom_1(9566) <= 16650518;
srom_1(9567) <= 16531744;
srom_1(9568) <= 16374785;
srom_1(9569) <= 16180375;
srom_1(9570) <= 15949428;
srom_1(9571) <= 15683025;
srom_1(9572) <= 15382415;
srom_1(9573) <= 15049010;
srom_1(9574) <= 14684372;
srom_1(9575) <= 14290210;
srom_1(9576) <= 13868374;
srom_1(9577) <= 13420842;
srom_1(9578) <= 12949711;
srom_1(9579) <= 12457192;
srom_1(9580) <= 11945594;
srom_1(9581) <= 11417316;
srom_1(9582) <= 10874835;
srom_1(9583) <= 10320696;
srom_1(9584) <= 9757496;
srom_1(9585) <= 9187878;
srom_1(9586) <= 8614511;
srom_1(9587) <= 8040084;
srom_1(9588) <= 7467293;
srom_1(9589) <= 6898821;
srom_1(9590) <= 6337336;
srom_1(9591) <= 5785469;
srom_1(9592) <= 5245810;
srom_1(9593) <= 4720888;
srom_1(9594) <= 4213166;
srom_1(9595) <= 3725024;
srom_1(9596) <= 3258750;
srom_1(9597) <= 2816533;
srom_1(9598) <= 2400445;
srom_1(9599) <= 2012437;
srom_1(9600) <= 1654329;
srom_1(9601) <= 1327801;
srom_1(9602) <= 1034383;
srom_1(9603) <= 775452;
srom_1(9604) <= 552221;
srom_1(9605) <= 365738;
srom_1(9606) <= 216877;
srom_1(9607) <= 106336;
srom_1(9608) <= 34634;
srom_1(9609) <= 2106;
srom_1(9610) <= 8905;
srom_1(9611) <= 54999;
srom_1(9612) <= 140173;
srom_1(9613) <= 264027;
srom_1(9614) <= 425979;
srom_1(9615) <= 625271;
srom_1(9616) <= 860968;
srom_1(9617) <= 1131964;
srom_1(9618) <= 1436989;
srom_1(9619) <= 1774613;
srom_1(9620) <= 2143253;
srom_1(9621) <= 2541178;
srom_1(9622) <= 2966525;
srom_1(9623) <= 3417297;
srom_1(9624) <= 3891382;
srom_1(9625) <= 4386555;
srom_1(9626) <= 4900496;
srom_1(9627) <= 5430793;
srom_1(9628) <= 5974961;
srom_1(9629) <= 6530447;
srom_1(9630) <= 7094647;
srom_1(9631) <= 7664915;
srom_1(9632) <= 8238576;
srom_1(9633) <= 8812940;
srom_1(9634) <= 9385315;
srom_1(9635) <= 9953016;
srom_1(9636) <= 10513381;
srom_1(9637) <= 11063782;
srom_1(9638) <= 11601639;
srom_1(9639) <= 12124428;
srom_1(9640) <= 12629699;
srom_1(9641) <= 13115081;
srom_1(9642) <= 13578300;
srom_1(9643) <= 14017183;
srom_1(9644) <= 14429671;
srom_1(9645) <= 14813830;
srom_1(9646) <= 15167860;
srom_1(9647) <= 15490099;
srom_1(9648) <= 15779037;
srom_1(9649) <= 16033318;
srom_1(9650) <= 16251751;
srom_1(9651) <= 16433311;
srom_1(9652) <= 16577147;
srom_1(9653) <= 16682583;
srom_1(9654) <= 16749127;
srom_1(9655) <= 16776465;
srom_1(9656) <= 16764469;
srom_1(9657) <= 16713196;
srom_1(9658) <= 16622886;
srom_1(9659) <= 16493963;
srom_1(9660) <= 16327032;
srom_1(9661) <= 16122874;
srom_1(9662) <= 15882447;
srom_1(9663) <= 15606879;
srom_1(9664) <= 15297463;
srom_1(9665) <= 14955648;
srom_1(9666) <= 14583038;
srom_1(9667) <= 14181381;
srom_1(9668) <= 13752559;
srom_1(9669) <= 13298583;
srom_1(9670) <= 12821584;
srom_1(9671) <= 12323796;
srom_1(9672) <= 11807555;
srom_1(9673) <= 11275281;
srom_1(9674) <= 10729471;
srom_1(9675) <= 10172683;
srom_1(9676) <= 9607530;
srom_1(9677) <= 9036660;
srom_1(9678) <= 8462752;
srom_1(9679) <= 7888495;
srom_1(9680) <= 7316584;
srom_1(9681) <= 6749700;
srom_1(9682) <= 6190502;
srom_1(9683) <= 5641611;
srom_1(9684) <= 5105602;
srom_1(9685) <= 4584988;
srom_1(9686) <= 4082210;
srom_1(9687) <= 3599627;
srom_1(9688) <= 3139500;
srom_1(9689) <= 2703989;
srom_1(9690) <= 2295135;
srom_1(9691) <= 1914855;
srom_1(9692) <= 1564932;
srom_1(9693) <= 1247009;
srom_1(9694) <= 962574;
srom_1(9695) <= 712963;
srom_1(9696) <= 499346;
srom_1(9697) <= 322724;
srom_1(9698) <= 183926;
srom_1(9699) <= 83602;
srom_1(9700) <= 22223;
srom_1(9701) <= 78;
srom_1(9702) <= 17269;
srom_1(9703) <= 73715;
srom_1(9704) <= 169154;
srom_1(9705) <= 303136;
srom_1(9706) <= 475034;
srom_1(9707) <= 684041;
srom_1(9708) <= 929178;
srom_1(9709) <= 1209294;
srom_1(9710) <= 1523077;
srom_1(9711) <= 1869054;
srom_1(9712) <= 2245604;
srom_1(9713) <= 2650961;
srom_1(9714) <= 3083223;
srom_1(9715) <= 3540364;
srom_1(9716) <= 4020240;
srom_1(9717) <= 4520601;
srom_1(9718) <= 5039100;
srom_1(9719) <= 5573307;
srom_1(9720) <= 6120715;
srom_1(9721) <= 6678758;
srom_1(9722) <= 7244819;
srom_1(9723) <= 7816244;
srom_1(9724) <= 8390353;
srom_1(9725) <= 8964454;
srom_1(9726) <= 9535854;
srom_1(9727) <= 10101875;
srom_1(9728) <= 10659861;
srom_1(9729) <= 11207197;
srom_1(9730) <= 11741315;
srom_1(9731) <= 12259711;
srom_1(9732) <= 12759955;
srom_1(9733) <= 13239699;
srom_1(9734) <= 13696696;
srom_1(9735) <= 14128800;
srom_1(9736) <= 14533987;
srom_1(9737) <= 14910357;
srom_1(9738) <= 15256143;
srom_1(9739) <= 15569725;
srom_1(9740) <= 15849633;
srom_1(9741) <= 16094553;
srom_1(9742) <= 16303337;
srom_1(9743) <= 16475007;
srom_1(9744) <= 16608756;
srom_1(9745) <= 16703959;
srom_1(9746) <= 16760168;
srom_1(9747) <= 16777120;
srom_1(9748) <= 16754735;
srom_1(9749) <= 16693118;
srom_1(9750) <= 16592559;
srom_1(9751) <= 16453529;
srom_1(9752) <= 16276679;
srom_1(9753) <= 16062840;
srom_1(9754) <= 15813013;
srom_1(9755) <= 15528371;
srom_1(9756) <= 15210248;
srom_1(9757) <= 14860136;
srom_1(9758) <= 14479677;
srom_1(9759) <= 14070655;
srom_1(9760) <= 13634987;
srom_1(9761) <= 13174718;
srom_1(9762) <= 12692005;
srom_1(9763) <= 12189111;
srom_1(9764) <= 11668396;
srom_1(9765) <= 11132301;
srom_1(9766) <= 10583340;
srom_1(9767) <= 10024086;
srom_1(9768) <= 9457164;
srom_1(9769) <= 8885230;
srom_1(9770) <= 8310968;
srom_1(9771) <= 7737070;
srom_1(9772) <= 7166227;
srom_1(9773) <= 6601117;
srom_1(9774) <= 6044388;
srom_1(9775) <= 5498652;
srom_1(9776) <= 4966469;
srom_1(9777) <= 4450332;
srom_1(9778) <= 3952664;
srom_1(9779) <= 3475798;
srom_1(9780) <= 3021969;
srom_1(9781) <= 2593306;
srom_1(9782) <= 2191820;
srom_1(9783) <= 1819392;
srom_1(9784) <= 1477770;
srom_1(9785) <= 1168554;
srom_1(9786) <= 893197;
srom_1(9787) <= 652987;
srom_1(9788) <= 449053;
srom_1(9789) <= 282350;
srom_1(9790) <= 153660;
srom_1(9791) <= 63587;
srom_1(9792) <= 12552;
srom_1(9793) <= 796;
srom_1(9794) <= 28373;
srom_1(9795) <= 95154;
srom_1(9796) <= 200826;
srom_1(9797) <= 344893;
srom_1(9798) <= 526679;
srom_1(9799) <= 745334;
srom_1(9800) <= 999830;
srom_1(9801) <= 1288974;
srom_1(9802) <= 1611411;
srom_1(9803) <= 1965629;
srom_1(9804) <= 2349967;
srom_1(9805) <= 2762621;
srom_1(9806) <= 3201658;
srom_1(9807) <= 3665018;
srom_1(9808) <= 4150529;
srom_1(9809) <= 4655913;
srom_1(9810) <= 5178802;
srom_1(9811) <= 5716742;
srom_1(9812) <= 6267211;
srom_1(9813) <= 6827629;
srom_1(9814) <= 7395366;
srom_1(9815) <= 7967761;
srom_1(9816) <= 8542130;
srom_1(9817) <= 9115779;
srom_1(9818) <= 9686017;
srom_1(9819) <= 10250172;
srom_1(9820) <= 10805597;
srom_1(9821) <= 11349688;
srom_1(9822) <= 11879894;
srom_1(9823) <= 12393728;
srom_1(9824) <= 12888780;
srom_1(9825) <= 13362729;
srom_1(9826) <= 13813353;
srom_1(9827) <= 14238539;
srom_1(9828) <= 14636292;
srom_1(9829) <= 15004748;
srom_1(9830) <= 15342178;
srom_1(9831) <= 15647001;
srom_1(9832) <= 15917786;
srom_1(9833) <= 16153265;
srom_1(9834) <= 16352332;
srom_1(9835) <= 16514055;
srom_1(9836) <= 16637675;
srom_1(9837) <= 16722612;
srom_1(9838) <= 16768468;
srom_1(9839) <= 16775028;
srom_1(9840) <= 16742261;
srom_1(9841) <= 16670322;
srom_1(9842) <= 16559546;
srom_1(9843) <= 16410454;
srom_1(9844) <= 16223744;
srom_1(9845) <= 16000293;
srom_1(9846) <= 15741149;
srom_1(9847) <= 15447525;
srom_1(9848) <= 15120800;
srom_1(9849) <= 14762506;
srom_1(9850) <= 14374322;
srom_1(9851) <= 13958068;
srom_1(9852) <= 13515698;
srom_1(9853) <= 13049285;
srom_1(9854) <= 12561017;
srom_1(9855) <= 12053183;
srom_1(9856) <= 11528164;
srom_1(9857) <= 10988423;
srom_1(9858) <= 10436490;
srom_1(9859) <= 9874954;
srom_1(9860) <= 9306448;
srom_1(9861) <= 8733638;
srom_1(9862) <= 8159210;
srom_1(9863) <= 7585858;
srom_1(9864) <= 7016270;
srom_1(9865) <= 6453118;
srom_1(9866) <= 5899041;
srom_1(9867) <= 5356640;
srom_1(9868) <= 4828456;
srom_1(9869) <= 4316966;
srom_1(9870) <= 3824571;
srom_1(9871) <= 3353577;
srom_1(9872) <= 2906194;
srom_1(9873) <= 2484521;
srom_1(9874) <= 2090533;
srom_1(9875) <= 1726080;
srom_1(9876) <= 1392869;
srom_1(9877) <= 1092464;
srom_1(9878) <= 826273;
srom_1(9879) <= 595544;
srom_1(9880) <= 401360;
srom_1(9881) <= 244630;
srom_1(9882) <= 126091;
srom_1(9883) <= 46297;
srom_1(9884) <= 5623;
srom_1(9885) <= 4260;
srom_1(9886) <= 42214;
srom_1(9887) <= 119307;
srom_1(9888) <= 235178;
srom_1(9889) <= 389283;
srom_1(9890) <= 580899;
srom_1(9891) <= 809129;
srom_1(9892) <= 1072901;
srom_1(9893) <= 1370979;
srom_1(9894) <= 1701965;
srom_1(9895) <= 2064307;
srom_1(9896) <= 2456306;
srom_1(9897) <= 2876124;
srom_1(9898) <= 3321791;
srom_1(9899) <= 3791219;
srom_1(9900) <= 4282205;
srom_1(9901) <= 4792447;
srom_1(9902) <= 5319554;
srom_1(9903) <= 5861052;
srom_1(9904) <= 6414402;
srom_1(9905) <= 6977011;
srom_1(9906) <= 7546238;
srom_1(9907) <= 8119416;
srom_1(9908) <= 8693857;
srom_1(9909) <= 9266865;
srom_1(9910) <= 9835756;
srom_1(9911) <= 10397860;
srom_1(9912) <= 10950542;
srom_1(9913) <= 11491210;
srom_1(9914) <= 12017330;
srom_1(9915) <= 12526432;
srom_1(9916) <= 13016132;
srom_1(9917) <= 13484131;
srom_1(9918) <= 13928235;
srom_1(9919) <= 14346362;
srom_1(9920) <= 14736551;
srom_1(9921) <= 15096973;
srom_1(9922) <= 15425937;
srom_1(9923) <= 15721900;
srom_1(9924) <= 15983475;
srom_1(9925) <= 16209435;
srom_1(9926) <= 16398720;
srom_1(9927) <= 16550443;
srom_1(9928) <= 16663893;
srom_1(9929) <= 16738537;
srom_1(9930) <= 16774025;
srom_1(9931) <= 16770191;
srom_1(9932) <= 16727053;
srom_1(9933) <= 16644813;
srom_1(9934) <= 16523857;
srom_1(9935) <= 16364752;
srom_1(9936) <= 16168244;
srom_1(9937) <= 15935255;
srom_1(9938) <= 15666877;
srom_1(9939) <= 15364368;
srom_1(9940) <= 15029148;
srom_1(9941) <= 14662788;
srom_1(9942) <= 14267006;
srom_1(9943) <= 13843659;
srom_1(9944) <= 13394731;
srom_1(9945) <= 12922327;
srom_1(9946) <= 12428663;
srom_1(9947) <= 11916054;
srom_1(9948) <= 11386904;
srom_1(9949) <= 10843693;
srom_1(9950) <= 10288970;
srom_1(9951) <= 9725335;
srom_1(9952) <= 9155432;
srom_1(9953) <= 8581933;
srom_1(9954) <= 8007527;
srom_1(9955) <= 7434909;
srom_1(9956) <= 6866763;
srom_1(9957) <= 6305753;
srom_1(9958) <= 5754510;
srom_1(9959) <= 5215619;
srom_1(9960) <= 4691608;
srom_1(9961) <= 4184933;
srom_1(9962) <= 3697971;
srom_1(9963) <= 3233005;
srom_1(9964) <= 2792215;
srom_1(9965) <= 2377668;
srom_1(9966) <= 1991309;
srom_1(9967) <= 1634949;
srom_1(9968) <= 1310259;
srom_1(9969) <= 1018762;
srom_1(9970) <= 761825;
srom_1(9971) <= 540652;
srom_1(9972) <= 356281;
srom_1(9973) <= 209577;
srom_1(9974) <= 101226;
srom_1(9975) <= 31739;
srom_1(9976) <= 1439;
srom_1(9977) <= 10469;
srom_1(9978) <= 58788;
srom_1(9979) <= 146168;
srom_1(9980) <= 272199;
srom_1(9981) <= 436292;
srom_1(9982) <= 637675;
srom_1(9983) <= 875405;
srom_1(9984) <= 1148367;
srom_1(9985) <= 1455281;
srom_1(9986) <= 1794708;
srom_1(9987) <= 2165056;
srom_1(9988) <= 2564588;
srom_1(9989) <= 2991431;
srom_1(9990) <= 3443583;
srom_1(9991) <= 3918924;
srom_1(9992) <= 4415225;
srom_1(9993) <= 4930159;
srom_1(9994) <= 5461311;
srom_1(9995) <= 6006189;
srom_1(9996) <= 6562240;
srom_1(9997) <= 7126855;
srom_1(9998) <= 7697386;
srom_1(9999) <= 8271159;
srom_1(10000) <= 8845483;
srom_1(10001) <= 9417665;
srom_1(10002) <= 9985021;
srom_1(10003) <= 10544890;
srom_1(10004) <= 11094648;
srom_1(10005) <= 11631717;
srom_1(10006) <= 12153577;
srom_1(10007) <= 12657783;
srom_1(10008) <= 13141968;
srom_1(10009) <= 13603864;
srom_1(10010) <= 14041303;
srom_1(10011) <= 14452235;
srom_1(10012) <= 14834733;
srom_1(10013) <= 15187002;
srom_1(10014) <= 15507391;
srom_1(10015) <= 15794398;
srom_1(10016) <= 16046677;
srom_1(10017) <= 16263044;
srom_1(10018) <= 16442486;
srom_1(10019) <= 16584159;
srom_1(10020) <= 16687402;
srom_1(10021) <= 16751728;
srom_1(10022) <= 16776837;
srom_1(10023) <= 16762610;
srom_1(10024) <= 16709115;
srom_1(10025) <= 16616602;
srom_1(10026) <= 16485505;
srom_1(10027) <= 16316440;
srom_1(10028) <= 16110197;
srom_1(10029) <= 15867746;
srom_1(10030) <= 15590222;
srom_1(10031) <= 15278928;
srom_1(10032) <= 14935322;
srom_1(10033) <= 14561017;
srom_1(10034) <= 14157767;
srom_1(10035) <= 13727463;
srom_1(10036) <= 13272124;
srom_1(10037) <= 12793884;
srom_1(10038) <= 12294987;
srom_1(10039) <= 11777771;
srom_1(10040) <= 11244662;
srom_1(10041) <= 10698160;
srom_1(10042) <= 10140828;
srom_1(10043) <= 9575279;
srom_1(10044) <= 9004165;
srom_1(10045) <= 8430165;
srom_1(10046) <= 7855969;
srom_1(10047) <= 7284272;
srom_1(10048) <= 6717753;
srom_1(10049) <= 6159069;
srom_1(10050) <= 5610841;
srom_1(10051) <= 5075638;
srom_1(10052) <= 4555971;
srom_1(10053) <= 4054277;
srom_1(10054) <= 3572907;
srom_1(10055) <= 3114121;
srom_1(10056) <= 2680068;
srom_1(10057) <= 2272784;
srom_1(10058) <= 1894179;
srom_1(10059) <= 1546029;
srom_1(10060) <= 1229967;
srom_1(10061) <= 947473;
srom_1(10062) <= 699874;
srom_1(10063) <= 488330;
srom_1(10064) <= 313833;
srom_1(10065) <= 177201;
srom_1(10066) <= 79075;
srom_1(10067) <= 19916;
srom_1(10068) <= 0;
srom_1(10069) <= 19422;
srom_1(10070) <= 78089;
srom_1(10071) <= 175727;
srom_1(10072) <= 311878;
srom_1(10073) <= 485904;
srom_1(10074) <= 696988;
srom_1(10075) <= 944141;
srom_1(10076) <= 1226204;
srom_1(10077) <= 1541853;
srom_1(10078) <= 1889610;
srom_1(10079) <= 2267842;
srom_1(10080) <= 2674777;
srom_1(10081) <= 3108505;
srom_1(10082) <= 3566994;
srom_1(10083) <= 4048094;
srom_1(10084) <= 4549547;
srom_1(10085) <= 5069003;
srom_1(10086) <= 5604026;
srom_1(10087) <= 6152106;
srom_1(10088) <= 6710675;
srom_1(10089) <= 7277111;
srom_1(10090) <= 7848760;
srom_1(10091) <= 8422941;
srom_1(10092) <= 8996960;
srom_1(10093) <= 9568127;
srom_1(10094) <= 10133763;
srom_1(10095) <= 10691214;
srom_1(10096) <= 11237869;
srom_1(10097) <= 11771162;
srom_1(10098) <= 12288593;
srom_1(10099) <= 12787735;
srom_1(10100) <= 13266249;
srom_1(10101) <= 13721889;
srom_1(10102) <= 14152521;
srom_1(10103) <= 14556123;
srom_1(10104) <= 14930803;
srom_1(10105) <= 15274805;
srom_1(10106) <= 15586515;
srom_1(10107) <= 15864472;
srom_1(10108) <= 16107372;
srom_1(10109) <= 16314075;
srom_1(10110) <= 16483614;
srom_1(10111) <= 16615192;
srom_1(10112) <= 16708193;
srom_1(10113) <= 16762181;
srom_1(10114) <= 16776902;
srom_1(10115) <= 16752288;
srom_1(10116) <= 16688453;
srom_1(10117) <= 16585697;
srom_1(10118) <= 16444503;
srom_1(10119) <= 16265531;
srom_1(10120) <= 16049622;
srom_1(10121) <= 15797788;
srom_1(10122) <= 15511210;
srom_1(10123) <= 15191231;
srom_1(10124) <= 14839353;
srom_1(10125) <= 14457224;
srom_1(10126) <= 14046638;
srom_1(10127) <= 13609520;
srom_1(10128) <= 13147919;
srom_1(10129) <= 12663999;
srom_1(10130) <= 12160031;
srom_1(10131) <= 11638378;
srom_1(10132) <= 11101485;
srom_1(10133) <= 10551870;
srom_1(10134) <= 9992112;
srom_1(10135) <= 9424833;
srom_1(10136) <= 8852696;
srom_1(10137) <= 8278382;
srom_1(10138) <= 7704586;
srom_1(10139) <= 7133997;
srom_1(10140) <= 6569291;
srom_1(10141) <= 6013116;
srom_1(10142) <= 5468081;
srom_1(10143) <= 4936742;
srom_1(10144) <= 4421589;
srom_1(10145) <= 3925039;
srom_1(10146) <= 3449420;
srom_1(10147) <= 2996963;
srom_1(10148) <= 2569789;
srom_1(10149) <= 2169902;
srom_1(10150) <= 1799176;
srom_1(10151) <= 1459350;
srom_1(10152) <= 1152018;
srom_1(10153) <= 878621;
srom_1(10154) <= 640440;
srom_1(10155) <= 438594;
srom_1(10156) <= 274028;
srom_1(10157) <= 147514;
srom_1(10158) <= 59645;
srom_1(10159) <= 10833;
srom_1(10160) <= 1308;
srom_1(10161) <= 31114;
srom_1(10162) <= 100111;
srom_1(10163) <= 207975;
srom_1(10164) <= 354201;
srom_1(10165) <= 538104;
srom_1(10166) <= 758820;
srom_1(10167) <= 1015315;
srom_1(10168) <= 1306385;
srom_1(10169) <= 1630667;
srom_1(10170) <= 1986639;
srom_1(10171) <= 2372632;
srom_1(10172) <= 2786836;
srom_1(10173) <= 3227308;
srom_1(10174) <= 3691984;
srom_1(10175) <= 4178684;
srom_1(10176) <= 4685125;
srom_1(10177) <= 5208934;
srom_1(10178) <= 5747653;
srom_1(10179) <= 6298756;
srom_1(10180) <= 6859659;
srom_1(10181) <= 7427732;
srom_1(10182) <= 8000311;
srom_1(10183) <= 8574711;
srom_1(10184) <= 9148238;
srom_1(10185) <= 9718203;
srom_1(10186) <= 10281933;
srom_1(10187) <= 10836785;
srom_1(10188) <= 11380156;
srom_1(10189) <= 11909499;
srom_1(10190) <= 12422331;
srom_1(10191) <= 12916247;
srom_1(10192) <= 13388932;
srom_1(10193) <= 13838169;
srom_1(10194) <= 14261851;
srom_1(10195) <= 14657991;
srom_1(10196) <= 15024732;
srom_1(10197) <= 15360354;
srom_1(10198) <= 15663283;
srom_1(10199) <= 15932098;
srom_1(10200) <= 16165539;
srom_1(10201) <= 16362512;
srom_1(10202) <= 16522092;
srom_1(10203) <= 16643532;
srom_1(10204) <= 16726261;
srom_1(10205) <= 16769893;
srom_1(10206) <= 16774221;
srom_1(10207) <= 16739227;
srom_1(10208) <= 16665073;
srom_1(10209) <= 16552109;
srom_1(10210) <= 16400863;
srom_1(10211) <= 16212044;
srom_1(10212) <= 15986539;
srom_1(10213) <= 15725405;
srom_1(10214) <= 15429866;
srom_1(10215) <= 15101308;
srom_1(10216) <= 14741271;
srom_1(10217) <= 14351445;
srom_1(10218) <= 13933658;
srom_1(10219) <= 13489867;
srom_1(10220) <= 13022155;
srom_1(10221) <= 12532715;
srom_1(10222) <= 12023841;
srom_1(10223) <= 11497921;
srom_1(10224) <= 10957420;
srom_1(10225) <= 10404873;
srom_1(10226) <= 9842871;
srom_1(10227) <= 9274049;
srom_1(10228) <= 8701075;
srom_1(10229) <= 8126636;
srom_1(10230) <= 7553426;
srom_1(10231) <= 6984132;
srom_1(10232) <= 6421424;
srom_1(10233) <= 5867941;
srom_1(10234) <= 5326278;
srom_1(10235) <= 4798975;
srom_1(10236) <= 4288505;
srom_1(10237) <= 3797263;
srom_1(10238) <= 3327550;
srom_1(10239) <= 2881571;
srom_1(10240) <= 2461416;
srom_1(10241) <= 2069055;
srom_1(10242) <= 1706330;
srom_1(10243) <= 1374939;
srom_1(10244) <= 1076438;
srom_1(10245) <= 812227;
srom_1(10246) <= 583543;
srom_1(10247) <= 391461;
srom_1(10248) <= 236879;
srom_1(10249) <= 120524;
srom_1(10250) <= 42941;
srom_1(10251) <= 4493;
srom_1(10252) <= 5362;
srom_1(10253) <= 45542;
srom_1(10254) <= 124846;
srom_1(10255) <= 242902;
srom_1(10256) <= 399155;
srom_1(10257) <= 592874;
srom_1(10258) <= 823149;
srom_1(10259) <= 1088902;
srom_1(10260) <= 1388886;
srom_1(10261) <= 1721693;
srom_1(10262) <= 2085764;
srom_1(10263) <= 2479391;
srom_1(10264) <= 2900729;
srom_1(10265) <= 3347801;
srom_1(10266) <= 3818511;
srom_1(10267) <= 4310652;
srom_1(10268) <= 4821916;
srom_1(10269) <= 5349905;
srom_1(10270) <= 5892144;
srom_1(10271) <= 6446090;
srom_1(10272) <= 7009144;
srom_1(10273) <= 7578668;
srom_1(10274) <= 8151989;
srom_1(10275) <= 8726420;
srom_1(10276) <= 9299267;
srom_1(10277) <= 9867844;
srom_1(10278) <= 10429484;
srom_1(10279) <= 10981554;
srom_1(10280) <= 11521464;
srom_1(10281) <= 12046683;
srom_1(10282) <= 12554749;
srom_1(10283) <= 13043277;
srom_1(10284) <= 13509979;
srom_1(10285) <= 13952665;
srom_1(10286) <= 14369258;
srom_1(10287) <= 14757807;
srom_1(10288) <= 15116488;
srom_1(10289) <= 15443620;
srom_1(10290) <= 15737668;
srom_1(10291) <= 15997254;
srom_1(10292) <= 16221161;
srom_1(10293) <= 16408338;
srom_1(10294) <= 16557908;
srom_1(10295) <= 16669169;
srom_1(10296) <= 16741600;
srom_1(10297) <= 16774860;
srom_1(10298) <= 16768795;
srom_1(10299) <= 16723432;
srom_1(10300) <= 16638984;
srom_1(10301) <= 16515847;
srom_1(10302) <= 16354599;
srom_1(10303) <= 16155996;
srom_1(10304) <= 15920969;
srom_1(10305) <= 15650619;
srom_1(10306) <= 15346216;
srom_1(10307) <= 15009186;
srom_1(10308) <= 14641110;
srom_1(10309) <= 14243714;
srom_1(10310) <= 13818861;
srom_1(10311) <= 13368544;
srom_1(10312) <= 12894874;
srom_1(10313) <= 12400073;
srom_1(10314) <= 11886461;
srom_1(10315) <= 11356446;
srom_1(10316) <= 10812514;
srom_1(10317) <= 10257215;
srom_1(10318) <= 9693154;
srom_1(10319) <= 9122975;
srom_1(10320) <= 8549352;
srom_1(10321) <= 7974976;
srom_1(10322) <= 7402540;
srom_1(10323) <= 6834727;
srom_1(10324) <= 6274201;
srom_1(10325) <= 5723590;
srom_1(10326) <= 5185477;
srom_1(10327) <= 4662384;
srom_1(10328) <= 4156764;
srom_1(10329) <= 3670989;
srom_1(10330) <= 3207337;
srom_1(10331) <= 2767981;
srom_1(10332) <= 2354983;
srom_1(10333) <= 1970278;
srom_1(10334) <= 1615671;
srom_1(10335) <= 1292825;
srom_1(10336) <= 1003253;
srom_1(10337) <= 748313;
srom_1(10338) <= 529202;
srom_1(10339) <= 346946;
srom_1(10340) <= 202400;
srom_1(10341) <= 96242;
srom_1(10342) <= 28969;
srom_1(10343) <= 898;
srom_1(10344) <= 12160;
srom_1(10345) <= 62702;
srom_1(10346) <= 152287;
srom_1(10347) <= 280495;
srom_1(10348) <= 446724;
srom_1(10349) <= 650196;
srom_1(10350) <= 889956;
srom_1(10351) <= 1164879;
srom_1(10352) <= 1473677;
srom_1(10353) <= 1814902;
srom_1(10354) <= 2186953;
srom_1(10355) <= 2588086;
srom_1(10356) <= 3016419;
srom_1(10357) <= 3469944;
srom_1(10358) <= 3946535;
srom_1(10359) <= 4443956;
srom_1(10360) <= 4959874;
srom_1(10361) <= 5491872;
srom_1(10362) <= 6037453;
srom_1(10363) <= 6594059;
srom_1(10364) <= 7159081;
srom_1(10365) <= 7729868;
srom_1(10366) <= 8303745;
srom_1(10367) <= 8878019;
srom_1(10368) <= 9449999;
srom_1(10369) <= 10017001;
srom_1(10370) <= 10576367;
srom_1(10371) <= 11125474;
srom_1(10372) <= 11661746;
srom_1(10373) <= 12182670;
srom_1(10374) <= 12685802;
srom_1(10375) <= 13168783;
srom_1(10376) <= 13629349;
srom_1(10377) <= 14065338;
srom_1(10378) <= 14474708;
srom_1(10379) <= 14855538;
srom_1(10380) <= 15206042;
srom_1(10381) <= 15524576;
srom_1(10382) <= 15809648;
srom_1(10383) <= 16059920;
srom_1(10384) <= 16274218;
srom_1(10385) <= 16451538;
srom_1(10386) <= 16591049;
srom_1(10387) <= 16692095;
srom_1(10388) <= 16754203;
srom_1(10389) <= 16777082;
srom_1(10390) <= 16760625;
srom_1(10391) <= 16704908;
srom_1(10392) <= 16610194;
srom_1(10393) <= 16476925;
srom_1(10394) <= 16305728;
srom_1(10395) <= 16097405;
srom_1(10396) <= 15852932;
srom_1(10397) <= 15573456;
srom_1(10398) <= 15260289;
srom_1(10399) <= 14914897;
srom_1(10400) <= 14538902;
srom_1(10401) <= 14134066;
srom_1(10402) <= 13702287;
srom_1(10403) <= 13245591;
srom_1(10404) <= 12766119;
srom_1(10405) <= 12266119;
srom_1(10406) <= 11747935;
srom_1(10407) <= 11213999;
srom_1(10408) <= 10666814;
srom_1(10409) <= 10108945;
srom_1(10410) <= 9543010;
srom_1(10411) <= 8971660;
srom_1(10412) <= 8397577;
srom_1(10413) <= 7823451;
srom_1(10414) <= 7251976;
srom_1(10415) <= 6685831;
srom_1(10416) <= 6127671;
srom_1(10417) <= 5580113;
srom_1(10418) <= 5045725;
srom_1(10419) <= 4527012;
srom_1(10420) <= 4026409;
srom_1(10421) <= 3546261;
srom_1(10422) <= 3088820;
srom_1(10423) <= 2656232;
srom_1(10424) <= 2250525;
srom_1(10425) <= 1873602;
srom_1(10426) <= 1527230;
srom_1(10427) <= 1213033;
srom_1(10428) <= 932485;
srom_1(10429) <= 686901;
srom_1(10430) <= 477433;
srom_1(10431) <= 305063;
srom_1(10432) <= 170600;
srom_1(10433) <= 74674;
srom_1(10434) <= 17735;
srom_1(10435) <= 50;
srom_1(10436) <= 21701;
srom_1(10437) <= 82588;
srom_1(10438) <= 182424;
srom_1(10439) <= 320743;
srom_1(10440) <= 496894;
srom_1(10441) <= 710052;
srom_1(10442) <= 959217;
srom_1(10443) <= 1243222;
srom_1(10444) <= 1560733;
srom_1(10445) <= 1910263;
srom_1(10446) <= 2290172;
srom_1(10447) <= 2698679;
srom_1(10448) <= 3133868;
srom_1(10449) <= 3593698;
srom_1(10450) <= 4076012;
srom_1(10451) <= 4578551;
srom_1(10452) <= 5098956;
srom_1(10453) <= 5634787;
srom_1(10454) <= 6183531;
srom_1(10455) <= 6742617;
srom_1(10456) <= 7309420;
srom_1(10457) <= 7881285;
srom_1(10458) <= 8455528;
srom_1(10459) <= 9029458;
srom_1(10460) <= 9600382;
srom_1(10461) <= 10165624;
srom_1(10462) <= 10722533;
srom_1(10463) <= 11268497;
srom_1(10464) <= 11800957;
srom_1(10465) <= 12317415;
srom_1(10466) <= 12815449;
srom_1(10467) <= 13292725;
srom_1(10468) <= 13747003;
srom_1(10469) <= 14176154;
srom_1(10470) <= 14578165;
srom_1(10471) <= 14951151;
srom_1(10472) <= 15293363;
srom_1(10473) <= 15603196;
srom_1(10474) <= 15879198;
srom_1(10475) <= 16120074;
srom_1(10476) <= 16324694;
srom_1(10477) <= 16492099;
srom_1(10478) <= 16621504;
srom_1(10479) <= 16712302;
srom_1(10480) <= 16764068;
srom_1(10481) <= 16776558;
srom_1(10482) <= 16749714;
srom_1(10483) <= 16683662;
srom_1(10484) <= 16578712;
srom_1(10485) <= 16435355;
srom_1(10486) <= 16254265;
srom_1(10487) <= 16036289;
srom_1(10488) <= 15782451;
srom_1(10489) <= 15493941;
srom_1(10490) <= 15172112;
srom_1(10491) <= 14818472;
srom_1(10492) <= 14434680;
srom_1(10493) <= 14022537;
srom_1(10494) <= 13583974;
srom_1(10495) <= 13121048;
srom_1(10496) <= 12635929;
srom_1(10497) <= 12130894;
srom_1(10498) <= 11608310;
srom_1(10499) <= 11070628;
srom_1(10500) <= 10520369;
srom_1(10501) <= 9960113;
srom_1(10502) <= 9392488;
srom_1(10503) <= 8820155;
srom_1(10504) <= 8245798;
srom_1(10505) <= 7672112;
srom_1(10506) <= 7101785;
srom_1(10507) <= 6537492;
srom_1(10508) <= 5981880;
srom_1(10509) <= 5437554;
srom_1(10510) <= 4907067;
srom_1(10511) <= 4392905;
srom_1(10512) <= 3897481;
srom_1(10513) <= 3423117;
srom_1(10514) <= 2972039;
srom_1(10515) <= 2546360;
srom_1(10516) <= 2148078;
srom_1(10517) <= 1779059;
srom_1(10518) <= 1441035;
srom_1(10519) <= 1135591;
srom_1(10520) <= 864158;
srom_1(10521) <= 628010;
srom_1(10522) <= 428255;
srom_1(10523) <= 265828;
srom_1(10524) <= 141491;
srom_1(10525) <= 55828;
srom_1(10526) <= 9241;
srom_1(10527) <= 1947;
srom_1(10528) <= 33981;
srom_1(10529) <= 105193;
srom_1(10530) <= 215248;
srom_1(10531) <= 363632;
srom_1(10532) <= 549647;
srom_1(10533) <= 772421;
srom_1(10534) <= 1030911;
srom_1(10535) <= 1323903;
srom_1(10536) <= 1650024;
srom_1(10537) <= 2007745;
srom_1(10538) <= 2395388;
srom_1(10539) <= 2811135;
srom_1(10540) <= 3253037;
srom_1(10541) <= 3719021;
srom_1(10542) <= 4206902;
srom_1(10543) <= 4714393;
srom_1(10544) <= 5239114;
srom_1(10545) <= 5778603;
srom_1(10546) <= 6330332;
srom_1(10547) <= 6891713;
srom_1(10548) <= 7460113;
srom_1(10549) <= 8032867;
srom_1(10550) <= 8607289;
srom_1(10551) <= 9180686;
srom_1(10552) <= 9750369;
srom_1(10553) <= 10313666;
srom_1(10554) <= 10867935;
srom_1(10555) <= 11410578;
srom_1(10556) <= 11939051;
srom_1(10557) <= 12450873;
srom_1(10558) <= 12943647;
srom_1(10559) <= 13415060;
srom_1(10560) <= 13862903;
srom_1(10561) <= 14285074;
srom_1(10562) <= 14679595;
srom_1(10563) <= 15044616;
srom_1(10564) <= 15378424;
srom_1(10565) <= 15679455;
srom_1(10566) <= 15946296;
srom_1(10567) <= 16177696;
srom_1(10568) <= 16372571;
srom_1(10569) <= 16530007;
srom_1(10570) <= 16649264;
srom_1(10571) <= 16729785;
srom_1(10572) <= 16771191;
srom_1(10573) <= 16773288;
srom_1(10574) <= 16736066;
srom_1(10575) <= 16659700;
srom_1(10576) <= 16544548;
srom_1(10577) <= 16391151;
srom_1(10578) <= 16200226;
srom_1(10579) <= 15972670;
srom_1(10580) <= 15709550;
srom_1(10581) <= 15412100;
srom_1(10582) <= 15081714;
srom_1(10583) <= 14719941;
srom_1(10584) <= 14328479;
srom_1(10585) <= 13909163;
srom_1(10586) <= 13463959;
srom_1(10587) <= 12994955;
srom_1(10588) <= 12504350;
srom_1(10589) <= 11994445;
srom_1(10590) <= 11467631;
srom_1(10591) <= 10926378;
srom_1(10592) <= 10373225;
srom_1(10593) <= 9810765;
srom_1(10594) <= 9241637;
srom_1(10595) <= 8668508;
srom_1(10596) <= 8094067;
srom_1(10597) <= 7521006;
srom_1(10598) <= 6952015;
srom_1(10599) <= 6389760;
srom_1(10600) <= 5836878;
srom_1(10601) <= 5295962;
srom_1(10602) <= 4769549;
srom_1(10603) <= 4260106;
srom_1(10604) <= 3770024;
srom_1(10605) <= 3301600;
srom_1(10606) <= 2857030;
srom_1(10607) <= 2438400;
srom_1(10608) <= 2047673;
srom_1(10609) <= 1686680;
srom_1(10610) <= 1357115;
srom_1(10611) <= 1060523;
srom_1(10612) <= 798295;
srom_1(10613) <= 571660;
srom_1(10614) <= 381682;
srom_1(10615) <= 229251;
srom_1(10616) <= 115082;
srom_1(10617) <= 39711;
srom_1(10618) <= 3490;
srom_1(10619) <= 6590;
srom_1(10620) <= 48996;
srom_1(10621) <= 130510;
srom_1(10622) <= 250748;
srom_1(10623) <= 409148;
srom_1(10624) <= 604966;
srom_1(10625) <= 837284;
srom_1(10626) <= 1105014;
srom_1(10627) <= 1406898;
srom_1(10628) <= 1741522;
srom_1(10629) <= 2107316;
srom_1(10630) <= 2502566;
srom_1(10631) <= 2925417;
srom_1(10632) <= 3373887;
srom_1(10633) <= 3845873;
srom_1(10634) <= 4339161;
srom_1(10635) <= 4851438;
srom_1(10636) <= 5380303;
srom_1(10637) <= 5923274;
srom_1(10638) <= 6477806;
srom_1(10639) <= 7041299;
srom_1(10640) <= 7611109;
srom_1(10641) <= 8184566;
srom_1(10642) <= 8758979;
srom_1(10643) <= 9331656;
srom_1(10644) <= 9899910;
srom_1(10645) <= 10461077;
srom_1(10646) <= 11012526;
srom_1(10647) <= 11551670;
srom_1(10648) <= 12075982;
srom_1(10649) <= 12583002;
srom_1(10650) <= 13070353;
srom_1(10651) <= 13535750;
srom_1(10652) <= 13977010;
srom_1(10653) <= 14392064;
srom_1(10654) <= 14778966;
srom_1(10655) <= 15135902;
srom_1(10656) <= 15461197;
srom_1(10657) <= 15753326;
srom_1(10658) <= 16010919;
srom_1(10659) <= 16232769;
srom_1(10660) <= 16417835;
srom_1(10661) <= 16565249;
srom_1(10662) <= 16674320;
srom_1(10663) <= 16744536;
srom_1(10664) <= 16775569;
srom_1(10665) <= 16767272;
srom_1(10666) <= 16719685;
srom_1(10667) <= 16633030;
srom_1(10668) <= 16507715;
srom_1(10669) <= 16344326;
srom_1(10670) <= 16143630;
srom_1(10671) <= 15906568;
srom_1(10672) <= 15634252;
srom_1(10673) <= 15327959;
srom_1(10674) <= 14989125;
srom_1(10675) <= 14619338;
srom_1(10676) <= 14220333;
srom_1(10677) <= 13793982;
srom_1(10678) <= 13342283;
srom_1(10679) <= 12867354;
srom_1(10680) <= 12371423;
srom_1(10681) <= 11856815;
srom_1(10682) <= 11325943;
srom_1(10683) <= 10781298;
srom_1(10684) <= 10225432;
srom_1(10685) <= 9660953;
srom_1(10686) <= 9090507;
srom_1(10687) <= 8516770;
srom_1(10688) <= 7942431;
srom_1(10689) <= 7370185;
srom_1(10690) <= 6802715;
srom_1(10691) <= 6242682;
srom_1(10692) <= 5692711;
srom_1(10693) <= 5155382;
srom_1(10694) <= 4633216;
srom_1(10695) <= 4128659;
srom_1(10696) <= 3644079;
srom_1(10697) <= 3181748;
srom_1(10698) <= 2743833;
srom_1(10699) <= 2332389;
srom_1(10700) <= 1949344;
srom_1(10701) <= 1596495;
srom_1(10702) <= 1275497;
srom_1(10703) <= 987854;
srom_1(10704) <= 734917;
srom_1(10705) <= 517870;
srom_1(10706) <= 337731;
srom_1(10707) <= 195346;
srom_1(10708) <= 91382;
srom_1(10709) <= 26327;
srom_1(10710) <= 485;
srom_1(10711) <= 13978;
srom_1(10712) <= 66742;
srom_1(10713) <= 158530;
srom_1(10714) <= 288912;
srom_1(10715) <= 457277;
srom_1(10716) <= 662834;
srom_1(10717) <= 904620;
srom_1(10718) <= 1181501;
srom_1(10719) <= 1492178;
srom_1(10720) <= 1835195;
srom_1(10721) <= 2208944;
srom_1(10722) <= 2611671;
srom_1(10723) <= 3041488;
srom_1(10724) <= 3496379;
srom_1(10725) <= 3974212;
srom_1(10726) <= 4472745;
srom_1(10727) <= 4989642;
srom_1(10728) <= 5522477;
srom_1(10729) <= 6068752;
srom_1(10730) <= 6625906;
srom_1(10731) <= 7191326;
srom_1(10732) <= 7762361;
srom_1(10733) <= 8336332;
srom_1(10734) <= 8910548;
srom_1(10735) <= 9482316;
srom_1(10736) <= 10048956;
srom_1(10737) <= 10607810;
srom_1(10738) <= 11156257;
srom_1(10739) <= 11691726;
srom_1(10740) <= 12211706;
srom_1(10741) <= 12713757;
srom_1(10742) <= 13195527;
srom_1(10743) <= 13654755;
srom_1(10744) <= 14089288;
srom_1(10745) <= 14497089;
srom_1(10746) <= 14876245;
srom_1(10747) <= 15224978;
srom_1(10748) <= 15541654;
srom_1(10749) <= 15824786;
srom_1(10750) <= 16073047;
srom_1(10751) <= 16285273;
srom_1(10752) <= 16460470;
srom_1(10753) <= 16597814;
srom_1(10754) <= 16696663;
srom_1(10755) <= 16756552;
srom_1(10756) <= 16777201;
srom_1(10757) <= 16758513;
srom_1(10758) <= 16700576;
srom_1(10759) <= 16603661;
srom_1(10760) <= 16468223;
srom_1(10761) <= 16294897;
srom_1(10762) <= 16084495;
srom_1(10763) <= 15838005;
srom_1(10764) <= 15556582;
srom_1(10765) <= 15241546;
srom_1(10766) <= 14894374;
srom_1(10767) <= 14516695;
srom_1(10768) <= 14110278;
srom_1(10769) <= 13677031;
srom_1(10770) <= 13218985;
srom_1(10771) <= 12738287;
srom_1(10772) <= 12237192;
srom_1(10773) <= 11718050;
srom_1(10774) <= 11183294;
srom_1(10775) <= 10635434;
srom_1(10776) <= 10077037;
srom_1(10777) <= 9510723;
srom_1(10778) <= 8939147;
srom_1(10779) <= 8364989;
srom_1(10780) <= 7790942;
srom_1(10781) <= 7219698;
srom_1(10782) <= 6653934;
srom_1(10783) <= 6096306;
srom_1(10784) <= 5549427;
srom_1(10785) <= 5015861;
srom_1(10786) <= 4498112;
srom_1(10787) <= 3998607;
srom_1(10788) <= 3519687;
srom_1(10789) <= 3063600;
srom_1(10790) <= 2632484;
srom_1(10791) <= 2228360;
srom_1(10792) <= 1853123;
srom_1(10793) <= 1508534;
srom_1(10794) <= 1196207;
srom_1(10795) <= 917609;
srom_1(10796) <= 674044;
srom_1(10797) <= 466656;
srom_1(10798) <= 296416;
srom_1(10799) <= 164123;
srom_1(10800) <= 70398;
srom_1(10801) <= 15680;
srom_1(10802) <= 225;
srom_1(10803) <= 24107;
srom_1(10804) <= 87212;
srom_1(10805) <= 189245;
srom_1(10806) <= 329728;
srom_1(10807) <= 508002;
srom_1(10808) <= 723231;
srom_1(10809) <= 974405;
srom_1(10810) <= 1260347;
srom_1(10811) <= 1579716;
srom_1(10812) <= 1931014;
srom_1(10813) <= 2312594;
srom_1(10814) <= 2722667;
srom_1(10815) <= 3159309;
srom_1(10816) <= 3620473;
srom_1(10817) <= 4103997;
srom_1(10818) <= 4607612;
srom_1(10819) <= 5128958;
srom_1(10820) <= 5665589;
srom_1(10821) <= 6214990;
srom_1(10822) <= 6774583;
srom_1(10823) <= 7341745;
srom_1(10824) <= 7913817;
srom_1(10825) <= 8488114;
srom_1(10826) <= 9061945;
srom_1(10827) <= 9632619;
srom_1(10828) <= 10197459;
srom_1(10829) <= 10753816;
srom_1(10830) <= 11299083;
srom_1(10831) <= 11830701;
srom_1(10832) <= 12346178;
srom_1(10833) <= 12843096;
srom_1(10834) <= 13319126;
srom_1(10835) <= 13772035;
srom_1(10836) <= 14199700;
srom_1(10837) <= 14600114;
srom_1(10838) <= 14971400;
srom_1(10839) <= 15311817;
srom_1(10840) <= 15619769;
srom_1(10841) <= 15893811;
srom_1(10842) <= 16132659;
srom_1(10843) <= 16335193;
srom_1(10844) <= 16500462;
srom_1(10845) <= 16627692;
srom_1(10846) <= 16716286;
srom_1(10847) <= 16765828;
srom_1(10848) <= 16776087;
srom_1(10849) <= 16747015;
srom_1(10850) <= 16678746;
srom_1(10851) <= 16571603;
srom_1(10852) <= 16426086;
srom_1(10853) <= 16242879;
srom_1(10854) <= 16022841;
srom_1(10855) <= 15767003;
srom_1(10856) <= 15476565;
srom_1(10857) <= 15152890;
srom_1(10858) <= 14797494;
srom_1(10859) <= 14412045;
srom_1(10860) <= 13998350;
srom_1(10861) <= 13558349;
srom_1(10862) <= 13094105;
srom_1(10863) <= 12607796;
srom_1(10864) <= 12101701;
srom_1(10865) <= 11578194;
srom_1(10866) <= 11039730;
srom_1(10867) <= 10488835;
srom_1(10868) <= 9928090;
srom_1(10869) <= 9360126;
srom_1(10870) <= 8787607;
srom_1(10871) <= 8213216;
srom_1(10872) <= 7639648;
srom_1(10873) <= 7069592;
srom_1(10874) <= 6505722;
srom_1(10875) <= 5950681;
srom_1(10876) <= 5407072;
srom_1(10877) <= 4877444;
srom_1(10878) <= 4364282;
srom_1(10879) <= 3869991;
srom_1(10880) <= 3396890;
srom_1(10881) <= 2947196;
srom_1(10882) <= 2523019;
srom_1(10883) <= 2126348;
srom_1(10884) <= 1759042;
srom_1(10885) <= 1422825;
srom_1(10886) <= 1119273;
srom_1(10887) <= 849809;
srom_1(10888) <= 615697;
srom_1(10889) <= 418035;
srom_1(10890) <= 257750;
srom_1(10891) <= 135593;
srom_1(10892) <= 52138;
srom_1(10893) <= 7775;
srom_1(10894) <= 2712;
srom_1(10895) <= 36974;
srom_1(10896) <= 110400;
srom_1(10897) <= 222645;
srom_1(10898) <= 373183;
srom_1(10899) <= 561308;
srom_1(10900) <= 786138;
srom_1(10901) <= 1046618;
srom_1(10902) <= 1341528;
srom_1(10903) <= 1669484;
srom_1(10904) <= 2028948;
srom_1(10905) <= 2418234;
srom_1(10906) <= 2835518;
srom_1(10907) <= 3278842;
srom_1(10908) <= 3746128;
srom_1(10909) <= 4235184;
srom_1(10910) <= 4743716;
srom_1(10911) <= 5269341;
srom_1(10912) <= 5809593;
srom_1(10913) <= 6361939;
srom_1(10914) <= 6923789;
srom_1(10915) <= 7492507;
srom_1(10916) <= 8065428;
srom_1(10917) <= 8639864;
srom_1(10918) <= 9213123;
srom_1(10919) <= 9782514;
srom_1(10920) <= 10345369;
srom_1(10921) <= 10899049;
srom_1(10922) <= 11440955;
srom_1(10923) <= 11968549;
srom_1(10924) <= 12479354;
srom_1(10925) <= 12970977;
srom_1(10926) <= 13441112;
srom_1(10927) <= 13887553;
srom_1(10928) <= 14308209;
srom_1(10929) <= 14701105;
srom_1(10930) <= 15064399;
srom_1(10931) <= 15396389;
srom_1(10932) <= 15695517;
srom_1(10933) <= 15960380;
srom_1(10934) <= 16189736;
srom_1(10935) <= 16382510;
srom_1(10936) <= 16537798;
srom_1(10937) <= 16654872;
srom_1(10938) <= 16733182;
srom_1(10939) <= 16772362;
srom_1(10940) <= 16772227;
srom_1(10941) <= 16732779;
srom_1(10942) <= 16654202;
srom_1(10943) <= 16536865;
srom_1(10944) <= 16381318;
srom_1(10945) <= 16188290;
srom_1(10946) <= 15958687;
srom_1(10947) <= 15693585;
srom_1(10948) <= 15394228;
srom_1(10949) <= 15062019;
srom_1(10950) <= 14698516;
srom_1(10951) <= 14305423;
srom_1(10952) <= 13884585;
srom_1(10953) <= 13437974;
srom_1(10954) <= 12967685;
srom_1(10955) <= 12475923;
srom_1(10956) <= 11964994;
srom_1(10957) <= 11437294;
srom_1(10958) <= 10895298;
srom_1(10959) <= 10341548;
srom_1(10960) <= 9778639;
srom_1(10961) <= 9209212;
srom_1(10962) <= 8635936;
srom_1(10963) <= 8061501;
srom_1(10964) <= 7488600;
srom_1(10965) <= 6919919;
srom_1(10966) <= 6358126;
srom_1(10967) <= 5805854;
srom_1(10968) <= 5265693;
srom_1(10969) <= 4740177;
srom_1(10970) <= 4231770;
srom_1(10971) <= 3742855;
srom_1(10972) <= 3275726;
srom_1(10973) <= 2832573;
srom_1(10974) <= 2415474;
srom_1(10975) <= 2026386;
srom_1(10976) <= 1667132;
srom_1(10977) <= 1339397;
srom_1(10978) <= 1044718;
srom_1(10979) <= 784478;
srom_1(10980) <= 559895;
srom_1(10981) <= 372025;
srom_1(10982) <= 221746;
srom_1(10983) <= 109765;
srom_1(10984) <= 36607;
srom_1(10985) <= 2613;
srom_1(10986) <= 7945;
srom_1(10987) <= 52576;
srom_1(10988) <= 136298;
srom_1(10989) <= 258718;
srom_1(10990) <= 419261;
srom_1(10991) <= 617176;
srom_1(10992) <= 851534;
srom_1(10993) <= 1121235;
srom_1(10994) <= 1425016;
srom_1(10995) <= 1761451;
srom_1(10996) <= 2128963;
srom_1(10997) <= 2525829;
srom_1(10998) <= 2950188;
srom_1(10999) <= 3400049;
srom_1(11000) <= 3873303;
srom_1(11001) <= 4367731;
srom_1(11002) <= 4881014;
srom_1(11003) <= 5410746;
srom_1(11004) <= 5954441;
srom_1(11005) <= 6509552;
srom_1(11006) <= 7073474;
srom_1(11007) <= 7643563;
srom_1(11008) <= 8217146;
srom_1(11009) <= 8791532;
srom_1(11010) <= 9364030;
srom_1(11011) <= 9931953;
srom_1(11012) <= 10492639;
srom_1(11013) <= 11043459;
srom_1(11014) <= 11581829;
srom_1(11015) <= 12105224;
srom_1(11016) <= 12611192;
srom_1(11017) <= 13097358;
srom_1(11018) <= 13561443;
srom_1(11019) <= 14001271;
srom_1(11020) <= 14414780;
srom_1(11021) <= 14800029;
srom_1(11022) <= 15155213;
srom_1(11023) <= 15478667;
srom_1(11024) <= 15768872;
srom_1(11025) <= 16024469;
srom_1(11026) <= 16244259;
srom_1(11027) <= 16427211;
srom_1(11028) <= 16572467;
srom_1(11029) <= 16679346;
srom_1(11030) <= 16747347;
srom_1(11031) <= 16776151;
srom_1(11032) <= 16765623;
srom_1(11033) <= 16715812;
srom_1(11034) <= 16626952;
srom_1(11035) <= 16499460;
srom_1(11036) <= 16333933;
srom_1(11037) <= 16131148;
srom_1(11038) <= 15892055;
srom_1(11039) <= 15617776;
srom_1(11040) <= 15309597;
srom_1(11041) <= 14968963;
srom_1(11042) <= 14597472;
srom_1(11043) <= 14196865;
srom_1(11044) <= 13769021;
srom_1(11045) <= 13315946;
srom_1(11046) <= 12839766;
srom_1(11047) <= 12342712;
srom_1(11048) <= 11827117;
srom_1(11049) <= 11295397;
srom_1(11050) <= 10750046;
srom_1(11051) <= 10193621;
srom_1(11052) <= 9628732;
srom_1(11053) <= 9058028;
srom_1(11054) <= 8484185;
srom_1(11055) <= 7909893;
srom_1(11056) <= 7337846;
srom_1(11057) <= 6770727;
srom_1(11058) <= 6211194;
srom_1(11059) <= 5661872;
srom_1(11060) <= 5125337;
srom_1(11061) <= 4604104;
srom_1(11062) <= 4100618;
srom_1(11063) <= 3617240;
srom_1(11064) <= 3156237;
srom_1(11065) <= 2719770;
srom_1(11066) <= 2309886;
srom_1(11067) <= 1928507;
srom_1(11068) <= 1577422;
srom_1(11069) <= 1258276;
srom_1(11070) <= 972568;
srom_1(11071) <= 721636;
srom_1(11072) <= 506656;
srom_1(11073) <= 328638;
srom_1(11074) <= 188416;
srom_1(11075) <= 86648;
srom_1(11076) <= 23810;
srom_1(11077) <= 197;
srom_1(11078) <= 15921;
srom_1(11079) <= 70907;
srom_1(11080) <= 164898;
srom_1(11081) <= 297452;
srom_1(11082) <= 467949;
srom_1(11083) <= 675588;
srom_1(11084) <= 919397;
srom_1(11085) <= 1198231;
srom_1(11086) <= 1510783;
srom_1(11087) <= 1855588;
srom_1(11088) <= 2231028;
srom_1(11089) <= 2635343;
srom_1(11090) <= 3066637;
srom_1(11091) <= 3522888;
srom_1(11092) <= 4001956;
srom_1(11093) <= 4501594;
srom_1(11094) <= 5019460;
srom_1(11095) <= 5553125;
srom_1(11096) <= 6100087;
srom_1(11097) <= 6657780;
srom_1(11098) <= 7223589;
srom_1(11099) <= 7794862;
srom_1(11100) <= 8368919;
srom_1(11101) <= 8943068;
srom_1(11102) <= 9514618;
srom_1(11103) <= 10080887;
srom_1(11104) <= 10639220;
srom_1(11105) <= 11187000;
srom_1(11106) <= 11721656;
srom_1(11107) <= 12240683;
srom_1(11108) <= 12741647;
srom_1(11109) <= 13222197;
srom_1(11110) <= 13680081;
srom_1(11111) <= 14113152;
srom_1(11112) <= 14519378;
srom_1(11113) <= 14896855;
srom_1(11114) <= 15243812;
srom_1(11115) <= 15558623;
srom_1(11116) <= 15839811;
srom_1(11117) <= 16086058;
srom_1(11118) <= 16296209;
srom_1(11119) <= 16469279;
srom_1(11120) <= 16604456;
srom_1(11121) <= 16701105;
srom_1(11122) <= 16758775;
srom_1(11123) <= 16777194;
srom_1(11124) <= 16756276;
srom_1(11125) <= 16696119;
srom_1(11126) <= 16597005;
srom_1(11127) <= 16459399;
srom_1(11128) <= 16283947;
srom_1(11129) <= 16071470;
srom_1(11130) <= 15822966;
srom_1(11131) <= 15539600;
srom_1(11132) <= 15222700;
srom_1(11133) <= 14873753;
srom_1(11134) <= 14494395;
srom_1(11135) <= 14086404;
srom_1(11136) <= 13651695;
srom_1(11137) <= 13192305;
srom_1(11138) <= 12710389;
srom_1(11139) <= 12208207;
srom_1(11140) <= 11688113;
srom_1(11141) <= 11152547;
srom_1(11142) <= 10604020;
srom_1(11143) <= 10045104;
srom_1(11144) <= 9478420;
srom_1(11145) <= 8906625;
srom_1(11146) <= 8332402;
srom_1(11147) <= 7758442;
srom_1(11148) <= 7187437;
srom_1(11149) <= 6622064;
srom_1(11150) <= 6064976;
srom_1(11151) <= 5518784;
srom_1(11152) <= 4986049;
srom_1(11153) <= 4469270;
srom_1(11154) <= 3970871;
srom_1(11155) <= 3493187;
srom_1(11156) <= 3038460;
srom_1(11157) <= 2608822;
srom_1(11158) <= 2206287;
srom_1(11159) <= 1832743;
srom_1(11160) <= 1489942;
srom_1(11161) <= 1179490;
srom_1(11162) <= 902845;
srom_1(11163) <= 661304;
srom_1(11164) <= 455998;
srom_1(11165) <= 287891;
srom_1(11166) <= 157771;
srom_1(11167) <= 66248;
srom_1(11168) <= 13752;
srom_1(11169) <= 528;
srom_1(11170) <= 26639;
srom_1(11171) <= 91962;
srom_1(11172) <= 196190;
srom_1(11173) <= 338836;
srom_1(11174) <= 519230;
srom_1(11175) <= 736526;
srom_1(11176) <= 989705;
srom_1(11177) <= 1277581;
srom_1(11178) <= 1598802;
srom_1(11179) <= 1951863;
srom_1(11180) <= 2335109;
srom_1(11181) <= 2746741;
srom_1(11182) <= 3184829;
srom_1(11183) <= 3647321;
srom_1(11184) <= 4132045;
srom_1(11185) <= 4636730;
srom_1(11186) <= 5159009;
srom_1(11187) <= 5696433;
srom_1(11188) <= 6246481;
srom_1(11189) <= 6806574;
srom_1(11190) <= 7374086;
srom_1(11191) <= 7946356;
srom_1(11192) <= 8520699;
srom_1(11193) <= 9094423;
srom_1(11194) <= 9664837;
srom_1(11195) <= 10229266;
srom_1(11196) <= 10785064;
srom_1(11197) <= 11329624;
srom_1(11198) <= 11860393;
srom_1(11199) <= 12374881;
srom_1(11200) <= 12870676;
srom_1(11201) <= 13345454;
srom_1(11202) <= 13796987;
srom_1(11203) <= 14223158;
srom_1(11204) <= 14621969;
srom_1(11205) <= 14991549;
srom_1(11206) <= 15330166;
srom_1(11207) <= 15636232;
srom_1(11208) <= 15908311;
srom_1(11209) <= 16145128;
srom_1(11210) <= 16345571;
srom_1(11211) <= 16508702;
srom_1(11212) <= 16633755;
srom_1(11213) <= 16720143;
srom_1(11214) <= 16767462;
srom_1(11215) <= 16775490;
srom_1(11216) <= 16744189;
srom_1(11217) <= 16673705;
srom_1(11218) <= 16564370;
srom_1(11219) <= 16416696;
srom_1(11220) <= 16231375;
srom_1(11221) <= 16009277;
srom_1(11222) <= 15751443;
srom_1(11223) <= 15459083;
srom_1(11224) <= 15133566;
srom_1(11225) <= 14776420;
srom_1(11226) <= 14389319;
srom_1(11227) <= 13974079;
srom_1(11228) <= 13532646;
srom_1(11229) <= 13067092;
srom_1(11230) <= 12579598;
srom_1(11231) <= 12072451;
srom_1(11232) <= 11548030;
srom_1(11233) <= 11008793;
srom_1(11234) <= 10457269;
srom_1(11235) <= 9896044;
srom_1(11236) <= 9327751;
srom_1(11237) <= 8755053;
srom_1(11238) <= 8180637;
srom_1(11239) <= 7607196;
srom_1(11240) <= 7037420;
srom_1(11241) <= 6473980;
srom_1(11242) <= 5919518;
srom_1(11243) <= 5376634;
srom_1(11244) <= 4847875;
srom_1(11245) <= 4335720;
srom_1(11246) <= 3842569;
srom_1(11247) <= 3370737;
srom_1(11248) <= 2922435;
srom_1(11249) <= 2499766;
srom_1(11250) <= 2104712;
srom_1(11251) <= 1739125;
srom_1(11252) <= 1404720;
srom_1(11253) <= 1103065;
srom_1(11254) <= 835574;
srom_1(11255) <= 603502;
srom_1(11256) <= 407937;
srom_1(11257) <= 249795;
srom_1(11258) <= 129820;
srom_1(11259) <= 48573;
srom_1(11260) <= 6435;
srom_1(11261) <= 3604;
srom_1(11262) <= 40094;
srom_1(11263) <= 115732;
srom_1(11264) <= 230165;
srom_1(11265) <= 382855;
srom_1(11266) <= 573087;
srom_1(11267) <= 799969;
srom_1(11268) <= 1062436;
srom_1(11269) <= 1359259;
srom_1(11270) <= 1689044;
srom_1(11271) <= 2050246;
srom_1(11272) <= 2441171;
srom_1(11273) <= 2859985;
srom_1(11274) <= 3304725;
srom_1(11275) <= 3773305;
srom_1(11276) <= 4263528;
srom_1(11277) <= 4773095;
srom_1(11278) <= 5299616;
srom_1(11279) <= 5840622;
srom_1(11280) <= 6393577;
srom_1(11281) <= 6955887;
srom_1(11282) <= 7524915;
srom_1(11283) <= 8097994;
srom_1(11284) <= 8672436;
srom_1(11285) <= 9245546;
srom_1(11286) <= 9814638;
srom_1(11287) <= 10377043;
srom_1(11288) <= 10930124;
srom_1(11289) <= 11471286;
srom_1(11290) <= 11997993;
srom_1(11291) <= 12507774;
srom_1(11292) <= 12998239;
srom_1(11293) <= 13467087;
srom_1(11294) <= 13912121;
srom_1(11295) <= 14331254;
srom_1(11296) <= 14722519;
srom_1(11297) <= 15084082;
srom_1(11298) <= 15414248;
srom_1(11299) <= 15711468;
srom_1(11300) <= 15974349;
srom_1(11301) <= 16201658;
srom_1(11302) <= 16392328;
srom_1(11303) <= 16545467;
srom_1(11304) <= 16660355;
srom_1(11305) <= 16736454;
srom_1(11306) <= 16773407;
srom_1(11307) <= 16771041;
srom_1(11308) <= 16729366;
srom_1(11309) <= 16648580;
srom_1(11310) <= 16529059;
srom_1(11311) <= 16371365;
srom_1(11312) <= 16176237;
srom_1(11313) <= 15944590;
srom_1(11314) <= 15677510;
srom_1(11315) <= 15376250;
srom_1(11316) <= 15042223;
srom_1(11317) <= 14676995;
srom_1(11318) <= 14282278;
srom_1(11319) <= 13859924;
srom_1(11320) <= 13411913;
srom_1(11321) <= 12940346;
srom_1(11322) <= 12447434;
srom_1(11323) <= 11935489;
srom_1(11324) <= 11406912;
srom_1(11325) <= 10864181;
srom_1(11326) <= 10309840;
srom_1(11327) <= 9746491;
srom_1(11328) <= 9176774;
srom_1(11329) <= 8603361;
srom_1(11330) <= 8028941;
srom_1(11331) <= 7456207;
srom_1(11332) <= 6887846;
srom_1(11333) <= 6326522;
srom_1(11334) <= 5774869;
srom_1(11335) <= 5235471;
srom_1(11336) <= 4710860;
srom_1(11337) <= 4203496;
srom_1(11338) <= 3715756;
srom_1(11339) <= 3249930;
srom_1(11340) <= 2808200;
srom_1(11341) <= 2392639;
srom_1(11342) <= 2005195;
srom_1(11343) <= 1647685;
srom_1(11344) <= 1321785;
srom_1(11345) <= 1029024;
srom_1(11346) <= 770775;
srom_1(11347) <= 548248;
srom_1(11348) <= 362488;
srom_1(11349) <= 214365;
srom_1(11350) <= 104573;
srom_1(11351) <= 33629;
srom_1(11352) <= 1863;
srom_1(11353) <= 9426;
srom_1(11354) <= 56282;
srom_1(11355) <= 142211;
srom_1(11356) <= 266810;
srom_1(11357) <= 429495;
srom_1(11358) <= 629503;
srom_1(11359) <= 865896;
srom_1(11360) <= 1137566;
srom_1(11361) <= 1443238;
srom_1(11362) <= 1781480;
srom_1(11363) <= 2150704;
srom_1(11364) <= 2549181;
srom_1(11365) <= 2975040;
srom_1(11366) <= 3426286;
srom_1(11367) <= 3900801;
srom_1(11368) <= 4396361;
srom_1(11369) <= 4910643;
srom_1(11370) <= 5441233;
srom_1(11371) <= 5985645;
srom_1(11372) <= 6541326;
srom_1(11373) <= 7105668;
srom_1(11374) <= 7676027;
srom_1(11375) <= 8249728;
srom_1(11376) <= 8824080;
srom_1(11377) <= 9396389;
srom_1(11378) <= 9963973;
srom_1(11379) <= 10524169;
srom_1(11380) <= 11074351;
srom_1(11381) <= 11611939;
srom_1(11382) <= 12134411;
srom_1(11383) <= 12639318;
srom_1(11384) <= 13124292;
srom_1(11385) <= 13587059;
srom_1(11386) <= 14025448;
srom_1(11387) <= 14437404;
srom_1(11388) <= 14820995;
srom_1(11389) <= 15174423;
srom_1(11390) <= 15496030;
srom_1(11391) <= 15784307;
srom_1(11392) <= 16037903;
srom_1(11393) <= 16255630;
srom_1(11394) <= 16436465;
srom_1(11395) <= 16579561;
srom_1(11396) <= 16684247;
srom_1(11397) <= 16750031;
srom_1(11398) <= 16776606;
srom_1(11399) <= 16763847;
srom_1(11400) <= 16711814;
srom_1(11401) <= 16620750;
srom_1(11402) <= 16491082;
srom_1(11403) <= 16323420;
srom_1(11404) <= 16118548;
srom_1(11405) <= 15877428;
srom_1(11406) <= 15601190;
srom_1(11407) <= 15291131;
srom_1(11408) <= 14948702;
srom_1(11409) <= 14575512;
srom_1(11410) <= 14173308;
srom_1(11411) <= 13743979;
srom_1(11412) <= 13289536;
srom_1(11413) <= 12812111;
srom_1(11414) <= 12313942;
srom_1(11415) <= 11797366;
srom_1(11416) <= 11264806;
srom_1(11417) <= 10718758;
srom_1(11418) <= 10161783;
srom_1(11419) <= 9596493;
srom_1(11420) <= 9025539;
srom_1(11421) <= 8451598;
srom_1(11422) <= 7877362;
srom_1(11423) <= 7305523;
srom_1(11424) <= 6738763;
srom_1(11425) <= 6179740;
srom_1(11426) <= 5631075;
srom_1(11427) <= 5095341;
srom_1(11428) <= 4575050;
srom_1(11429) <= 4072642;
srom_1(11430) <= 3590473;
srom_1(11431) <= 3130805;
srom_1(11432) <= 2695792;
srom_1(11433) <= 2287474;
srom_1(11434) <= 1907767;
srom_1(11435) <= 1558451;
srom_1(11436) <= 1241164;
srom_1(11437) <= 957393;
srom_1(11438) <= 708470;
srom_1(11439) <= 495562;
srom_1(11440) <= 319667;
srom_1(11441) <= 181610;
srom_1(11442) <= 82039;
srom_1(11443) <= 21419;
srom_1(11444) <= 37;
srom_1(11445) <= 17991;
srom_1(11446) <= 75198;
srom_1(11447) <= 171390;
srom_1(11448) <= 306115;
srom_1(11449) <= 478741;
srom_1(11450) <= 688459;
srom_1(11451) <= 934286;
srom_1(11452) <= 1215069;
srom_1(11453) <= 1529492;
srom_1(11454) <= 1876078;
srom_1(11455) <= 2253205;
srom_1(11456) <= 2659102;
srom_1(11457) <= 3091867;
srom_1(11458) <= 3549470;
srom_1(11459) <= 4029766;
srom_1(11460) <= 4530502;
srom_1(11461) <= 5049329;
srom_1(11462) <= 5583816;
srom_1(11463) <= 6131455;
srom_1(11464) <= 6689679;
srom_1(11465) <= 7255870;
srom_1(11466) <= 7827373;
srom_1(11467) <= 8401507;
srom_1(11468) <= 8975581;
srom_1(11469) <= 9546902;
srom_1(11470) <= 10112792;
srom_1(11471) <= 10670596;
srom_1(11472) <= 11217699;
srom_1(11473) <= 11751536;
srom_1(11474) <= 12269603;
srom_1(11475) <= 12769471;
srom_1(11476) <= 13248795;
srom_1(11477) <= 13705328;
srom_1(11478) <= 14136929;
srom_1(11479) <= 14541574;
srom_1(11480) <= 14917366;
srom_1(11481) <= 15262542;
srom_1(11482) <= 15575484;
srom_1(11483) <= 15854724;
srom_1(11484) <= 16098954;
srom_1(11485) <= 16307026;
srom_1(11486) <= 16477967;
srom_1(11487) <= 16610973;
srom_1(11488) <= 16705422;
srom_1(11489) <= 16760871;
srom_1(11490) <= 16777059;
srom_1(11491) <= 16753911;
srom_1(11492) <= 16691536;
srom_1(11493) <= 16590224;
srom_1(11494) <= 16450453;
srom_1(11495) <= 16272877;
srom_1(11496) <= 16058329;
srom_1(11497) <= 15807815;
srom_1(11498) <= 15522510;
srom_1(11499) <= 15203751;
srom_1(11500) <= 14853034;
srom_1(11501) <= 14472003;
srom_1(11502) <= 14062444;
srom_1(11503) <= 13626280;
srom_1(11504) <= 13165553;
srom_1(11505) <= 12682427;
srom_1(11506) <= 12179165;
srom_1(11507) <= 11658127;
srom_1(11508) <= 11121758;
srom_1(11509) <= 10572572;
srom_1(11510) <= 10013145;
srom_1(11511) <= 9446100;
srom_1(11512) <= 8874096;
srom_1(11513) <= 8299815;
srom_1(11514) <= 7725951;
srom_1(11515) <= 7155194;
srom_1(11516) <= 6590221;
srom_1(11517) <= 6033681;
srom_1(11518) <= 5488184;
srom_1(11519) <= 4956288;
srom_1(11520) <= 4440488;
srom_1(11521) <= 3943201;
srom_1(11522) <= 3466761;
srom_1(11523) <= 3013401;
srom_1(11524) <= 2585247;
srom_1(11525) <= 2184307;
srom_1(11526) <= 1812461;
srom_1(11527) <= 1471453;
srom_1(11528) <= 1162882;
srom_1(11529) <= 888195;
srom_1(11530) <= 648680;
srom_1(11531) <= 445460;
srom_1(11532) <= 279488;
srom_1(11533) <= 151542;
srom_1(11534) <= 62223;
srom_1(11535) <= 11950;
srom_1(11536) <= 957;
srom_1(11537) <= 29297;
srom_1(11538) <= 96836;
srom_1(11539) <= 203259;
srom_1(11540) <= 348065;
srom_1(11541) <= 530576;
srom_1(11542) <= 749937;
srom_1(11543) <= 1005117;
srom_1(11544) <= 1294921;
srom_1(11545) <= 1617990;
srom_1(11546) <= 1972809;
srom_1(11547) <= 2357714;
srom_1(11548) <= 2770899;
srom_1(11549) <= 3210428;
srom_1(11550) <= 3674240;
srom_1(11551) <= 4160158;
srom_1(11552) <= 4665905;
srom_1(11553) <= 5189109;
srom_1(11554) <= 5727317;
srom_1(11555) <= 6278004;
srom_1(11556) <= 6838589;
srom_1(11557) <= 7406442;
srom_1(11558) <= 7978901;
srom_1(11559) <= 8553282;
srom_1(11560) <= 9126890;
srom_1(11561) <= 9697036;
srom_1(11562) <= 10261046;
srom_1(11563) <= 10816276;
srom_1(11564) <= 11360121;
srom_1(11565) <= 11890033;
srom_1(11566) <= 12403524;
srom_1(11567) <= 12898189;
srom_1(11568) <= 13371706;
srom_1(11569) <= 13821856;
srom_1(11570) <= 14246528;
srom_1(11571) <= 14643730;
srom_1(11572) <= 15011599;
srom_1(11573) <= 15348411;
srom_1(11574) <= 15652586;
srom_1(11575) <= 15922698;
srom_1(11576) <= 16157479;
srom_1(11577) <= 16355830;
srom_1(11578) <= 16516820;
srom_1(11579) <= 16639694;
srom_1(11580) <= 16723875;
srom_1(11581) <= 16768970;
srom_1(11582) <= 16774766;
srom_1(11583) <= 16741237;
srom_1(11584) <= 16668539;
srom_1(11585) <= 16557014;
srom_1(11586) <= 16407185;
srom_1(11587) <= 16219753;
srom_1(11588) <= 15995599;
srom_1(11589) <= 15735773;
srom_1(11590) <= 15441493;
srom_1(11591) <= 15114140;
srom_1(11592) <= 14755249;
srom_1(11593) <= 14366502;
srom_1(11594) <= 13949723;
srom_1(11595) <= 13506866;
srom_1(11596) <= 13040007;
srom_1(11597) <= 12551337;
srom_1(11598) <= 12043146;
srom_1(11599) <= 11517818;
srom_1(11600) <= 10977816;
srom_1(11601) <= 10425672;
srom_1(11602) <= 9863976;
srom_1(11603) <= 9295361;
srom_1(11604) <= 8722494;
srom_1(11605) <= 8148061;
srom_1(11606) <= 7574756;
srom_1(11607) <= 7005268;
srom_1(11608) <= 6442267;
srom_1(11609) <= 5888392;
srom_1(11610) <= 5346243;
srom_1(11611) <= 4818359;
srom_1(11612) <= 4307218;
srom_1(11613) <= 3815216;
srom_1(11614) <= 3344660;
srom_1(11615) <= 2897757;
srom_1(11616) <= 2476603;
srom_1(11617) <= 2083172;
srom_1(11618) <= 1719309;
srom_1(11619) <= 1386720;
srom_1(11620) <= 1086967;
srom_1(11621) <= 821453;
srom_1(11622) <= 591423;
srom_1(11623) <= 397958;
srom_1(11624) <= 241964;
srom_1(11625) <= 124172;
srom_1(11626) <= 45134;
srom_1(11627) <= 5222;
srom_1(11628) <= 4623;
srom_1(11629) <= 43339;
srom_1(11630) <= 121189;
srom_1(11631) <= 237808;
srom_1(11632) <= 392648;
srom_1(11633) <= 584984;
srom_1(11634) <= 813915;
srom_1(11635) <= 1078365;
srom_1(11636) <= 1377096;
srom_1(11637) <= 1708706;
srom_1(11638) <= 2071641;
srom_1(11639) <= 2464197;
srom_1(11640) <= 2884536;
srom_1(11641) <= 3330685;
srom_1(11642) <= 3800552;
srom_1(11643) <= 4291935;
srom_1(11644) <= 4802527;
srom_1(11645) <= 5329937;
srom_1(11646) <= 5871689;
srom_1(11647) <= 6425244;
srom_1(11648) <= 6988007;
srom_1(11649) <= 7557337;
srom_1(11650) <= 8130565;
srom_1(11651) <= 8705003;
srom_1(11652) <= 9277957;
srom_1(11653) <= 9846741;
srom_1(11654) <= 10408687;
srom_1(11655) <= 10961161;
srom_1(11656) <= 11501571;
srom_1(11657) <= 12027383;
srom_1(11658) <= 12536131;
srom_1(11659) <= 13025431;
srom_1(11660) <= 13492986;
srom_1(11661) <= 13936606;
srom_1(11662) <= 14354209;
srom_1(11663) <= 14743837;
srom_1(11664) <= 15103664;
srom_1(11665) <= 15432001;
srom_1(11666) <= 15727309;
srom_1(11667) <= 15988204;
srom_1(11668) <= 16213462;
srom_1(11669) <= 16402026;
srom_1(11670) <= 16553012;
srom_1(11671) <= 16665713;
srom_1(11672) <= 16739599;
srom_1(11673) <= 16774325;
srom_1(11674) <= 16769728;
srom_1(11675) <= 16725828;
srom_1(11676) <= 16642832;
srom_1(11677) <= 16521130;
srom_1(11678) <= 16361291;
srom_1(11679) <= 16164065;
srom_1(11680) <= 15930378;
srom_1(11681) <= 15661325;
srom_1(11682) <= 15358167;
srom_1(11683) <= 15022327;
srom_1(11684) <= 14655379;
srom_1(11685) <= 14259044;
srom_1(11686) <= 13835181;
srom_1(11687) <= 13385776;
srom_1(11688) <= 12912939;
srom_1(11689) <= 12418885;
srom_1(11690) <= 11905931;
srom_1(11691) <= 11376484;
srom_1(11692) <= 10833026;
srom_1(11693) <= 10278104;
srom_1(11694) <= 9714323;
srom_1(11695) <= 9144324;
srom_1(11696) <= 8570782;
srom_1(11697) <= 7996386;
srom_1(11698) <= 7423828;
srom_1(11699) <= 6855795;
srom_1(11700) <= 6294950;
srom_1(11701) <= 5743923;
srom_1(11702) <= 5205297;
srom_1(11703) <= 4681599;
srom_1(11704) <= 4175285;
srom_1(11705) <= 3688728;
srom_1(11706) <= 3224211;
srom_1(11707) <= 2783911;
srom_1(11708) <= 2369894;
srom_1(11709) <= 1984100;
srom_1(11710) <= 1628339;
srom_1(11711) <= 1304280;
srom_1(11712) <= 1013441;
srom_1(11713) <= 757187;
srom_1(11714) <= 536720;
srom_1(11715) <= 353072;
srom_1(11716) <= 207106;
srom_1(11717) <= 99506;
srom_1(11718) <= 30777;
srom_1(11719) <= 1240;
srom_1(11720) <= 11034;
srom_1(11721) <= 60113;
srom_1(11722) <= 148248;
srom_1(11723) <= 275025;
srom_1(11724) <= 439849;
srom_1(11725) <= 641947;
srom_1(11726) <= 880373;
srom_1(11727) <= 1154006;
srom_1(11728) <= 1461566;
srom_1(11729) <= 1801609;
srom_1(11730) <= 2172540;
srom_1(11731) <= 2572621;
srom_1(11732) <= 2999974;
srom_1(11733) <= 3452597;
srom_1(11734) <= 3928367;
srom_1(11735) <= 4425052;
srom_1(11736) <= 4940324;
srom_1(11737) <= 5471766;
srom_1(11738) <= 6016886;
srom_1(11739) <= 6573127;
srom_1(11740) <= 7137882;
srom_1(11741) <= 7708503;
srom_1(11742) <= 8282312;
srom_1(11743) <= 8856620;
srom_1(11744) <= 9428733;
srom_1(11745) <= 9995969;
srom_1(11746) <= 10555667;
srom_1(11747) <= 11105203;
srom_1(11748) <= 11642000;
srom_1(11749) <= 12163541;
srom_1(11750) <= 12667380;
srom_1(11751) <= 13151154;
srom_1(11752) <= 13612595;
srom_1(11753) <= 14049539;
srom_1(11754) <= 14459937;
srom_1(11755) <= 14841864;
srom_1(11756) <= 15193530;
srom_1(11757) <= 15513285;
srom_1(11758) <= 15799630;
srom_1(11759) <= 16051223;
srom_1(11760) <= 16266882;
srom_1(11761) <= 16445598;
srom_1(11762) <= 16586531;
srom_1(11763) <= 16689022;
srom_1(11764) <= 16752589;
srom_1(11765) <= 16776935;
srom_1(11766) <= 16761945;
srom_1(11767) <= 16707689;
srom_1(11768) <= 16614423;
srom_1(11769) <= 16482583;
srom_1(11770) <= 16312787;
srom_1(11771) <= 16105832;
srom_1(11772) <= 15862688;
srom_1(11773) <= 15584496;
srom_1(11774) <= 15272560;
srom_1(11775) <= 14928343;
srom_1(11776) <= 14553458;
srom_1(11777) <= 14149665;
srom_1(11778) <= 13718855;
srom_1(11779) <= 13263051;
srom_1(11780) <= 12784388;
srom_1(11781) <= 12285113;
srom_1(11782) <= 11767565;
srom_1(11783) <= 11234172;
srom_1(11784) <= 10687435;
srom_1(11785) <= 10129918;
srom_1(11786) <= 9564236;
srom_1(11787) <= 8993041;
srom_1(11788) <= 8419011;
srom_1(11789) <= 7844839;
srom_1(11790) <= 7273216;
srom_1(11791) <= 6706824;
srom_1(11792) <= 6148319;
srom_1(11793) <= 5600319;
srom_1(11794) <= 5065394;
srom_1(11795) <= 4546053;
srom_1(11796) <= 4044731;
srom_1(11797) <= 3563779;
srom_1(11798) <= 3105452;
srom_1(11799) <= 2671900;
srom_1(11800) <= 2265155;
srom_1(11801) <= 1887125;
srom_1(11802) <= 1539583;
srom_1(11803) <= 1224159;
srom_1(11804) <= 942331;
srom_1(11805) <= 695421;
srom_1(11806) <= 484587;
srom_1(11807) <= 310818;
srom_1(11808) <= 174928;
srom_1(11809) <= 77555;
srom_1(11810) <= 19155;
srom_1(11811) <= 3;
srom_1(11812) <= 20188;
srom_1(11813) <= 79615;
srom_1(11814) <= 178005;
srom_1(11815) <= 314899;
srom_1(11816) <= 489652;
srom_1(11817) <= 701446;
srom_1(11818) <= 949289;
srom_1(11819) <= 1232016;
srom_1(11820) <= 1548304;
srom_1(11821) <= 1896668;
srom_1(11822) <= 2275474;
srom_1(11823) <= 2682948;
srom_1(11824) <= 3117177;
srom_1(11825) <= 3576126;
srom_1(11826) <= 4057642;
srom_1(11827) <= 4559467;
srom_1(11828) <= 5079249;
srom_1(11829) <= 5614549;
srom_1(11830) <= 6162858;
srom_1(11831) <= 6721605;
srom_1(11832) <= 7288168;
srom_1(11833) <= 7859892;
srom_1(11834) <= 8434094;
srom_1(11835) <= 9008084;
srom_1(11836) <= 9579169;
srom_1(11837) <= 10144671;
srom_1(11838) <= 10701938;
srom_1(11839) <= 11248357;
srom_1(11840) <= 11781365;
srom_1(11841) <= 12298464;
srom_1(11842) <= 12797228;
srom_1(11843) <= 13275319;
srom_1(11844) <= 13730494;
srom_1(11845) <= 14160619;
srom_1(11846) <= 14563677;
srom_1(11847) <= 14937779;
srom_1(11848) <= 15281169;
srom_1(11849) <= 15592237;
srom_1(11850) <= 15869525;
srom_1(11851) <= 16111732;
srom_1(11852) <= 16317723;
srom_1(11853) <= 16486532;
srom_1(11854) <= 16617367;
srom_1(11855) <= 16709614;
srom_1(11856) <= 16762841;
srom_1(11857) <= 16776799;
srom_1(11858) <= 16751421;
srom_1(11859) <= 16686827;
srom_1(11860) <= 16583320;
srom_1(11861) <= 16441386;
srom_1(11862) <= 16261689;
srom_1(11863) <= 16045072;
srom_1(11864) <= 15792552;
srom_1(11865) <= 15505312;
srom_1(11866) <= 15184699;
srom_1(11867) <= 14832217;
srom_1(11868) <= 14449519;
srom_1(11869) <= 14038399;
srom_1(11870) <= 13600785;
srom_1(11871) <= 13138730;
srom_1(11872) <= 12654399;
srom_1(11873) <= 12150065;
srom_1(11874) <= 11628092;
srom_1(11875) <= 11090928;
srom_1(11876) <= 10541092;
srom_1(11877) <= 9981162;
srom_1(11878) <= 9413764;
srom_1(11879) <= 8841559;
srom_1(11880) <= 8267230;
srom_1(11881) <= 7693470;
srom_1(11882) <= 7122969;
srom_1(11883) <= 6558404;
srom_1(11884) <= 6002421;
srom_1(11885) <= 5457628;
srom_1(11886) <= 4926579;
srom_1(11887) <= 4411765;
srom_1(11888) <= 3915599;
srom_1(11889) <= 3440409;
srom_1(11890) <= 2988423;
srom_1(11891) <= 2561760;
srom_1(11892) <= 2162421;
srom_1(11893) <= 1792279;
srom_1(11894) <= 1453070;
srom_1(11895) <= 1146383;
srom_1(11896) <= 873658;
srom_1(11897) <= 636173;
srom_1(11898) <= 435042;
srom_1(11899) <= 271207;
srom_1(11900) <= 145438;
srom_1(11901) <= 58324;
srom_1(11902) <= 10274;
srom_1(11903) <= 1513;
srom_1(11904) <= 32081;
srom_1(11905) <= 101836;
srom_1(11906) <= 210451;
srom_1(11907) <= 357415;
srom_1(11908) <= 542041;
srom_1(11909) <= 763462;
srom_1(11910) <= 1020640;
srom_1(11911) <= 1312369;
srom_1(11912) <= 1637281;
srom_1(11913) <= 1993852;
srom_1(11914) <= 2380410;
srom_1(11915) <= 2795143;
srom_1(11916) <= 3236106;
srom_1(11917) <= 3701230;
srom_1(11918) <= 4188335;
srom_1(11919) <= 4695136;
srom_1(11920) <= 5219258;
srom_1(11921) <= 5758241;
srom_1(11922) <= 6309560;
srom_1(11923) <= 6870627;
srom_1(11924) <= 7438814;
srom_1(11925) <= 8011453;
srom_1(11926) <= 8585862;
srom_1(11927) <= 9159345;
srom_1(11928) <= 9729215;
srom_1(11929) <= 10292797;
srom_1(11930) <= 10847451;
srom_1(11931) <= 11390574;
srom_1(11932) <= 11919619;
srom_1(11933) <= 12432107;
srom_1(11934) <= 12925633;
srom_1(11935) <= 13397884;
srom_1(11936) <= 13846644;
srom_1(11937) <= 14269809;
srom_1(11938) <= 14665396;
srom_1(11939) <= 15031549;
srom_1(11940) <= 15366550;
srom_1(11941) <= 15668830;
srom_1(11942) <= 15936970;
srom_1(11943) <= 16169714;
srom_1(11944) <= 16365969;
srom_1(11945) <= 16524815;
srom_1(11946) <= 16645508;
srom_1(11947) <= 16727481;
srom_1(11948) <= 16770351;
srom_1(11949) <= 16773916;
srom_1(11950) <= 16738159;
srom_1(11951) <= 16663248;
srom_1(11952) <= 16549535;
srom_1(11953) <= 16397552;
srom_1(11954) <= 16208013;
srom_1(11955) <= 15981805;
srom_1(11956) <= 15719991;
srom_1(11957) <= 15423797;
srom_1(11958) <= 15094613;
srom_1(11959) <= 14733982;
srom_1(11960) <= 14343595;
srom_1(11961) <= 13925283;
srom_1(11962) <= 13481008;
srom_1(11963) <= 13012853;
srom_1(11964) <= 12523013;
srom_1(11965) <= 12013786;
srom_1(11966) <= 11487559;
srom_1(11967) <= 10946800;
srom_1(11968) <= 10394044;
srom_1(11969) <= 9831885;
srom_1(11970) <= 9262957;
srom_1(11971) <= 8689929;
srom_1(11972) <= 8115488;
srom_1(11973) <= 7542328;
srom_1(11974) <= 6973137;
srom_1(11975) <= 6410583;
srom_1(11976) <= 5857305;
srom_1(11977) <= 5315896;
srom_1(11978) <= 4788897;
srom_1(11979) <= 4278778;
srom_1(11980) <= 3787932;
srom_1(11981) <= 3318660;
srom_1(11982) <= 2873162;
srom_1(11983) <= 2453528;
srom_1(11984) <= 2061726;
srom_1(11985) <= 1699593;
srom_1(11986) <= 1368827;
srom_1(11987) <= 1070979;
srom_1(11988) <= 807445;
srom_1(11989) <= 579463;
srom_1(11990) <= 388100;
srom_1(11991) <= 234255;
srom_1(11992) <= 118648;
srom_1(11993) <= 41821;
srom_1(11994) <= 4136;
srom_1(11995) <= 5768;
srom_1(11996) <= 46710;
srom_1(11997) <= 126771;
srom_1(11998) <= 245573;
srom_1(11999) <= 402562;
srom_1(12000) <= 596999;
srom_1(12001) <= 827975;
srom_1(12002) <= 1094404;
srom_1(12003) <= 1395039;
srom_1(12004) <= 1728469;
srom_1(12005) <= 2093130;
srom_1(12006) <= 2487313;
srom_1(12007) <= 2909170;
srom_1(12008) <= 3356721;
srom_1(12009) <= 3827868;
srom_1(12010) <= 4320403;
srom_1(12011) <= 4832014;
srom_1(12012) <= 5360304;
srom_1(12013) <= 5902795;
srom_1(12014) <= 6456942;
srom_1(12015) <= 7020147;
srom_1(12016) <= 7589770;
srom_1(12017) <= 8163139;
srom_1(12018) <= 8737565;
srom_1(12019) <= 9310354;
srom_1(12020) <= 9878822;
srom_1(12021) <= 10440301;
srom_1(12022) <= 10992159;
srom_1(12023) <= 11531808;
srom_1(12024) <= 12056717;
srom_1(12025) <= 12564426;
srom_1(12026) <= 13052552;
srom_1(12027) <= 13518808;
srom_1(12028) <= 13961007;
srom_1(12029) <= 14377074;
srom_1(12030) <= 14765060;
srom_1(12031) <= 15123144;
srom_1(12032) <= 15449648;
srom_1(12033) <= 15743040;
srom_1(12034) <= 16001944;
srom_1(12035) <= 16225147;
srom_1(12036) <= 16411602;
srom_1(12037) <= 16560434;
srom_1(12038) <= 16670946;
srom_1(12039) <= 16742619;
srom_1(12040) <= 16775117;
srom_1(12041) <= 16768288;
srom_1(12042) <= 16722164;
srom_1(12043) <= 16636960;
srom_1(12044) <= 16513078;
srom_1(12045) <= 16351097;
srom_1(12046) <= 16151777;
srom_1(12047) <= 15916053;
srom_1(12048) <= 15645030;
srom_1(12049) <= 15339979;
srom_1(12050) <= 15002331;
srom_1(12051) <= 14633669;
srom_1(12052) <= 14235722;
srom_1(12053) <= 13810355;
srom_1(12054) <= 13359564;
srom_1(12055) <= 12885463;
srom_1(12056) <= 12390274;
srom_1(12057) <= 11876320;
srom_1(12058) <= 11346011;
srom_1(12059) <= 10801834;
srom_1(12060) <= 10246340;
srom_1(12061) <= 9682135;
srom_1(12062) <= 9111863;
srom_1(12063) <= 8538201;
srom_1(12064) <= 7963836;
srom_1(12065) <= 7391464;
srom_1(12066) <= 6823768;
srom_1(12067) <= 6263409;
srom_1(12068) <= 5713017;
srom_1(12069) <= 5175171;
srom_1(12070) <= 4652394;
srom_1(12071) <= 4147138;
srom_1(12072) <= 3661771;
srom_1(12073) <= 3198570;
srom_1(12074) <= 2759707;
srom_1(12075) <= 2347239;
srom_1(12076) <= 1963102;
srom_1(12077) <= 1609096;
srom_1(12078) <= 1286882;
srom_1(12079) <= 997970;
srom_1(12080) <= 743715;
srom_1(12081) <= 525310;
srom_1(12082) <= 343778;
srom_1(12083) <= 199972;
srom_1(12084) <= 94564;
srom_1(12085) <= 28051;
srom_1(12086) <= 743;
srom_1(12087) <= 12768;
srom_1(12088) <= 64071;
srom_1(12089) <= 154410;
srom_1(12090) <= 283362;
srom_1(12091) <= 450323;
srom_1(12092) <= 654508;
srom_1(12093) <= 894962;
srom_1(12094) <= 1170556;
srom_1(12095) <= 1479998;
srom_1(12096) <= 1821837;
srom_1(12097) <= 2194469;
srom_1(12098) <= 2596148;
srom_1(12099) <= 3024990;
srom_1(12100) <= 3478984;
srom_1(12101) <= 3956000;
srom_1(12102) <= 4453803;
srom_1(12103) <= 4970057;
srom_1(12104) <= 5502342;
srom_1(12105) <= 6048162;
srom_1(12106) <= 6604956;
srom_1(12107) <= 7170115;
srom_1(12108) <= 7740988;
srom_1(12109) <= 8314898;
srom_1(12110) <= 8889153;
srom_1(12111) <= 9461062;
srom_1(12112) <= 10027941;
srom_1(12113) <= 10587132;
srom_1(12114) <= 11136014;
srom_1(12115) <= 11672013;
srom_1(12116) <= 12192614;
srom_1(12117) <= 12695378;
srom_1(12118) <= 13177945;
srom_1(12119) <= 13638053;
srom_1(12120) <= 14073545;
srom_1(12121) <= 14482379;
srom_1(12122) <= 14862636;
srom_1(12123) <= 15212535;
srom_1(12124) <= 15530433;
srom_1(12125) <= 15814842;
srom_1(12126) <= 16064426;
srom_1(12127) <= 16278016;
srom_1(12128) <= 16454609;
srom_1(12129) <= 16593378;
srom_1(12130) <= 16693672;
srom_1(12131) <= 16755021;
srom_1(12132) <= 16777137;
srom_1(12133) <= 16759916;
srom_1(12134) <= 16703440;
srom_1(12135) <= 16607972;
srom_1(12136) <= 16473961;
srom_1(12137) <= 16302034;
srom_1(12138) <= 16092999;
srom_1(12139) <= 15847836;
srom_1(12140) <= 15567693;
srom_1(12141) <= 15253886;
srom_1(12142) <= 14907884;
srom_1(12143) <= 14531312;
srom_1(12144) <= 14125934;
srom_1(12145) <= 13693652;
srom_1(12146) <= 13236493;
srom_1(12147) <= 12756600;
srom_1(12148) <= 12256224;
srom_1(12149) <= 11737712;
srom_1(12150) <= 11203495;
srom_1(12151) <= 10656078;
srom_1(12152) <= 10098027;
srom_1(12153) <= 9531961;
srom_1(12154) <= 8960533;
srom_1(12155) <= 8386423;
srom_1(12156) <= 7812324;
srom_1(12157) <= 7240926;
srom_1(12158) <= 6674911;
srom_1(12159) <= 6116932;
srom_1(12160) <= 5569605;
srom_1(12161) <= 5035498;
srom_1(12162) <= 4517114;
srom_1(12163) <= 4016886;
srom_1(12164) <= 3537157;
srom_1(12165) <= 3080179;
srom_1(12166) <= 2648094;
srom_1(12167) <= 2242928;
srom_1(12168) <= 1866582;
srom_1(12169) <= 1520819;
srom_1(12170) <= 1207262;
srom_1(12171) <= 927381;
srom_1(12172) <= 682487;
srom_1(12173) <= 473731;
srom_1(12174) <= 302090;
srom_1(12175) <= 168370;
srom_1(12176) <= 73197;
srom_1(12177) <= 17017;
srom_1(12178) <= 95;
srom_1(12179) <= 22510;
srom_1(12180) <= 84156;
srom_1(12181) <= 184745;
srom_1(12182) <= 323804;
srom_1(12183) <= 500682;
srom_1(12184) <= 714550;
srom_1(12185) <= 964403;
srom_1(12186) <= 1249071;
srom_1(12187) <= 1567219;
srom_1(12188) <= 1917355;
srom_1(12189) <= 2297836;
srom_1(12190) <= 2706880;
srom_1(12191) <= 3142566;
srom_1(12192) <= 3602854;
srom_1(12193) <= 4085583;
srom_1(12194) <= 4588491;
srom_1(12195) <= 5109219;
srom_1(12196) <= 5645325;
srom_1(12197) <= 6194295;
srom_1(12198) <= 6753555;
srom_1(12199) <= 7320482;
srom_1(12200) <= 7892418;
srom_1(12201) <= 8466681;
srom_1(12202) <= 9040578;
srom_1(12203) <= 9611418;
srom_1(12204) <= 10176523;
srom_1(12205) <= 10733244;
srom_1(12206) <= 11278971;
srom_1(12207) <= 11811143;
srom_1(12208) <= 12327266;
srom_1(12209) <= 12824919;
srom_1(12210) <= 13301769;
srom_1(12211) <= 13755580;
srom_1(12212) <= 14184223;
srom_1(12213) <= 14585688;
srom_1(12214) <= 14958093;
srom_1(12215) <= 15299691;
srom_1(12216) <= 15608881;
srom_1(12217) <= 15884212;
srom_1(12218) <= 16124394;
srom_1(12219) <= 16328301;
srom_1(12220) <= 16494975;
srom_1(12221) <= 16623636;
srom_1(12222) <= 16713680;
srom_1(12223) <= 16764685;
srom_1(12224) <= 16776411;
srom_1(12225) <= 16748804;
srom_1(12226) <= 16681994;
srom_1(12227) <= 16576293;
srom_1(12228) <= 16432196;
srom_1(12229) <= 16250381;
srom_1(12230) <= 16031699;
srom_1(12231) <= 15777177;
srom_1(12232) <= 15488006;
srom_1(12233) <= 15165544;
srom_1(12234) <= 14811303;
srom_1(12235) <= 14426943;
srom_1(12236) <= 14014268;
srom_1(12237) <= 13575212;
srom_1(12238) <= 13111834;
srom_1(12239) <= 12626307;
srom_1(12240) <= 12120909;
srom_1(12241) <= 11598008;
srom_1(12242) <= 11060057;
srom_1(12243) <= 10509579;
srom_1(12244) <= 9949155;
srom_1(12245) <= 9381413;
srom_1(12246) <= 8809015;
srom_1(12247) <= 8234646;
srom_1(12248) <= 7660999;
srom_1(12249) <= 7090764;
srom_1(12250) <= 6526615;
srom_1(12251) <= 5971198;
srom_1(12252) <= 5427116;
srom_1(12253) <= 4896922;
srom_1(12254) <= 4383102;
srom_1(12255) <= 3888065;
srom_1(12256) <= 3414132;
srom_1(12257) <= 2963527;
srom_1(12258) <= 2538361;
srom_1(12259) <= 2140629;
srom_1(12260) <= 1772197;
srom_1(12261) <= 1434791;
srom_1(12262) <= 1129993;
srom_1(12263) <= 859234;
srom_1(12264) <= 623783;
srom_1(12265) <= 424743;
srom_1(12266) <= 263049;
srom_1(12267) <= 139459;
srom_1(12268) <= 54551;
srom_1(12269) <= 8725;
srom_1(12270) <= 2195;
srom_1(12271) <= 34991;
srom_1(12272) <= 106961;
srom_1(12273) <= 217766;
srom_1(12274) <= 366887;
srom_1(12275) <= 553625;
srom_1(12276) <= 777103;
srom_1(12277) <= 1036275;
srom_1(12278) <= 1329924;
srom_1(12279) <= 1656673;
srom_1(12280) <= 2014991;
srom_1(12281) <= 2403197;
srom_1(12282) <= 2819471;
srom_1(12283) <= 3261860;
srom_1(12284) <= 3728291;
srom_1(12285) <= 4216575;
srom_1(12286) <= 4724423;
srom_1(12287) <= 5249454;
srom_1(12288) <= 5789206;
srom_1(12289) <= 6341147;
srom_1(12290) <= 6902689;
srom_1(12291) <= 7471199;
srom_1(12292) <= 8044011;
srom_1(12293) <= 8618439;
srom_1(12294) <= 9191790;
srom_1(12295) <= 9761374;
srom_1(12296) <= 10324520;
srom_1(12297) <= 10878589;
srom_1(12298) <= 11420981;
srom_1(12299) <= 11949153;
srom_1(12300) <= 12460628;
srom_1(12301) <= 12953009;
srom_1(12302) <= 13423985;
srom_1(12303) <= 13871349;
srom_1(12304) <= 14293002;
srom_1(12305) <= 14686968;
srom_1(12306) <= 15051398;
srom_1(12307) <= 15384585;
srom_1(12308) <= 15684964;
srom_1(12309) <= 15951129;
srom_1(12310) <= 16181830;
srom_1(12311) <= 16375987;
srom_1(12312) <= 16532687;
srom_1(12313) <= 16651198;
srom_1(12314) <= 16730962;
srom_1(12315) <= 16771606;
srom_1(12316) <= 16772939;
srom_1(12317) <= 16734955;
srom_1(12318) <= 16657832;
srom_1(12319) <= 16541933;
srom_1(12320) <= 16387799;
srom_1(12321) <= 16196154;
srom_1(12322) <= 15967897;
srom_1(12323) <= 15704098;
srom_1(12324) <= 15405995;
srom_1(12325) <= 15074984;
srom_1(12326) <= 14712619;
srom_1(12327) <= 14320598;
srom_1(12328) <= 13900760;
srom_1(12329) <= 13455074;
srom_1(12330) <= 12985629;
srom_1(12331) <= 12494627;
srom_1(12332) <= 11984371;
srom_1(12333) <= 11457253;
srom_1(12334) <= 10915745;
srom_1(12335) <= 10362386;
srom_1(12336) <= 9799772;
srom_1(12337) <= 9230540;
srom_1(12338) <= 8657360;
srom_1(12339) <= 8082920;
srom_1(12340) <= 7509913;
srom_1(12341) <= 6941027;
srom_1(12342) <= 6378929;
srom_1(12343) <= 5826255;
srom_1(12344) <= 5285597;
srom_1(12345) <= 4759490;
srom_1(12346) <= 4250401;
srom_1(12347) <= 3760717;
srom_1(12348) <= 3292735;
srom_1(12349) <= 2848650;
srom_1(12350) <= 2430543;
srom_1(12351) <= 2040376;
srom_1(12352) <= 1679978;
srom_1(12353) <= 1351039;
srom_1(12354) <= 1055101;
srom_1(12355) <= 793553;
srom_1(12356) <= 567620;
srom_1(12357) <= 378363;
srom_1(12358) <= 226669;
srom_1(12359) <= 113248;
srom_1(12360) <= 38634;
srom_1(12361) <= 3176;
srom_1(12362) <= 7040;
srom_1(12363) <= 50207;
srom_1(12364) <= 132477;
srom_1(12365) <= 253462;
srom_1(12366) <= 412596;
srom_1(12367) <= 609132;
srom_1(12368) <= 842149;
srom_1(12369) <= 1110553;
srom_1(12370) <= 1413087;
srom_1(12371) <= 1748332;
srom_1(12372) <= 2114715;
srom_1(12373) <= 2510518;
srom_1(12374) <= 2933886;
srom_1(12375) <= 3382833;
srom_1(12376) <= 3855253;
srom_1(12377) <= 4348933;
srom_1(12378) <= 4861555;
srom_1(12379) <= 5390717;
srom_1(12380) <= 5933937;
srom_1(12381) <= 6488668;
srom_1(12382) <= 7052309;
srom_1(12383) <= 7622216;
srom_1(12384) <= 8195717;
srom_1(12385) <= 8770122;
srom_1(12386) <= 9342738;
srom_1(12387) <= 9910880;
srom_1(12388) <= 10471883;
srom_1(12389) <= 11023118;
srom_1(12390) <= 11561998;
srom_1(12391) <= 12085997;
srom_1(12392) <= 12592657;
srom_1(12393) <= 13079604;
srom_1(12394) <= 13544553;
srom_1(12395) <= 13985323;
srom_1(12396) <= 14399849;
srom_1(12397) <= 14786186;
srom_1(12398) <= 15142523;
srom_1(12399) <= 15467188;
srom_1(12400) <= 15758659;
srom_1(12401) <= 16015570;
srom_1(12402) <= 16236715;
srom_1(12403) <= 16421057;
srom_1(12404) <= 16567733;
srom_1(12405) <= 16676054;
srom_1(12406) <= 16745512;
srom_1(12407) <= 16775782;
srom_1(12408) <= 16766722;
srom_1(12409) <= 16718373;
srom_1(12410) <= 16630964;
srom_1(12411) <= 16504903;
srom_1(12412) <= 16340782;
srom_1(12413) <= 16139371;
srom_1(12414) <= 15901614;
srom_1(12415) <= 15628625;
srom_1(12416) <= 15321686;
srom_1(12417) <= 14982235;
srom_1(12418) <= 14611864;
srom_1(12419) <= 14212311;
srom_1(12420) <= 13785448;
srom_1(12421) <= 13333277;
srom_1(12422) <= 12857919;
srom_1(12423) <= 12361603;
srom_1(12424) <= 11846656;
srom_1(12425) <= 11315493;
srom_1(12426) <= 10770605;
srom_1(12427) <= 10214547;
srom_1(12428) <= 9649927;
srom_1(12429) <= 9079392;
srom_1(12430) <= 8505617;
srom_1(12431) <= 7931294;
srom_1(12432) <= 7359115;
srom_1(12433) <= 6791764;
srom_1(12434) <= 6231901;
srom_1(12435) <= 5682151;
srom_1(12436) <= 5145093;
srom_1(12437) <= 4623245;
srom_1(12438) <= 4119054;
srom_1(12439) <= 3634885;
srom_1(12440) <= 3173007;
srom_1(12441) <= 2735587;
srom_1(12442) <= 2324676;
srom_1(12443) <= 1942201;
srom_1(12444) <= 1589955;
srom_1(12445) <= 1269591;
srom_1(12446) <= 982610;
srom_1(12447) <= 730358;
srom_1(12448) <= 514018;
srom_1(12449) <= 334605;
srom_1(12450) <= 192960;
srom_1(12451) <= 89748;
srom_1(12452) <= 25451;
srom_1(12453) <= 372;
srom_1(12454) <= 14629;
srom_1(12455) <= 68153;
srom_1(12456) <= 160696;
srom_1(12457) <= 291822;
srom_1(12458) <= 460916;
srom_1(12459) <= 667186;
srom_1(12460) <= 909665;
srom_1(12461) <= 1187215;
srom_1(12462) <= 1498534;
srom_1(12463) <= 1842164;
srom_1(12464) <= 2216492;
srom_1(12465) <= 2619763;
srom_1(12466) <= 3050087;
srom_1(12467) <= 3505444;
srom_1(12468) <= 3983700;
srom_1(12469) <= 4482613;
srom_1(12470) <= 4999842;
srom_1(12471) <= 5532962;
srom_1(12472) <= 6079473;
srom_1(12473) <= 6636812;
srom_1(12474) <= 7202367;
srom_1(12475) <= 7773484;
srom_1(12476) <= 8347485;
srom_1(12477) <= 8921679;
srom_1(12478) <= 9493374;
srom_1(12479) <= 10059888;
srom_1(12480) <= 10618564;
srom_1(12481) <= 11166784;
srom_1(12482) <= 11701976;
srom_1(12483) <= 12221630;
srom_1(12484) <= 12723310;
srom_1(12485) <= 13204663;
srom_1(12486) <= 13663432;
srom_1(12487) <= 14097465;
srom_1(12488) <= 14504728;
srom_1(12489) <= 14883310;
srom_1(12490) <= 15231436;
srom_1(12491) <= 15547474;
srom_1(12492) <= 15829941;
srom_1(12493) <= 16077514;
srom_1(12494) <= 16289030;
srom_1(12495) <= 16463499;
srom_1(12496) <= 16600101;
srom_1(12497) <= 16698197;
srom_1(12498) <= 16757327;
srom_1(12499) <= 16777213;
srom_1(12500) <= 16757762;
srom_1(12501) <= 16699065;
srom_1(12502) <= 16601397;
srom_1(12503) <= 16465217;
srom_1(12504) <= 16291162;
srom_1(12505) <= 16080050;
srom_1(12506) <= 15832871;
srom_1(12507) <= 15550782;
srom_1(12508) <= 15235107;
srom_1(12509) <= 14887327;
srom_1(12510) <= 14509073;
srom_1(12511) <= 14102117;
srom_1(12512) <= 13668368;
srom_1(12513) <= 13209861;
srom_1(12514) <= 12728746;
srom_1(12515) <= 12227278;
srom_1(12516) <= 11707809;
srom_1(12517) <= 11172775;
srom_1(12518) <= 10624686;
srom_1(12519) <= 10066110;
srom_1(12520) <= 9499669;
srom_1(12521) <= 8928017;
srom_1(12522) <= 8353835;
srom_1(12523) <= 7779817;
srom_1(12524) <= 7208654;
srom_1(12525) <= 6643023;
srom_1(12526) <= 6085579;
srom_1(12527) <= 5538934;
srom_1(12528) <= 5005652;
srom_1(12529) <= 4488234;
srom_1(12530) <= 3989106;
srom_1(12531) <= 3510609;
srom_1(12532) <= 3054986;
srom_1(12533) <= 2624375;
srom_1(12534) <= 2220794;
srom_1(12535) <= 1846137;
srom_1(12536) <= 1502159;
srom_1(12537) <= 1190474;
srom_1(12538) <= 912543;
srom_1(12539) <= 669670;
srom_1(12540) <= 462994;
srom_1(12541) <= 293484;
srom_1(12542) <= 161935;
srom_1(12543) <= 68964;
srom_1(12544) <= 15006;
srom_1(12545) <= 315;
srom_1(12546) <= 24959;
srom_1(12547) <= 88824;
srom_1(12548) <= 191608;
srom_1(12549) <= 332832;
srom_1(12550) <= 511832;
srom_1(12551) <= 727769;
srom_1(12552) <= 979630;
srom_1(12553) <= 1266234;
srom_1(12554) <= 1586237;
srom_1(12555) <= 1938139;
srom_1(12556) <= 2320290;
srom_1(12557) <= 2730897;
srom_1(12558) <= 3168035;
srom_1(12559) <= 3629654;
srom_1(12560) <= 4113589;
srom_1(12561) <= 4617572;
srom_1(12562) <= 5139238;
srom_1(12563) <= 5676141;
srom_1(12564) <= 6225765;
srom_1(12565) <= 6785530;
srom_1(12566) <= 7352813;
srom_1(12567) <= 7924953;
srom_1(12568) <= 8499267;
srom_1(12569) <= 9073063;
srom_1(12570) <= 9643648;
srom_1(12571) <= 10208349;
srom_1(12572) <= 10764516;
srom_1(12573) <= 11309541;
srom_1(12574) <= 11840869;
srom_1(12575) <= 12356009;
srom_1(12576) <= 12852544;
srom_1(12577) <= 13328146;
srom_1(12578) <= 13780584;
srom_1(12579) <= 14207738;
srom_1(12580) <= 14607604;
srom_1(12581) <= 14978307;
srom_1(12582) <= 15318109;
srom_1(12583) <= 15625416;
srom_1(12584) <= 15898787;
srom_1(12585) <= 16136940;
srom_1(12586) <= 16338758;
srom_1(12587) <= 16503296;
srom_1(12588) <= 16629781;
srom_1(12589) <= 16717620;
srom_1(12590) <= 16766402;
srom_1(12591) <= 16775897;
srom_1(12592) <= 16746062;
srom_1(12593) <= 16677035;
srom_1(12594) <= 16569141;
srom_1(12595) <= 16422886;
srom_1(12596) <= 16238955;
srom_1(12597) <= 16018212;
srom_1(12598) <= 15761690;
srom_1(12599) <= 15470594;
srom_1(12600) <= 15146287;
srom_1(12601) <= 14790292;
srom_1(12602) <= 14404277;
srom_1(12603) <= 13990052;
srom_1(12604) <= 13549560;
srom_1(12605) <= 13084867;
srom_1(12606) <= 12598152;
srom_1(12607) <= 12091696;
srom_1(12608) <= 11567875;
srom_1(12609) <= 11029146;
srom_1(12610) <= 10478034;
srom_1(12611) <= 9917124;
srom_1(12612) <= 9349047;
srom_1(12613) <= 8776465;
srom_1(12614) <= 8202065;
srom_1(12615) <= 7628540;
srom_1(12616) <= 7058579;
srom_1(12617) <= 6494854;
srom_1(12618) <= 5940011;
srom_1(12619) <= 5396649;
srom_1(12620) <= 4867318;
srom_1(12621) <= 4354499;
srom_1(12622) <= 3860598;
srom_1(12623) <= 3387930;
srom_1(12624) <= 2938712;
srom_1(12625) <= 2515050;
srom_1(12626) <= 2118932;
srom_1(12627) <= 1752214;
srom_1(12628) <= 1416616;
srom_1(12629) <= 1113713;
srom_1(12630) <= 844924;
srom_1(12631) <= 611510;
srom_1(12632) <= 414565;
srom_1(12633) <= 255014;
srom_1(12634) <= 133603;
srom_1(12635) <= 50904;
srom_1(12636) <= 7302;
srom_1(12637) <= 3003;
srom_1(12638) <= 38028;
srom_1(12639) <= 112211;
srom_1(12640) <= 225205;
srom_1(12641) <= 376480;
srom_1(12642) <= 565326;
srom_1(12643) <= 790859;
srom_1(12644) <= 1052020;
srom_1(12645) <= 1347585;
srom_1(12646) <= 1676167;
srom_1(12647) <= 2036227;
srom_1(12648) <= 2426075;
srom_1(12649) <= 2843883;
srom_1(12650) <= 3287693;
srom_1(12651) <= 3755422;
srom_1(12652) <= 4244878;
srom_1(12653) <= 4753765;
srom_1(12654) <= 5279698;
srom_1(12655) <= 5820209;
srom_1(12656) <= 6372764;
srom_1(12657) <= 6934772;
srom_1(12658) <= 7503598;
srom_1(12659) <= 8076574;
srom_1(12660) <= 8651013;
srom_1(12661) <= 9224222;
srom_1(12662) <= 9793512;
srom_1(12663) <= 10356214;
srom_1(12664) <= 10909689;
srom_1(12665) <= 11451342;
srom_1(12666) <= 11978633;
srom_1(12667) <= 12489088;
srom_1(12668) <= 12980316;
srom_1(12669) <= 13450011;
srom_1(12670) <= 13895972;
srom_1(12671) <= 14316106;
srom_1(12672) <= 14708445;
srom_1(12673) <= 15071147;
srom_1(12674) <= 15402513;
srom_1(12675) <= 15700989;
srom_1(12676) <= 15965174;
srom_1(12677) <= 16193830;
srom_1(12678) <= 16385884;
srom_1(12679) <= 16540437;
srom_1(12680) <= 16656763;
srom_1(12681) <= 16734316;
srom_1(12682) <= 16772734;
srom_1(12683) <= 16771835;
srom_1(12684) <= 16731625;
srom_1(12685) <= 16652292;
srom_1(12686) <= 16534207;
srom_1(12687) <= 16377925;
srom_1(12688) <= 16184178;
srom_1(12689) <= 15953875;
srom_1(12690) <= 15688096;
srom_1(12691) <= 15388087;
srom_1(12692) <= 15055255;
srom_1(12693) <= 14691161;
srom_1(12694) <= 14297512;
srom_1(12695) <= 13876154;
srom_1(12696) <= 13429063;
srom_1(12697) <= 12958336;
srom_1(12698) <= 12466179;
srom_1(12699) <= 11954902;
srom_1(12700) <= 11426901;
srom_1(12701) <= 10884652;
srom_1(12702) <= 10330699;
srom_1(12703) <= 9767638;
srom_1(12704) <= 9198111;
srom_1(12705) <= 8624787;
srom_1(12706) <= 8050356;
srom_1(12707) <= 7477511;
srom_1(12708) <= 6908939;
srom_1(12709) <= 6347305;
srom_1(12710) <= 5795244;
srom_1(12711) <= 5255344;
srom_1(12712) <= 4730137;
srom_1(12713) <= 4222085;
srom_1(12714) <= 3733572;
srom_1(12715) <= 3266888;
srom_1(12716) <= 2824222;
srom_1(12717) <= 2407648;
srom_1(12718) <= 2019122;
srom_1(12719) <= 1660464;
srom_1(12720) <= 1333357;
srom_1(12721) <= 1039334;
srom_1(12722) <= 779775;
srom_1(12723) <= 555896;
srom_1(12724) <= 368747;
srom_1(12725) <= 219206;
srom_1(12726) <= 107974;
srom_1(12727) <= 35573;
srom_1(12728) <= 2342;
srom_1(12729) <= 8438;
srom_1(12730) <= 53830;
srom_1(12731) <= 138308;
srom_1(12732) <= 261474;
srom_1(12733) <= 422751;
srom_1(12734) <= 621382;
srom_1(12735) <= 856437;
srom_1(12736) <= 1126812;
srom_1(12737) <= 1431241;
srom_1(12738) <= 1768295;
srom_1(12739) <= 2136394;
srom_1(12740) <= 2533812;
srom_1(12741) <= 2958685;
srom_1(12742) <= 3409020;
srom_1(12743) <= 3882707;
srom_1(12744) <= 4377523;
srom_1(12745) <= 4891149;
srom_1(12746) <= 5421176;
srom_1(12747) <= 5965117;
srom_1(12748) <= 6520424;
srom_1(12749) <= 7084491;
srom_1(12750) <= 7654673;
srom_1(12751) <= 8228297;
srom_1(12752) <= 8802673;
srom_1(12753) <= 9375107;
srom_1(12754) <= 9942915;
srom_1(12755) <= 10503434;
srom_1(12756) <= 11054037;
srom_1(12757) <= 11592140;
srom_1(12758) <= 12115220;
srom_1(12759) <= 12620826;
srom_1(12760) <= 13106585;
srom_1(12761) <= 13570219;
srom_1(12762) <= 14009556;
srom_1(12763) <= 14422533;
srom_1(12764) <= 14807216;
srom_1(12765) <= 15161800;
srom_1(12766) <= 15484621;
srom_1(12767) <= 15774167;
srom_1(12768) <= 16029080;
srom_1(12769) <= 16248164;
srom_1(12770) <= 16430392;
srom_1(12771) <= 16574909;
srom_1(12772) <= 16681037;
srom_1(12773) <= 16748280;
srom_1(12774) <= 16776321;
srom_1(12775) <= 16765029;
srom_1(12776) <= 16714458;
srom_1(12777) <= 16624843;
srom_1(12778) <= 16496606;
srom_1(12779) <= 16330348;
srom_1(12780) <= 16126848;
srom_1(12781) <= 15887061;
srom_1(12782) <= 15612112;
srom_1(12783) <= 15303288;
srom_1(12784) <= 14962040;
srom_1(12785) <= 14589966;
srom_1(12786) <= 14188812;
srom_1(12787) <= 13760459;
srom_1(12788) <= 13306915;
srom_1(12789) <= 12830308;
srom_1(12790) <= 12332872;
srom_1(12791) <= 11816940;
srom_1(12792) <= 11284931;
srom_1(12793) <= 10739341;
srom_1(12794) <= 10182727;
srom_1(12795) <= 9617700;
srom_1(12796) <= 9046909;
srom_1(12797) <= 8473032;
srom_1(12798) <= 7898758;
srom_1(12799) <= 7326781;
srom_1(12800) <= 6759784;
srom_1(12801) <= 6200425;
srom_1(12802) <= 5651327;
srom_1(12803) <= 5115065;
srom_1(12804) <= 4594153;
srom_1(12805) <= 4091036;
srom_1(12806) <= 3608071;
srom_1(12807) <= 3147523;
srom_1(12808) <= 2711553;
srom_1(12809) <= 2302205;
srom_1(12810) <= 1921397;
srom_1(12811) <= 1570917;
srom_1(12812) <= 1252407;
srom_1(12813) <= 967361;
srom_1(12814) <= 717116;
srom_1(12815) <= 502846;
srom_1(12816) <= 325554;
srom_1(12817) <= 186073;
srom_1(12818) <= 85056;
srom_1(12819) <= 22978;
srom_1(12820) <= 128;
srom_1(12821) <= 16615;
srom_1(12822) <= 72362;
srom_1(12823) <= 167106;
srom_1(12824) <= 300403;
srom_1(12825) <= 471629;
srom_1(12826) <= 679981;
srom_1(12827) <= 924480;
srom_1(12828) <= 1203982;
srom_1(12829) <= 1517175;
srom_1(12830) <= 1862590;
srom_1(12831) <= 2238608;
srom_1(12832) <= 2643465;
srom_1(12833) <= 3075264;
srom_1(12834) <= 3531978;
srom_1(12835) <= 4011467;
srom_1(12836) <= 4511482;
srom_1(12837) <= 5029678;
srom_1(12838) <= 5563625;
srom_1(12839) <= 6110819;
srom_1(12840) <= 6668695;
srom_1(12841) <= 7234636;
srom_1(12842) <= 7805988;
srom_1(12843) <= 8380073;
srom_1(12844) <= 8954197;
srom_1(12845) <= 9525669;
srom_1(12846) <= 10091810;
srom_1(12847) <= 10649963;
srom_1(12848) <= 11197512;
srom_1(12849) <= 11731889;
srom_1(12850) <= 12250588;
srom_1(12851) <= 12751177;
srom_1(12852) <= 13231309;
srom_1(12853) <= 13688731;
srom_1(12854) <= 14121299;
srom_1(12855) <= 14526985;
srom_1(12856) <= 14903886;
srom_1(12857) <= 15250234;
srom_1(12858) <= 15564406;
srom_1(12859) <= 15844928;
srom_1(12860) <= 16090485;
srom_1(12861) <= 16299925;
srom_1(12862) <= 16472266;
srom_1(12863) <= 16606700;
srom_1(12864) <= 16702597;
srom_1(12865) <= 16759506;
srom_1(12866) <= 16777162;
srom_1(12867) <= 16755481;
srom_1(12868) <= 16694564;
srom_1(12869) <= 16594698;
srom_1(12870) <= 16456351;
srom_1(12871) <= 16280171;
srom_1(12872) <= 16066985;
srom_1(12873) <= 15817793;
srom_1(12874) <= 15533763;
srom_1(12875) <= 15216226;
srom_1(12876) <= 14866672;
srom_1(12877) <= 14486741;
srom_1(12878) <= 14078213;
srom_1(12879) <= 13643005;
srom_1(12880) <= 13183157;
srom_1(12881) <= 12700826;
srom_1(12882) <= 12198273;
srom_1(12883) <= 11677856;
srom_1(12884) <= 11142014;
srom_1(12885) <= 10593260;
srom_1(12886) <= 10034168;
srom_1(12887) <= 9467360;
srom_1(12888) <= 8895492;
srom_1(12889) <= 8321248;
srom_1(12890) <= 7747320;
srom_1(12891) <= 7176399;
srom_1(12892) <= 6611162;
srom_1(12893) <= 6054261;
srom_1(12894) <= 5508305;
srom_1(12895) <= 4975857;
srom_1(12896) <= 4459412;
srom_1(12897) <= 3961393;
srom_1(12898) <= 3484134;
srom_1(12899) <= 3029874;
srom_1(12900) <= 2600743;
srom_1(12901) <= 2198753;
srom_1(12902) <= 1825790;
srom_1(12903) <= 1483602;
srom_1(12904) <= 1173794;
srom_1(12905) <= 897818;
srom_1(12906) <= 656970;
srom_1(12907) <= 452378;
srom_1(12908) <= 285001;
srom_1(12909) <= 155625;
srom_1(12910) <= 64856;
srom_1(12911) <= 13121;
srom_1(12912) <= 660;
srom_1(12913) <= 27534;
srom_1(12914) <= 93616;
srom_1(12915) <= 198596;
srom_1(12916) <= 341981;
srom_1(12917) <= 523100;
srom_1(12918) <= 741103;
srom_1(12919) <= 994968;
srom_1(12920) <= 1283504;
srom_1(12921) <= 1605358;
srom_1(12922) <= 1959021;
srom_1(12923) <= 2342835;
srom_1(12924) <= 2755000;
srom_1(12925) <= 3193582;
srom_1(12926) <= 3656526;
srom_1(12927) <= 4141660;
srom_1(12928) <= 4646710;
srom_1(12929) <= 5169306;
srom_1(12930) <= 5706999;
srom_1(12931) <= 6257267;
srom_1(12932) <= 6817529;
srom_1(12933) <= 7385159;
srom_1(12934) <= 7957494;
srom_1(12935) <= 8531851;
srom_1(12936) <= 9105536;
srom_1(12937) <= 9675860;
srom_1(12938) <= 10240147;
srom_1(12939) <= 10795751;
srom_1(12940) <= 11340067;
srom_1(12941) <= 11870544;
srom_1(12942) <= 12384692;
srom_1(12943) <= 12880101;
srom_1(12944) <= 13354447;
srom_1(12945) <= 13805508;
srom_1(12946) <= 14231166;
srom_1(12947) <= 14629427;
srom_1(12948) <= 14998423;
srom_1(12949) <= 15336423;
srom_1(12950) <= 15641842;
srom_1(12951) <= 15913248;
srom_1(12952) <= 16149368;
srom_1(12953) <= 16349096;
srom_1(12954) <= 16511494;
srom_1(12955) <= 16635802;
srom_1(12956) <= 16721435;
srom_1(12957) <= 16767993;
srom_1(12958) <= 16775257;
srom_1(12959) <= 16743193;
srom_1(12960) <= 16671951;
srom_1(12961) <= 16561866;
srom_1(12962) <= 16413454;
srom_1(12963) <= 16227411;
srom_1(12964) <= 16004609;
srom_1(12965) <= 15746092;
srom_1(12966) <= 15453074;
srom_1(12967) <= 15126928;
srom_1(12968) <= 14769184;
srom_1(12969) <= 14381520;
srom_1(12970) <= 13965752;
srom_1(12971) <= 13523831;
srom_1(12972) <= 13057829;
srom_1(12973) <= 12569932;
srom_1(12974) <= 12062427;
srom_1(12975) <= 11537695;
srom_1(12976) <= 10998195;
srom_1(12977) <= 10446458;
srom_1(12978) <= 9885071;
srom_1(12979) <= 9316666;
srom_1(12980) <= 8743910;
srom_1(12981) <= 8169487;
srom_1(12982) <= 7596092;
srom_1(12983) <= 7026413;
srom_1(12984) <= 6463122;
srom_1(12985) <= 5908861;
srom_1(12986) <= 5366227;
srom_1(12987) <= 4837767;
srom_1(12988) <= 4325958;
srom_1(12989) <= 3833200;
srom_1(12990) <= 3361803;
srom_1(12991) <= 2913980;
srom_1(12992) <= 2491828;
srom_1(12993) <= 2097329;
srom_1(12994) <= 1732331;
srom_1(12995) <= 1398548;
srom_1(12996) <= 1097542;
srom_1(12997) <= 830728;
srom_1(12998) <= 599354;
srom_1(12999) <= 404508;
srom_1(13000) <= 247101;
srom_1(13001) <= 127873;
srom_1(13002) <= 47382;
srom_1(13003) <= 6006;
srom_1(13004) <= 3939;
srom_1(13005) <= 41190;
srom_1(13006) <= 117586;
srom_1(13007) <= 232767;
srom_1(13008) <= 386193;
srom_1(13009) <= 577146;
srom_1(13010) <= 804729;
srom_1(13011) <= 1067876;
srom_1(13012) <= 1365352;
srom_1(13013) <= 1695762;
srom_1(13014) <= 2057558;
srom_1(13015) <= 2449042;
srom_1(13016) <= 2868379;
srom_1(13017) <= 3313602;
srom_1(13018) <= 3782623;
srom_1(13019) <= 4273244;
srom_1(13020) <= 4783162;
srom_1(13021) <= 5309988;
srom_1(13022) <= 5851251;
srom_1(13023) <= 6404412;
srom_1(13024) <= 6966878;
srom_1(13025) <= 7536011;
srom_1(13026) <= 8109141;
srom_1(13027) <= 8683583;
srom_1(13028) <= 9256641;
srom_1(13029) <= 9825628;
srom_1(13030) <= 10387877;
srom_1(13031) <= 10940751;
srom_1(13032) <= 11481657;
srom_1(13033) <= 12008058;
srom_1(13034) <= 12517487;
srom_1(13035) <= 13007553;
srom_1(13036) <= 13475960;
srom_1(13037) <= 13920511;
srom_1(13038) <= 14339121;
srom_1(13039) <= 14729826;
srom_1(13040) <= 15090796;
srom_1(13041) <= 15420336;
srom_1(13042) <= 15716903;
srom_1(13043) <= 15979104;
srom_1(13044) <= 16205711;
srom_1(13045) <= 16395661;
srom_1(13046) <= 16548063;
srom_1(13047) <= 16662203;
srom_1(13048) <= 16737545;
srom_1(13049) <= 16773735;
srom_1(13050) <= 16770606;
srom_1(13051) <= 16728170;
srom_1(13052) <= 16646626;
srom_1(13053) <= 16526359;
srom_1(13054) <= 16367930;
srom_1(13055) <= 16172084;
srom_1(13056) <= 15939738;
srom_1(13057) <= 15671983;
srom_1(13058) <= 15370073;
srom_1(13059) <= 15035425;
srom_1(13060) <= 14669607;
srom_1(13061) <= 14274336;
srom_1(13062) <= 13851465;
srom_1(13063) <= 13402976;
srom_1(13064) <= 12930973;
srom_1(13065) <= 12437670;
srom_1(13066) <= 11925379;
srom_1(13067) <= 11396503;
srom_1(13068) <= 10853521;
srom_1(13069) <= 10298982;
srom_1(13070) <= 9735483;
srom_1(13071) <= 9165669;
srom_1(13072) <= 8592211;
srom_1(13073) <= 8017798;
srom_1(13074) <= 7445123;
srom_1(13075) <= 6876873;
srom_1(13076) <= 6315713;
srom_1(13077) <= 5764272;
srom_1(13078) <= 5225138;
srom_1(13079) <= 4700839;
srom_1(13080) <= 4193833;
srom_1(13081) <= 3706498;
srom_1(13082) <= 3241118;
srom_1(13083) <= 2799877;
srom_1(13084) <= 2384844;
srom_1(13085) <= 1997964;
srom_1(13086) <= 1641052;
srom_1(13087) <= 1315782;
srom_1(13088) <= 1023678;
srom_1(13089) <= 766111;
srom_1(13090) <= 544289;
srom_1(13091) <= 359252;
srom_1(13092) <= 211867;
srom_1(13093) <= 102825;
srom_1(13094) <= 32638;
srom_1(13095) <= 1636;
srom_1(13096) <= 9962;
srom_1(13097) <= 57579;
srom_1(13098) <= 144263;
srom_1(13099) <= 269608;
srom_1(13100) <= 433025;
srom_1(13101) <= 633749;
srom_1(13102) <= 870838;
srom_1(13103) <= 1143181;
srom_1(13104) <= 1449499;
srom_1(13105) <= 1788358;
srom_1(13106) <= 2158167;
srom_1(13107) <= 2557194;
srom_1(13108) <= 2983565;
srom_1(13109) <= 3435283;
srom_1(13110) <= 3910228;
srom_1(13111) <= 4406174;
srom_1(13112) <= 4920796;
srom_1(13113) <= 5451679;
srom_1(13114) <= 5996334;
srom_1(13115) <= 6552207;
srom_1(13116) <= 7116692;
srom_1(13117) <= 7687141;
srom_1(13118) <= 8260880;
srom_1(13119) <= 8835218;
srom_1(13120) <= 9407461;
srom_1(13121) <= 9974927;
srom_1(13122) <= 10534954;
srom_1(13123) <= 11084915;
srom_1(13124) <= 11622233;
srom_1(13125) <= 12144388;
srom_1(13126) <= 12648930;
srom_1(13127) <= 13133494;
srom_1(13128) <= 13595808;
srom_1(13129) <= 14033703;
srom_1(13130) <= 14445127;
srom_1(13131) <= 14828149;
srom_1(13132) <= 15180974;
srom_1(13133) <= 15501948;
srom_1(13134) <= 15789564;
srom_1(13135) <= 16042475;
srom_1(13136) <= 16259494;
srom_1(13137) <= 16439604;
srom_1(13138) <= 16581961;
srom_1(13139) <= 16685895;
srom_1(13140) <= 16750921;
srom_1(13141) <= 16776733;
srom_1(13142) <= 16763210;
srom_1(13143) <= 16710416;
srom_1(13144) <= 16618598;
srom_1(13145) <= 16488187;
srom_1(13146) <= 16319794;
srom_1(13147) <= 16114209;
srom_1(13148) <= 15872396;
srom_1(13149) <= 15595489;
srom_1(13150) <= 15284786;
srom_1(13151) <= 14941745;
srom_1(13152) <= 14567974;
srom_1(13153) <= 14165226;
srom_1(13154) <= 13735389;
srom_1(13155) <= 13280479;
srom_1(13156) <= 12802630;
srom_1(13157) <= 12304081;
srom_1(13158) <= 11787172;
srom_1(13159) <= 11254326;
srom_1(13160) <= 10708041;
srom_1(13161) <= 10150880;
srom_1(13162) <= 9585455;
srom_1(13163) <= 9014417;
srom_1(13164) <= 8440445;
srom_1(13165) <= 7866229;
srom_1(13166) <= 7294464;
srom_1(13167) <= 6727829;
srom_1(13168) <= 6168982;
srom_1(13169) <= 5620543;
srom_1(13170) <= 5085085;
srom_1(13171) <= 4565119;
srom_1(13172) <= 4063082;
srom_1(13173) <= 3581329;
srom_1(13174) <= 3122118;
srom_1(13175) <= 2687605;
srom_1(13176) <= 2279825;
srom_1(13177) <= 1900691;
srom_1(13178) <= 1551982;
srom_1(13179) <= 1235331;
srom_1(13180) <= 952225;
srom_1(13181) <= 703991;
srom_1(13182) <= 491792;
srom_1(13183) <= 316624;
srom_1(13184) <= 179309;
srom_1(13185) <= 80490;
srom_1(13186) <= 20630;
srom_1(13187) <= 11;
srom_1(13188) <= 18729;
srom_1(13189) <= 76696;
srom_1(13190) <= 173640;
srom_1(13191) <= 309107;
srom_1(13192) <= 482462;
srom_1(13193) <= 692891;
srom_1(13194) <= 939409;
srom_1(13195) <= 1220858;
srom_1(13196) <= 1535919;
srom_1(13197) <= 1883114;
srom_1(13198) <= 2260817;
srom_1(13199) <= 2667254;
srom_1(13200) <= 3100521;
srom_1(13201) <= 3558585;
srom_1(13202) <= 4039300;
srom_1(13203) <= 4540409;
srom_1(13204) <= 5059564;
srom_1(13205) <= 5594330;
srom_1(13206) <= 6142200;
srom_1(13207) <= 6700603;
srom_1(13208) <= 7266923;
srom_1(13209) <= 7838502;
srom_1(13210) <= 8412661;
srom_1(13211) <= 8986707;
srom_1(13212) <= 9557948;
srom_1(13213) <= 10123706;
srom_1(13214) <= 10681327;
srom_1(13215) <= 11228197;
srom_1(13216) <= 11761751;
srom_1(13217) <= 12279488;
srom_1(13218) <= 12778979;
srom_1(13219) <= 13257881;
srom_1(13220) <= 13713950;
srom_1(13221) <= 14145047;
srom_1(13222) <= 14549150;
srom_1(13223) <= 14924364;
srom_1(13224) <= 15268929;
srom_1(13225) <= 15581230;
srom_1(13226) <= 15859803;
srom_1(13227) <= 16103340;
srom_1(13228) <= 16310701;
srom_1(13229) <= 16480912;
srom_1(13230) <= 16613175;
srom_1(13231) <= 16706871;
srom_1(13232) <= 16761560;
srom_1(13233) <= 16776984;
srom_1(13234) <= 16753073;
srom_1(13235) <= 16689938;
srom_1(13236) <= 16587875;
srom_1(13237) <= 16447363;
srom_1(13238) <= 16269061;
srom_1(13239) <= 16053805;
srom_1(13240) <= 15802603;
srom_1(13241) <= 15516635;
srom_1(13242) <= 15197242;
srom_1(13243) <= 14845920;
srom_1(13244) <= 14464317;
srom_1(13245) <= 14054224;
srom_1(13246) <= 13617563;
srom_1(13247) <= 13156381;
srom_1(13248) <= 12672841;
srom_1(13249) <= 12169211;
srom_1(13250) <= 11647853;
srom_1(13251) <= 11111211;
srom_1(13252) <= 10561801;
srom_1(13253) <= 10002201;
srom_1(13254) <= 9435034;
srom_1(13255) <= 8862960;
srom_1(13256) <= 8288662;
srom_1(13257) <= 7714832;
srom_1(13258) <= 7144162;
srom_1(13259) <= 6579328;
srom_1(13260) <= 6022978;
srom_1(13261) <= 5477721;
srom_1(13262) <= 4946114;
srom_1(13263) <= 4430650;
srom_1(13264) <= 3933747;
srom_1(13265) <= 3457733;
srom_1(13266) <= 3004843;
srom_1(13267) <= 2577199;
srom_1(13268) <= 2176806;
srom_1(13269) <= 1805543;
srom_1(13270) <= 1465150;
srom_1(13271) <= 1157223;
srom_1(13272) <= 883207;
srom_1(13273) <= 644386;
srom_1(13274) <= 441880;
srom_1(13275) <= 276640;
srom_1(13276) <= 149439;
srom_1(13277) <= 60875;
srom_1(13278) <= 11362;
srom_1(13279) <= 1133;
srom_1(13280) <= 30235;
srom_1(13281) <= 98533;
srom_1(13282) <= 205706;
srom_1(13283) <= 351252;
srom_1(13284) <= 534487;
srom_1(13285) <= 754553;
srom_1(13286) <= 1010418;
srom_1(13287) <= 1300881;
srom_1(13288) <= 1624581;
srom_1(13289) <= 1980001;
srom_1(13290) <= 2365472;
srom_1(13291) <= 2779188;
srom_1(13292) <= 3219208;
srom_1(13293) <= 3683469;
srom_1(13294) <= 4169795;
srom_1(13295) <= 4675904;
srom_1(13296) <= 5199423;
srom_1(13297) <= 5737897;
srom_1(13298) <= 6288801;
srom_1(13299) <= 6849552;
srom_1(13300) <= 7417520;
srom_1(13301) <= 7990042;
srom_1(13302) <= 8564433;
srom_1(13303) <= 9138000;
srom_1(13304) <= 9708052;
srom_1(13305) <= 10271917;
srom_1(13306) <= 10826950;
srom_1(13307) <= 11370549;
srom_1(13308) <= 11900165;
srom_1(13309) <= 12413314;
srom_1(13310) <= 12907590;
srom_1(13311) <= 13380674;
srom_1(13312) <= 13830349;
srom_1(13313) <= 14254506;
srom_1(13314) <= 14651156;
srom_1(13315) <= 15018438;
srom_1(13316) <= 15354631;
srom_1(13317) <= 15658158;
srom_1(13318) <= 15927595;
srom_1(13319) <= 16161680;
srom_1(13320) <= 16359314;
srom_1(13321) <= 16519570;
srom_1(13322) <= 16641698;
srom_1(13323) <= 16725124;
srom_1(13324) <= 16769457;
srom_1(13325) <= 16774489;
srom_1(13326) <= 16740198;
srom_1(13327) <= 16666742;
srom_1(13328) <= 16554468;
srom_1(13329) <= 16403901;
srom_1(13330) <= 16215748;
srom_1(13331) <= 15990891;
srom_1(13332) <= 15730383;
srom_1(13333) <= 15435448;
srom_1(13334) <= 15107468;
srom_1(13335) <= 14747980;
srom_1(13336) <= 14358672;
srom_1(13337) <= 13941367;
srom_1(13338) <= 13498024;
srom_1(13339) <= 13030721;
srom_1(13340) <= 12541650;
srom_1(13341) <= 12033103;
srom_1(13342) <= 11507467;
srom_1(13343) <= 10967204;
srom_1(13344) <= 10414850;
srom_1(13345) <= 9852994;
srom_1(13346) <= 9284271;
srom_1(13347) <= 8711348;
srom_1(13348) <= 8136912;
srom_1(13349) <= 7563656;
srom_1(13350) <= 6994268;
srom_1(13351) <= 6431419;
srom_1(13352) <= 5877748;
srom_1(13353) <= 5335851;
srom_1(13354) <= 4808269;
srom_1(13355) <= 4297477;
srom_1(13356) <= 3805870;
srom_1(13357) <= 3335753;
srom_1(13358) <= 2889330;
srom_1(13359) <= 2468695;
srom_1(13360) <= 2075821;
srom_1(13361) <= 1712549;
srom_1(13362) <= 1380584;
srom_1(13363) <= 1081482;
srom_1(13364) <= 816646;
srom_1(13365) <= 587317;
srom_1(13366) <= 394570;
srom_1(13367) <= 239311;
srom_1(13368) <= 122267;
srom_1(13369) <= 43986;
srom_1(13370) <= 4836;
srom_1(13371) <= 5001;
srom_1(13372) <= 44479;
srom_1(13373) <= 123085;
srom_1(13374) <= 240452;
srom_1(13375) <= 396028;
srom_1(13376) <= 589083;
srom_1(13377) <= 818714;
srom_1(13378) <= 1083842;
srom_1(13379) <= 1383225;
srom_1(13380) <= 1715459;
srom_1(13381) <= 2078985;
srom_1(13382) <= 2472099;
srom_1(13383) <= 2892958;
srom_1(13384) <= 3339588;
srom_1(13385) <= 3809894;
srom_1(13386) <= 4301671;
srom_1(13387) <= 4812614;
srom_1(13388) <= 5340325;
srom_1(13389) <= 5882331;
srom_1(13390) <= 6436090;
srom_1(13391) <= 6999005;
srom_1(13392) <= 7568436;
srom_1(13393) <= 8141713;
srom_1(13394) <= 8716148;
srom_1(13395) <= 9289047;
srom_1(13396) <= 9857724;
srom_1(13397) <= 10419511;
srom_1(13398) <= 10971775;
srom_1(13399) <= 11511925;
srom_1(13400) <= 12037429;
srom_1(13401) <= 12545823;
srom_1(13402) <= 13034721;
srom_1(13403) <= 13501833;
srom_1(13404) <= 13944967;
srom_1(13405) <= 14362045;
srom_1(13406) <= 14751112;
srom_1(13407) <= 15110343;
srom_1(13408) <= 15438053;
srom_1(13409) <= 15732706;
srom_1(13410) <= 15992920;
srom_1(13411) <= 16217475;
srom_1(13412) <= 16405317;
srom_1(13413) <= 16555566;
srom_1(13414) <= 16667518;
srom_1(13415) <= 16740647;
srom_1(13416) <= 16774610;
srom_1(13417) <= 16769249;
srom_1(13418) <= 16724588;
srom_1(13419) <= 16640836;
srom_1(13420) <= 16518388;
srom_1(13421) <= 16357815;
srom_1(13422) <= 16159873;
srom_1(13423) <= 15925488;
srom_1(13424) <= 15655760;
srom_1(13425) <= 15351954;
srom_1(13426) <= 15015494;
srom_1(13427) <= 14647959;
srom_1(13428) <= 14251072;
srom_1(13429) <= 13826693;
srom_1(13430) <= 13376813;
srom_1(13431) <= 12903542;
srom_1(13432) <= 12409099;
srom_1(13433) <= 11895802;
srom_1(13434) <= 11366059;
srom_1(13435) <= 10822354;
srom_1(13436) <= 10267236;
srom_1(13437) <= 9703308;
srom_1(13438) <= 9133215;
srom_1(13439) <= 8559631;
srom_1(13440) <= 7985244;
srom_1(13441) <= 7412749;
srom_1(13442) <= 6844831;
srom_1(13443) <= 6284151;
srom_1(13444) <= 5733340;
srom_1(13445) <= 5194981;
srom_1(13446) <= 4671597;
srom_1(13447) <= 4165644;
srom_1(13448) <= 3679494;
srom_1(13449) <= 3215426;
srom_1(13450) <= 2775617;
srom_1(13451) <= 2362130;
srom_1(13452) <= 1976902;
srom_1(13453) <= 1621742;
srom_1(13454) <= 1298313;
srom_1(13455) <= 1008133;
srom_1(13456) <= 752563;
srom_1(13457) <= 532801;
srom_1(13458) <= 349878;
srom_1(13459) <= 204651;
srom_1(13460) <= 97801;
srom_1(13461) <= 29829;
srom_1(13462) <= 1055;
srom_1(13463) <= 11613;
srom_1(13464) <= 61454;
srom_1(13465) <= 150343;
srom_1(13466) <= 277865;
srom_1(13467) <= 443420;
srom_1(13468) <= 646233;
srom_1(13469) <= 885353;
srom_1(13470) <= 1159659;
srom_1(13471) <= 1467863;
srom_1(13472) <= 1808521;
srom_1(13473) <= 2180035;
srom_1(13474) <= 2580663;
srom_1(13475) <= 3008527;
srom_1(13476) <= 3461620;
srom_1(13477) <= 3937817;
srom_1(13478) <= 4434886;
srom_1(13479) <= 4950495;
srom_1(13480) <= 5482226;
srom_1(13481) <= 6027586;
srom_1(13482) <= 6584018;
srom_1(13483) <= 7148913;
srom_1(13484) <= 7719620;
srom_1(13485) <= 8293465;
srom_1(13486) <= 8867756;
srom_1(13487) <= 9439800;
srom_1(13488) <= 10006915;
srom_1(13489) <= 10566440;
srom_1(13490) <= 11115754;
srom_1(13491) <= 11652278;
srom_1(13492) <= 12173498;
srom_1(13493) <= 12676970;
srom_1(13494) <= 13160332;
srom_1(13495) <= 13621318;
srom_1(13496) <= 14057765;
srom_1(13497) <= 14467628;
srom_1(13498) <= 14848985;
srom_1(13499) <= 15200046;
srom_1(13500) <= 15519167;
srom_1(13501) <= 15804849;
srom_1(13502) <= 16055755;
srom_1(13503) <= 16270706;
srom_1(13504) <= 16448696;
srom_1(13505) <= 16588889;
srom_1(13506) <= 16690628;
srom_1(13507) <= 16753436;
srom_1(13508) <= 16777019;
srom_1(13509) <= 16761265;
srom_1(13510) <= 16706249;
srom_1(13511) <= 16612229;
srom_1(13512) <= 16479645;
srom_1(13513) <= 16309120;
srom_1(13514) <= 16101453;
srom_1(13515) <= 15857617;
srom_1(13516) <= 15578757;
srom_1(13517) <= 15266180;
srom_1(13518) <= 14921351;
srom_1(13519) <= 14545889;
srom_1(13520) <= 14141552;
srom_1(13521) <= 13710238;
srom_1(13522) <= 13253969;
srom_1(13523) <= 12774885;
srom_1(13524) <= 12275232;
srom_1(13525) <= 11757353;
srom_1(13526) <= 11223677;
srom_1(13527) <= 10676706;
srom_1(13528) <= 10119006;
srom_1(13529) <= 9553191;
srom_1(13530) <= 8981915;
srom_1(13531) <= 8407857;
srom_1(13532) <= 7833709;
srom_1(13533) <= 7262163;
srom_1(13534) <= 6695899;
srom_1(13535) <= 6137572;
srom_1(13536) <= 5589802;
srom_1(13537) <= 5055156;
srom_1(13538) <= 4536142;
srom_1(13539) <= 4035193;
srom_1(13540) <= 3554659;
srom_1(13541) <= 3096793;
srom_1(13542) <= 2663742;
srom_1(13543) <= 2257537;
srom_1(13544) <= 1880083;
srom_1(13545) <= 1533149;
srom_1(13546) <= 1218363;
srom_1(13547) <= 937201;
srom_1(13548) <= 690981;
srom_1(13549) <= 480858;
srom_1(13550) <= 307817;
srom_1(13551) <= 172669;
srom_1(13552) <= 76049;
srom_1(13553) <= 18409;
srom_1(13554) <= 20;
srom_1(13555) <= 20968;
srom_1(13556) <= 81155;
srom_1(13557) <= 180298;
srom_1(13558) <= 317933;
srom_1(13559) <= 493414;
srom_1(13560) <= 705918;
srom_1(13561) <= 954449;
srom_1(13562) <= 1237841;
srom_1(13563) <= 1554766;
srom_1(13564) <= 1903737;
srom_1(13565) <= 2283118;
srom_1(13566) <= 2691129;
srom_1(13567) <= 3125858;
srom_1(13568) <= 3585266;
srom_1(13569) <= 4067198;
srom_1(13570) <= 4569395;
srom_1(13571) <= 5089501;
srom_1(13572) <= 5625078;
srom_1(13573) <= 6173614;
srom_1(13574) <= 6732537;
srom_1(13575) <= 7299226;
srom_1(13576) <= 7871024;
srom_1(13577) <= 8445248;
srom_1(13578) <= 9019207;
srom_1(13579) <= 9590209;
srom_1(13580) <= 10155576;
srom_1(13581) <= 10712657;
srom_1(13582) <= 11258840;
srom_1(13583) <= 11791563;
srom_1(13584) <= 12308329;
srom_1(13585) <= 12806714;
srom_1(13586) <= 13284380;
srom_1(13587) <= 13739089;
srom_1(13588) <= 14168708;
srom_1(13589) <= 14571221;
srom_1(13590) <= 14944743;
srom_1(13591) <= 15287520;
srom_1(13592) <= 15597946;
srom_1(13593) <= 15874565;
srom_1(13594) <= 16116079;
srom_1(13595) <= 16321357;
srom_1(13596) <= 16489436;
srom_1(13597) <= 16619526;
srom_1(13598) <= 16711020;
srom_1(13599) <= 16763486;
srom_1(13600) <= 16776680;
srom_1(13601) <= 16750540;
srom_1(13602) <= 16685187;
srom_1(13603) <= 16580929;
srom_1(13604) <= 16438254;
srom_1(13605) <= 16257832;
srom_1(13606) <= 16040508;
srom_1(13607) <= 15787302;
srom_1(13608) <= 15499401;
srom_1(13609) <= 15178154;
srom_1(13610) <= 14825070;
srom_1(13611) <= 14441802;
srom_1(13612) <= 14030149;
srom_1(13613) <= 13592041;
srom_1(13614) <= 13129532;
srom_1(13615) <= 12644792;
srom_1(13616) <= 12140092;
srom_1(13617) <= 11617801;
srom_1(13618) <= 11080367;
srom_1(13619) <= 10530310;
srom_1(13620) <= 9970210;
srom_1(13621) <= 9402693;
srom_1(13622) <= 8830421;
srom_1(13623) <= 8256077;
srom_1(13624) <= 7682355;
srom_1(13625) <= 7111944;
srom_1(13626) <= 6547521;
srom_1(13627) <= 5991730;
srom_1(13628) <= 5447180;
srom_1(13629) <= 4916423;
srom_1(13630) <= 4401948;
srom_1(13631) <= 3906167;
srom_1(13632) <= 3431407;
srom_1(13633) <= 2979893;
srom_1(13634) <= 2553742;
srom_1(13635) <= 2154952;
srom_1(13636) <= 1785394;
srom_1(13637) <= 1446802;
srom_1(13638) <= 1140761;
srom_1(13639) <= 868708;
srom_1(13640) <= 631919;
srom_1(13641) <= 431503;
srom_1(13642) <= 268401;
srom_1(13643) <= 143378;
srom_1(13644) <= 57019;
srom_1(13645) <= 9730;
srom_1(13646) <= 1732;
srom_1(13647) <= 33063;
srom_1(13648) <= 103576;
srom_1(13649) <= 212941;
srom_1(13650) <= 360644;
srom_1(13651) <= 545993;
srom_1(13652) <= 768118;
srom_1(13653) <= 1025979;
srom_1(13654) <= 1318365;
srom_1(13655) <= 1643907;
srom_1(13656) <= 2001076;
srom_1(13657) <= 2388199;
srom_1(13658) <= 2803460;
srom_1(13659) <= 3244912;
srom_1(13660) <= 3710484;
srom_1(13661) <= 4197993;
srom_1(13662) <= 4705154;
srom_1(13663) <= 5229588;
srom_1(13664) <= 5768835;
srom_1(13665) <= 6320367;
srom_1(13666) <= 6881598;
srom_1(13667) <= 7449896;
srom_1(13668) <= 8022596;
srom_1(13669) <= 8597012;
srom_1(13670) <= 9170451;
srom_1(13671) <= 9740224;
srom_1(13672) <= 10303658;
srom_1(13673) <= 10858112;
srom_1(13674) <= 11400986;
srom_1(13675) <= 11929734;
srom_1(13676) <= 12441876;
srom_1(13677) <= 12935011;
srom_1(13678) <= 13406826;
srom_1(13679) <= 13855109;
srom_1(13680) <= 14277758;
srom_1(13681) <= 14672790;
srom_1(13682) <= 15038354;
srom_1(13683) <= 15372735;
srom_1(13684) <= 15674365;
srom_1(13685) <= 15941829;
srom_1(13686) <= 16173874;
srom_1(13687) <= 16369411;
srom_1(13688) <= 16527523;
srom_1(13689) <= 16647469;
srom_1(13690) <= 16728687;
srom_1(13691) <= 16770795;
srom_1(13692) <= 16773596;
srom_1(13693) <= 16737077;
srom_1(13694) <= 16661409;
srom_1(13695) <= 16546947;
srom_1(13696) <= 16394228;
srom_1(13697) <= 16203967;
srom_1(13698) <= 15977058;
srom_1(13699) <= 15714564;
srom_1(13700) <= 15417716;
srom_1(13701) <= 15087906;
srom_1(13702) <= 14726681;
srom_1(13703) <= 14335734;
srom_1(13704) <= 13916899;
srom_1(13705) <= 13472140;
srom_1(13706) <= 13003543;
srom_1(13707) <= 12513305;
srom_1(13708) <= 12003724;
srom_1(13709) <= 11477191;
srom_1(13710) <= 10936175;
srom_1(13711) <= 10383212;
srom_1(13712) <= 9820896;
srom_1(13713) <= 9251863;
srom_1(13714) <= 8678782;
srom_1(13715) <= 8104341;
srom_1(13716) <= 7531232;
srom_1(13717) <= 6962144;
srom_1(13718) <= 6399745;
srom_1(13719) <= 5846673;
srom_1(13720) <= 5305521;
srom_1(13721) <= 4778826;
srom_1(13722) <= 4269059;
srom_1(13723) <= 3778609;
srom_1(13724) <= 3309778;
srom_1(13725) <= 2864763;
srom_1(13726) <= 2445651;
srom_1(13727) <= 2054408;
srom_1(13728) <= 1692868;
srom_1(13729) <= 1362726;
srom_1(13730) <= 1065532;
srom_1(13731) <= 802678;
srom_1(13732) <= 575396;
srom_1(13733) <= 384754;
srom_1(13734) <= 231644;
srom_1(13735) <= 116786;
srom_1(13736) <= 40716;
srom_1(13737) <= 3793;
srom_1(13738) <= 6189;
srom_1(13739) <= 47893;
srom_1(13740) <= 128710;
srom_1(13741) <= 248260;
srom_1(13742) <= 405983;
srom_1(13743) <= 601139;
srom_1(13744) <= 832813;
srom_1(13745) <= 1099919;
srom_1(13746) <= 1401204;
srom_1(13747) <= 1735256;
srom_1(13748) <= 2100507;
srom_1(13749) <= 2495245;
srom_1(13750) <= 2917620;
srom_1(13751) <= 3365650;
srom_1(13752) <= 3837234;
srom_1(13753) <= 4330161;
srom_1(13754) <= 4842119;
srom_1(13755) <= 5370708;
srom_1(13756) <= 5913450;
srom_1(13757) <= 6467798;
srom_1(13758) <= 7031153;
srom_1(13759) <= 7600874;
srom_1(13760) <= 8174289;
srom_1(13761) <= 8748709;
srom_1(13762) <= 9321440;
srom_1(13763) <= 9889797;
srom_1(13764) <= 10451114;
srom_1(13765) <= 11002759;
srom_1(13766) <= 11542146;
srom_1(13767) <= 12066745;
srom_1(13768) <= 12574096;
srom_1(13769) <= 13061819;
srom_1(13770) <= 13527628;
srom_1(13771) <= 13969339;
srom_1(13772) <= 14384880;
srom_1(13773) <= 14772302;
srom_1(13774) <= 15129788;
srom_1(13775) <= 15455663;
srom_1(13776) <= 15748398;
srom_1(13777) <= 16006621;
srom_1(13778) <= 16229120;
srom_1(13779) <= 16414852;
srom_1(13780) <= 16562946;
srom_1(13781) <= 16672708;
srom_1(13782) <= 16743623;
srom_1(13783) <= 16775359;
srom_1(13784) <= 16767766;
srom_1(13785) <= 16720880;
srom_1(13786) <= 16634922;
srom_1(13787) <= 16510294;
srom_1(13788) <= 16347580;
srom_1(13789) <= 16147544;
srom_1(13790) <= 15911124;
srom_1(13791) <= 15639427;
srom_1(13792) <= 15333730;
srom_1(13793) <= 14995464;
srom_1(13794) <= 14626217;
srom_1(13795) <= 14227719;
srom_1(13796) <= 13801839;
srom_1(13797) <= 13350575;
srom_1(13798) <= 12876043;
srom_1(13799) <= 12380468;
srom_1(13800) <= 11866173;
srom_1(13801) <= 11335571;
srom_1(13802) <= 10791149;
srom_1(13803) <= 10235461;
srom_1(13804) <= 9671113;
srom_1(13805) <= 9100751;
srom_1(13806) <= 8527049;
srom_1(13807) <= 7952697;
srom_1(13808) <= 7380390;
srom_1(13809) <= 6812811;
srom_1(13810) <= 6252621;
srom_1(13811) <= 5702448;
srom_1(13812) <= 5164871;
srom_1(13813) <= 4642411;
srom_1(13814) <= 4137519;
srom_1(13815) <= 3652561;
srom_1(13816) <= 3189812;
srom_1(13817) <= 2751442;
srom_1(13818) <= 2339506;
srom_1(13819) <= 1955937;
srom_1(13820) <= 1602533;
srom_1(13821) <= 1280952;
srom_1(13822) <= 992700;
srom_1(13823) <= 739130;
srom_1(13824) <= 521432;
srom_1(13825) <= 340625;
srom_1(13826) <= 197558;
srom_1(13827) <= 92902;
srom_1(13828) <= 27147;
srom_1(13829) <= 602;
srom_1(13830) <= 13391;
srom_1(13831) <= 65454;
srom_1(13832) <= 156547;
srom_1(13833) <= 286244;
srom_1(13834) <= 453935;
srom_1(13835) <= 658835;
srom_1(13836) <= 899982;
srom_1(13837) <= 1176245;
srom_1(13838) <= 1486331;
srom_1(13839) <= 1828783;
srom_1(13840) <= 2201996;
srom_1(13841) <= 2604221;
srom_1(13842) <= 3033571;
srom_1(13843) <= 3488032;
srom_1(13844) <= 3965474;
srom_1(13845) <= 4463657;
srom_1(13846) <= 4980246;
srom_1(13847) <= 5512817;
srom_1(13848) <= 6058875;
srom_1(13849) <= 6615857;
srom_1(13850) <= 7181152;
srom_1(13851) <= 7752109;
srom_1(13852) <= 8326051;
srom_1(13853) <= 8900287;
srom_1(13854) <= 9472123;
srom_1(13855) <= 10038878;
srom_1(13856) <= 10597894;
srom_1(13857) <= 11146551;
srom_1(13858) <= 11682274;
srom_1(13859) <= 12202552;
srom_1(13860) <= 12704945;
srom_1(13861) <= 13187098;
srom_1(13862) <= 13646749;
srom_1(13863) <= 14081742;
srom_1(13864) <= 14490038;
srom_1(13865) <= 14869723;
srom_1(13866) <= 15219016;
srom_1(13867) <= 15536278;
srom_1(13868) <= 15820022;
srom_1(13869) <= 16068918;
srom_1(13870) <= 16281799;
srom_1(13871) <= 16457665;
srom_1(13872) <= 16595693;
srom_1(13873) <= 16695235;
srom_1(13874) <= 16755825;
srom_1(13875) <= 16777177;
srom_1(13876) <= 16759193;
srom_1(13877) <= 16701956;
srom_1(13878) <= 16605735;
srom_1(13879) <= 16470982;
srom_1(13880) <= 16298327;
srom_1(13881) <= 16088580;
srom_1(13882) <= 15842726;
srom_1(13883) <= 15561917;
srom_1(13884) <= 15247470;
srom_1(13885) <= 14900859;
srom_1(13886) <= 14523710;
srom_1(13887) <= 14117792;
srom_1(13888) <= 13685007;
srom_1(13889) <= 13227386;
srom_1(13890) <= 12747074;
srom_1(13891) <= 12246324;
srom_1(13892) <= 11727483;
srom_1(13893) <= 11192985;
srom_1(13894) <= 10645337;
srom_1(13895) <= 10087106;
srom_1(13896) <= 9520910;
srom_1(13897) <= 8949405;
srom_1(13898) <= 8375269;
srom_1(13899) <= 7801197;
srom_1(13900) <= 7229878;
srom_1(13901) <= 6663994;
srom_1(13902) <= 6106197;
srom_1(13903) <= 5559102;
srom_1(13904) <= 5025277;
srom_1(13905) <= 4507223;
srom_1(13906) <= 4007370;
srom_1(13907) <= 3528062;
srom_1(13908) <= 3071548;
srom_1(13909) <= 2639966;
srom_1(13910) <= 2235342;
srom_1(13911) <= 1859573;
srom_1(13912) <= 1514421;
srom_1(13913) <= 1201504;
srom_1(13914) <= 922290;
srom_1(13915) <= 678087;
srom_1(13916) <= 470043;
srom_1(13917) <= 299131;
srom_1(13918) <= 166153;
srom_1(13919) <= 71734;
srom_1(13920) <= 16315;
srom_1(13921) <= 156;
srom_1(13922) <= 23334;
srom_1(13923) <= 85740;
srom_1(13924) <= 187080;
srom_1(13925) <= 326881;
srom_1(13926) <= 504485;
srom_1(13927) <= 719061;
srom_1(13928) <= 969602;
srom_1(13929) <= 1254933;
srom_1(13930) <= 1573717;
srom_1(13931) <= 1924458;
srom_1(13932) <= 2305511;
srom_1(13933) <= 2715090;
srom_1(13934) <= 3151275;
srom_1(13935) <= 3612018;
srom_1(13936) <= 4095161;
srom_1(13937) <= 4598438;
srom_1(13938) <= 5119488;
srom_1(13939) <= 5655868;
srom_1(13940) <= 6205062;
srom_1(13941) <= 6764496;
srom_1(13942) <= 7331546;
srom_1(13943) <= 7903553;
srom_1(13944) <= 8477835;
srom_1(13945) <= 9051698;
srom_1(13946) <= 9622451;
srom_1(13947) <= 10187419;
srom_1(13948) <= 10743951;
srom_1(13949) <= 11289439;
srom_1(13950) <= 11821323;
srom_1(13951) <= 12337111;
srom_1(13952) <= 12834382;
srom_1(13953) <= 13310805;
srom_1(13954) <= 13764147;
srom_1(13955) <= 14192281;
srom_1(13956) <= 14593200;
srom_1(13957) <= 14965023;
srom_1(13958) <= 15306007;
srom_1(13959) <= 15614553;
srom_1(13960) <= 15889213;
srom_1(13961) <= 16128702;
srom_1(13962) <= 16331894;
srom_1(13963) <= 16497837;
srom_1(13964) <= 16625753;
srom_1(13965) <= 16715043;
srom_1(13966) <= 16765287;
srom_1(13967) <= 16776249;
srom_1(13968) <= 16747880;
srom_1(13969) <= 16680311;
srom_1(13970) <= 16573859;
srom_1(13971) <= 16429023;
srom_1(13972) <= 16246484;
srom_1(13973) <= 16027096;
srom_1(13974) <= 15771889;
srom_1(13975) <= 15482058;
srom_1(13976) <= 15158965;
srom_1(13977) <= 14804122;
srom_1(13978) <= 14419196;
srom_1(13979) <= 14005989;
srom_1(13980) <= 13566441;
srom_1(13981) <= 13102612;
srom_1(13982) <= 12616678;
srom_1(13983) <= 12110916;
srom_1(13984) <= 11587700;
srom_1(13985) <= 11049482;
srom_1(13986) <= 10498786;
srom_1(13987) <= 9938195;
srom_1(13988) <= 9370337;
srom_1(13989) <= 8797875;
srom_1(13990) <= 8223495;
srom_1(13991) <= 7649888;
srom_1(13992) <= 7079746;
srom_1(13993) <= 6515741;
srom_1(13994) <= 5960519;
srom_1(13995) <= 5416683;
srom_1(13996) <= 4886784;
srom_1(13997) <= 4373305;
srom_1(13998) <= 3878656;
srom_1(13999) <= 3405156;
srom_1(14000) <= 2955024;
srom_1(14001) <= 2530373;
srom_1(14002) <= 2133192;
srom_1(14003) <= 1765346;
srom_1(14004) <= 1428558;
srom_1(14005) <= 1124409;
srom_1(14006) <= 854323;
srom_1(14007) <= 619569;
srom_1(14008) <= 421246;
srom_1(14009) <= 260285;
srom_1(14010) <= 137441;
srom_1(14011) <= 53289;
srom_1(14012) <= 8224;
srom_1(14013) <= 2457;
srom_1(14014) <= 36016;
srom_1(14015) <= 108744;
srom_1(14016) <= 220298;
srom_1(14017) <= 370157;
srom_1(14018) <= 557616;
srom_1(14019) <= 781798;
srom_1(14020) <= 1041651;
srom_1(14021) <= 1335956;
srom_1(14022) <= 1663334;
srom_1(14023) <= 2022249;
srom_1(14024) <= 2411017;
srom_1(14025) <= 2827817;
srom_1(14026) <= 3270693;
srom_1(14027) <= 3737569;
srom_1(14028) <= 4226255;
srom_1(14029) <= 4734460;
srom_1(14030) <= 5259800;
srom_1(14031) <= 5799813;
srom_1(14032) <= 6351965;
srom_1(14033) <= 6913667;
srom_1(14034) <= 7482286;
srom_1(14035) <= 8055156;
srom_1(14036) <= 8629589;
srom_1(14037) <= 9202891;
srom_1(14038) <= 9772376;
srom_1(14039) <= 10335371;
srom_1(14040) <= 10889237;
srom_1(14041) <= 11431377;
srom_1(14042) <= 11959249;
srom_1(14043) <= 12470376;
srom_1(14044) <= 12962363;
srom_1(14045) <= 13432902;
srom_1(14046) <= 13879786;
srom_1(14047) <= 14300920;
srom_1(14048) <= 14694329;
srom_1(14049) <= 15058169;
srom_1(14050) <= 15390733;
srom_1(14051) <= 15690461;
srom_1(14052) <= 15955949;
srom_1(14053) <= 16185951;
srom_1(14054) <= 16379388;
srom_1(14055) <= 16535354;
srom_1(14056) <= 16653116;
srom_1(14057) <= 16732124;
srom_1(14058) <= 16772006;
srom_1(14059) <= 16772576;
srom_1(14060) <= 16733830;
srom_1(14061) <= 16655950;
srom_1(14062) <= 16539302;
srom_1(14063) <= 16384433;
srom_1(14064) <= 16192068;
srom_1(14065) <= 15963111;
srom_1(14066) <= 15698634;
srom_1(14067) <= 15399877;
srom_1(14068) <= 15068243;
srom_1(14069) <= 14705285;
srom_1(14070) <= 14312706;
srom_1(14071) <= 13892348;
srom_1(14072) <= 13446180;
srom_1(14073) <= 12976295;
srom_1(14074) <= 12484897;
srom_1(14075) <= 11974291;
srom_1(14076) <= 11446870;
srom_1(14077) <= 10905107;
srom_1(14078) <= 10351544;
srom_1(14079) <= 9788776;
srom_1(14080) <= 9219442;
srom_1(14081) <= 8646212;
srom_1(14082) <= 8071774;
srom_1(14083) <= 7498822;
srom_1(14084) <= 6930042;
srom_1(14085) <= 6368102;
srom_1(14086) <= 5815637;
srom_1(14087) <= 5275237;
srom_1(14088) <= 4749437;
srom_1(14089) <= 4240702;
srom_1(14090) <= 3751419;
srom_1(14091) <= 3283880;
srom_1(14092) <= 2840280;
srom_1(14093) <= 2422697;
srom_1(14094) <= 2033091;
srom_1(14095) <= 1673288;
srom_1(14096) <= 1344975;
srom_1(14097) <= 1049692;
srom_1(14098) <= 788824;
srom_1(14099) <= 563594;
srom_1(14100) <= 375058;
srom_1(14101) <= 224101;
srom_1(14102) <= 111429;
srom_1(14103) <= 37572;
srom_1(14104) <= 2876;
srom_1(14105) <= 7504;
srom_1(14106) <= 51433;
srom_1(14107) <= 134459;
srom_1(14108) <= 256190;
srom_1(14109) <= 416058;
srom_1(14110) <= 613312;
srom_1(14111) <= 847026;
srom_1(14112) <= 1116106;
srom_1(14113) <= 1419289;
srom_1(14114) <= 1755153;
srom_1(14115) <= 2122124;
srom_1(14116) <= 2518481;
srom_1(14117) <= 2942364;
srom_1(14118) <= 3391787;
srom_1(14119) <= 3864642;
srom_1(14120) <= 4358711;
srom_1(14121) <= 4871678;
srom_1(14122) <= 5401137;
srom_1(14123) <= 5944605;
srom_1(14124) <= 6499534;
srom_1(14125) <= 7063321;
srom_1(14126) <= 7633324;
srom_1(14127) <= 8206867;
srom_1(14128) <= 8781264;
srom_1(14129) <= 9353818;
srom_1(14130) <= 9921847;
srom_1(14131) <= 10482686;
srom_1(14132) <= 11033705;
srom_1(14133) <= 11572320;
srom_1(14134) <= 12096005;
srom_1(14135) <= 12602306;
srom_1(14136) <= 13088846;
srom_1(14137) <= 13553346;
srom_1(14138) <= 13993627;
srom_1(14139) <= 14407623;
srom_1(14140) <= 14793395;
srom_1(14141) <= 15149132;
srom_1(14142) <= 15473167;
srom_1(14143) <= 15763980;
srom_1(14144) <= 16020207;
srom_1(14145) <= 16240647;
srom_1(14146) <= 16424266;
srom_1(14147) <= 16570203;
srom_1(14148) <= 16677774;
srom_1(14149) <= 16746474;
srom_1(14150) <= 16775981;
srom_1(14151) <= 16766157;
srom_1(14152) <= 16717047;
srom_1(14153) <= 16628883;
srom_1(14154) <= 16502077;
srom_1(14155) <= 16337225;
srom_1(14156) <= 16135098;
srom_1(14157) <= 15896646;
srom_1(14158) <= 15622986;
srom_1(14159) <= 15315401;
srom_1(14160) <= 14975334;
srom_1(14161) <= 14604380;
srom_1(14162) <= 14204278;
srom_1(14163) <= 13776904;
srom_1(14164) <= 13324263;
srom_1(14165) <= 12848476;
srom_1(14166) <= 12351776;
srom_1(14167) <= 11836491;
srom_1(14168) <= 11305038;
srom_1(14169) <= 10759909;
srom_1(14170) <= 10203659;
srom_1(14171) <= 9638899;
srom_1(14172) <= 9068275;
srom_1(14173) <= 8494464;
srom_1(14174) <= 7920157;
srom_1(14175) <= 7348046;
srom_1(14176) <= 6780815;
srom_1(14177) <= 6221124;
srom_1(14178) <= 5671596;
srom_1(14179) <= 5134810;
srom_1(14180) <= 4613282;
srom_1(14181) <= 4109457;
srom_1(14182) <= 3625699;
srom_1(14183) <= 3164276;
srom_1(14184) <= 2727352;
srom_1(14185) <= 2316975;
srom_1(14186) <= 1935070;
srom_1(14187) <= 1583428;
srom_1(14188) <= 1263697;
srom_1(14189) <= 977378;
srom_1(14190) <= 725813;
srom_1(14191) <= 510181;
srom_1(14192) <= 331494;
srom_1(14193) <= 190589;
srom_1(14194) <= 88128;
srom_1(14195) <= 24590;
srom_1(14196) <= 274;
srom_1(14197) <= 15294;
srom_1(14198) <= 69580;
srom_1(14199) <= 162876;
srom_1(14200) <= 294745;
srom_1(14201) <= 464569;
srom_1(14202) <= 671552;
srom_1(14203) <= 914723;
srom_1(14204) <= 1192941;
srom_1(14205) <= 1504903;
srom_1(14206) <= 1849144;
srom_1(14207) <= 2224051;
srom_1(14208) <= 2627866;
srom_1(14209) <= 3058695;
srom_1(14210) <= 3514517;
srom_1(14211) <= 3993196;
srom_1(14212) <= 4492487;
srom_1(14213) <= 5010048;
srom_1(14214) <= 5543452;
srom_1(14215) <= 6090198;
srom_1(14216) <= 6647722;
srom_1(14217) <= 7213409;
srom_1(14218) <= 7784608;
srom_1(14219) <= 8358639;
srom_1(14220) <= 8932810;
srom_1(14221) <= 9504430;
srom_1(14222) <= 10070816;
srom_1(14223) <= 10629315;
srom_1(14224) <= 11177306;
srom_1(14225) <= 11712220;
srom_1(14226) <= 12231548;
srom_1(14227) <= 12732856;
srom_1(14228) <= 13213791;
srom_1(14229) <= 13672100;
srom_1(14230) <= 14105633;
srom_1(14231) <= 14512356;
srom_1(14232) <= 14890364;
srom_1(14233) <= 15237882;
srom_1(14234) <= 15553281;
srom_1(14235) <= 15835083;
srom_1(14236) <= 16081966;
srom_1(14237) <= 16292772;
srom_1(14238) <= 16466513;
srom_1(14239) <= 16602374;
srom_1(14240) <= 16699717;
srom_1(14241) <= 16758087;
srom_1(14242) <= 16777210;
srom_1(14243) <= 16756995;
srom_1(14244) <= 16697538;
srom_1(14245) <= 16599118;
srom_1(14246) <= 16462196;
srom_1(14247) <= 16287414;
srom_1(14248) <= 16075592;
srom_1(14249) <= 15827723;
srom_1(14250) <= 15544969;
srom_1(14251) <= 15228657;
srom_1(14252) <= 14880269;
srom_1(14253) <= 14501440;
srom_1(14254) <= 14093945;
srom_1(14255) <= 13659696;
srom_1(14256) <= 13200730;
srom_1(14257) <= 12719197;
srom_1(14258) <= 12217357;
srom_1(14259) <= 11697563;
srom_1(14260) <= 11162251;
srom_1(14261) <= 10613934;
srom_1(14262) <= 10055181;
srom_1(14263) <= 9488612;
srom_1(14264) <= 8916886;
srom_1(14265) <= 8342682;
srom_1(14266) <= 7768693;
srom_1(14267) <= 7197612;
srom_1(14268) <= 6632115;
srom_1(14269) <= 6074856;
srom_1(14270) <= 5528446;
srom_1(14271) <= 4995448;
srom_1(14272) <= 4478363;
srom_1(14273) <= 3979613;
srom_1(14274) <= 3501539;
srom_1(14275) <= 3046382;
srom_1(14276) <= 2616277;
srom_1(14277) <= 2213240;
srom_1(14278) <= 1839161;
srom_1(14279) <= 1495796;
srom_1(14280) <= 1184752;
srom_1(14281) <= 907491;
srom_1(14282) <= 665310;
srom_1(14283) <= 459347;
srom_1(14284) <= 290567;
srom_1(14285) <= 159761;
srom_1(14286) <= 67544;
srom_1(14287) <= 14346;
srom_1(14288) <= 419;
srom_1(14289) <= 25826;
srom_1(14290) <= 90450;
srom_1(14291) <= 193986;
srom_1(14292) <= 335950;
srom_1(14293) <= 515675;
srom_1(14294) <= 732319;
srom_1(14295) <= 984867;
srom_1(14296) <= 1272133;
srom_1(14297) <= 1592770;
srom_1(14298) <= 1945276;
srom_1(14299) <= 2327996;
srom_1(14300) <= 2739137;
srom_1(14301) <= 3176770;
srom_1(14302) <= 3638843;
srom_1(14303) <= 4123190;
srom_1(14304) <= 4627538;
srom_1(14305) <= 5149524;
srom_1(14306) <= 5686698;
srom_1(14307) <= 6236543;
srom_1(14308) <= 6796480;
srom_1(14309) <= 7363882;
srom_1(14310) <= 7936090;
srom_1(14311) <= 8510420;
srom_1(14312) <= 9084178;
srom_1(14313) <= 9654675;
srom_1(14314) <= 10219235;
srom_1(14315) <= 10775210;
srom_1(14316) <= 11319994;
srom_1(14317) <= 11851032;
srom_1(14318) <= 12365833;
srom_1(14319) <= 12861983;
srom_1(14320) <= 13337156;
srom_1(14321) <= 13789124;
srom_1(14322) <= 14215767;
srom_1(14323) <= 14615084;
srom_1(14324) <= 14985203;
srom_1(14325) <= 15324389;
srom_1(14326) <= 15631050;
srom_1(14327) <= 15903749;
srom_1(14328) <= 16141207;
srom_1(14329) <= 16342310;
srom_1(14330) <= 16506116;
srom_1(14331) <= 16631856;
srom_1(14332) <= 16718940;
srom_1(14333) <= 16766961;
srom_1(14334) <= 16775692;
srom_1(14335) <= 16745094;
srom_1(14336) <= 16675309;
srom_1(14337) <= 16566665;
srom_1(14338) <= 16419671;
srom_1(14339) <= 16235017;
srom_1(14340) <= 16013569;
srom_1(14341) <= 15756364;
srom_1(14342) <= 15464609;
srom_1(14343) <= 15139673;
srom_1(14344) <= 14783078;
srom_1(14345) <= 14396498;
srom_1(14346) <= 13981745;
srom_1(14347) <= 13540763;
srom_1(14348) <= 13075621;
srom_1(14349) <= 12588500;
srom_1(14350) <= 12081685;
srom_1(14351) <= 11557551;
srom_1(14352) <= 11018557;
srom_1(14353) <= 10467230;
srom_1(14354) <= 9906156;
srom_1(14355) <= 9337966;
srom_1(14356) <= 8765323;
srom_1(14357) <= 8190914;
srom_1(14358) <= 7617433;
srom_1(14359) <= 7047567;
srom_1(14360) <= 6483990;
srom_1(14361) <= 5929345;
srom_1(14362) <= 5386232;
srom_1(14363) <= 4857198;
srom_1(14364) <= 4344724;
srom_1(14365) <= 3851213;
srom_1(14366) <= 3378979;
srom_1(14367) <= 2930238;
srom_1(14368) <= 2507092;
srom_1(14369) <= 2111527;
srom_1(14370) <= 1745398;
srom_1(14371) <= 1410420;
srom_1(14372) <= 1108166;
srom_1(14373) <= 840052;
srom_1(14374) <= 607336;
srom_1(14375) <= 411109;
srom_1(14376) <= 252292;
srom_1(14377) <= 131628;
srom_1(14378) <= 49684;
srom_1(14379) <= 6844;
srom_1(14380) <= 3309;
srom_1(14381) <= 39096;
srom_1(14382) <= 114036;
srom_1(14383) <= 227779;
srom_1(14384) <= 379791;
srom_1(14385) <= 569358;
srom_1(14386) <= 795593;
srom_1(14387) <= 1057434;
srom_1(14388) <= 1353654;
srom_1(14389) <= 1682863;
srom_1(14390) <= 2043517;
srom_1(14391) <= 2433926;
srom_1(14392) <= 2852258;
srom_1(14393) <= 3296552;
srom_1(14394) <= 3764724;
srom_1(14395) <= 4254580;
srom_1(14396) <= 4763821;
srom_1(14397) <= 5290060;
srom_1(14398) <= 5830829;
srom_1(14399) <= 6383593;
srom_1(14400) <= 6945759;
srom_1(14401) <= 7514690;
srom_1(14402) <= 8087720;
srom_1(14403) <= 8662161;
srom_1(14404) <= 9235319;
srom_1(14405) <= 9804507;
srom_1(14406) <= 10367054;
srom_1(14407) <= 10920325;
srom_1(14408) <= 11461723;
srom_1(14409) <= 11988710;
srom_1(14410) <= 12498815;
srom_1(14411) <= 12989646;
srom_1(14412) <= 13458901;
srom_1(14413) <= 13904380;
srom_1(14414) <= 14323993;
srom_1(14415) <= 14715774;
srom_1(14416) <= 15077884;
srom_1(14417) <= 15408625;
srom_1(14418) <= 15706448;
srom_1(14419) <= 15969954;
srom_1(14420) <= 16197910;
srom_1(14421) <= 16389244;
srom_1(14422) <= 16543061;
srom_1(14423) <= 16658639;
srom_1(14424) <= 16735435;
srom_1(14425) <= 16773091;
srom_1(14426) <= 16771429;
srom_1(14427) <= 16730457;
srom_1(14428) <= 16650367;
srom_1(14429) <= 16531535;
srom_1(14430) <= 16374518;
srom_1(14431) <= 16180052;
srom_1(14432) <= 15949049;
srom_1(14433) <= 15682593;
srom_1(14434) <= 15381933;
srom_1(14435) <= 15048479;
srom_1(14436) <= 14683794;
srom_1(14437) <= 14289589;
srom_1(14438) <= 13867713;
srom_1(14439) <= 13420143;
srom_1(14440) <= 12948978;
srom_1(14441) <= 12456428;
srom_1(14442) <= 11944803;
srom_1(14443) <= 11416502;
srom_1(14444) <= 10874001;
srom_1(14445) <= 10319846;
srom_1(14446) <= 9756635;
srom_1(14447) <= 9187008;
srom_1(14448) <= 8613638;
srom_1(14449) <= 8039212;
srom_1(14450) <= 7466425;
srom_1(14451) <= 6897962;
srom_1(14452) <= 6336489;
srom_1(14453) <= 5784639;
srom_1(14454) <= 5245000;
srom_1(14455) <= 4720103;
srom_1(14456) <= 4212408;
srom_1(14457) <= 3724298;
srom_1(14458) <= 3258059;
srom_1(14459) <= 2815880;
srom_1(14460) <= 2399833;
srom_1(14461) <= 2011869;
srom_1(14462) <= 1653809;
srom_1(14463) <= 1327329;
srom_1(14464) <= 1033963;
srom_1(14465) <= 775085;
srom_1(14466) <= 551910;
srom_1(14467) <= 365483;
srom_1(14468) <= 216680;
srom_1(14469) <= 106198;
srom_1(14470) <= 34554;
srom_1(14471) <= 2086;
srom_1(14472) <= 8945;
srom_1(14473) <= 55099;
srom_1(14474) <= 140332;
srom_1(14475) <= 264244;
srom_1(14476) <= 426254;
srom_1(14477) <= 625602;
srom_1(14478) <= 861353;
srom_1(14479) <= 1132402;
srom_1(14480) <= 1437478;
srom_1(14481) <= 1775151;
srom_1(14482) <= 2143836;
srom_1(14483) <= 2541805;
srom_1(14484) <= 2967191;
srom_1(14485) <= 3418001;
srom_1(14486) <= 3892119;
srom_1(14487) <= 4387323;
srom_1(14488) <= 4901290;
srom_1(14489) <= 5431611;
srom_1(14490) <= 5975798;
srom_1(14491) <= 6531299;
srom_1(14492) <= 7095510;
srom_1(14493) <= 7665785;
srom_1(14494) <= 8239449;
srom_1(14495) <= 8813813;
srom_1(14496) <= 9386182;
srom_1(14497) <= 9953874;
srom_1(14498) <= 10514226;
srom_1(14499) <= 11064610;
srom_1(14500) <= 11602445;
srom_1(14501) <= 12125210;
srom_1(14502) <= 12630452;
srom_1(14503) <= 13115803;
srom_1(14504) <= 13578986;
srom_1(14505) <= 14017830;
srom_1(14506) <= 14430277;
srom_1(14507) <= 14814392;
srom_1(14508) <= 15168374;
srom_1(14509) <= 15490564;
srom_1(14510) <= 15779450;
srom_1(14511) <= 16033678;
srom_1(14512) <= 16252055;
srom_1(14513) <= 16433559;
srom_1(14514) <= 16577336;
srom_1(14515) <= 16682714;
srom_1(14516) <= 16749198;
srom_1(14517) <= 16776476;
srom_1(14518) <= 16764421;
srom_1(14519) <= 16713088;
srom_1(14520) <= 16622720;
srom_1(14521) <= 16493738;
srom_1(14522) <= 16326749;
srom_1(14523) <= 16122535;
srom_1(14524) <= 15882055;
srom_1(14525) <= 15606434;
srom_1(14526) <= 15296967;
srom_1(14527) <= 14955105;
srom_1(14528) <= 14582449;
srom_1(14529) <= 14180749;
srom_1(14530) <= 13751887;
srom_1(14531) <= 13297875;
srom_1(14532) <= 12820842;
srom_1(14533) <= 12323025;
srom_1(14534) <= 11806757;
srom_1(14535) <= 11274461;
srom_1(14536) <= 10728632;
srom_1(14537) <= 10171830;
srom_1(14538) <= 9606666;
srom_1(14539) <= 9035789;
srom_1(14540) <= 8461878;
srom_1(14541) <= 7887624;
srom_1(14542) <= 7315718;
srom_1(14543) <= 6748844;
srom_1(14544) <= 6189659;
srom_1(14545) <= 5640786;
srom_1(14546) <= 5104798;
srom_1(14547) <= 4584209;
srom_1(14548) <= 4081461;
srom_1(14549) <= 3598910;
srom_1(14550) <= 3138819;
srom_1(14551) <= 2703347;
srom_1(14552) <= 2294534;
srom_1(14553) <= 1914299;
srom_1(14554) <= 1564424;
srom_1(14555) <= 1246551;
srom_1(14556) <= 962168;
srom_1(14557) <= 712611;
srom_1(14558) <= 499049;
srom_1(14559) <= 322484;
srom_1(14560) <= 183744;
srom_1(14561) <= 83479;
srom_1(14562) <= 22160;
srom_1(14563) <= 74;
srom_1(14564) <= 17325;
srom_1(14565) <= 73831;
srom_1(14566) <= 169328;
srom_1(14567) <= 303369;
srom_1(14568) <= 475324;
srom_1(14569) <= 684386;
srom_1(14570) <= 929577;
srom_1(14571) <= 1209746;
srom_1(14572) <= 1523578;
srom_1(14573) <= 1869604;
srom_1(14574) <= 2246199;
srom_1(14575) <= 2651598;
srom_1(14576) <= 3083899;
srom_1(14577) <= 3541077;
srom_1(14578) <= 4020986;
srom_1(14579) <= 4521376;
srom_1(14580) <= 5039901;
srom_1(14581) <= 5574129;
srom_1(14582) <= 6121556;
srom_1(14583) <= 6679613;
srom_1(14584) <= 7245685;
srom_1(14585) <= 7817116;
srom_1(14586) <= 8391226;
srom_1(14587) <= 8965325;
srom_1(14588) <= 9536719;
srom_1(14589) <= 10102730;
srom_1(14590) <= 10660702;
srom_1(14591) <= 11208019;
srom_1(14592) <= 11742116;
srom_1(14593) <= 12260486;
srom_1(14594) <= 12760700;
srom_1(14595) <= 13240412;
srom_1(14596) <= 13697372;
srom_1(14597) <= 14129437;
srom_1(14598) <= 14534582;
srom_1(14599) <= 14910906;
srom_1(14600) <= 15256645;
srom_1(14601) <= 15570177;
srom_1(14602) <= 15850032;
srom_1(14603) <= 16094898;
srom_1(14604) <= 16303627;
srom_1(14605) <= 16475239;
srom_1(14606) <= 16608931;
srom_1(14607) <= 16704074;
srom_1(14608) <= 16760223;
srom_1(14609) <= 16777115;
srom_1(14610) <= 16754671;
srom_1(14611) <= 16692995;
srom_1(14612) <= 16592377;
srom_1(14613) <= 16453288;
srom_1(14614) <= 16276382;
srom_1(14615) <= 16062487;
srom_1(14616) <= 15812607;
srom_1(14617) <= 15527913;
srom_1(14618) <= 15209740;
srom_1(14619) <= 14859580;
srom_1(14620) <= 14479076;
srom_1(14621) <= 14070012;
srom_1(14622) <= 13634306;
srom_1(14623) <= 13174001;
srom_1(14624) <= 12691255;
srom_1(14625) <= 12188333;
srom_1(14626) <= 11667592;
srom_1(14627) <= 11131476;
srom_1(14628) <= 10582497;
srom_1(14629) <= 10023230;
srom_1(14630) <= 9456298;
srom_1(14631) <= 8884359;
srom_1(14632) <= 8310095;
srom_1(14633) <= 7736199;
srom_1(14634) <= 7165363;
srom_1(14635) <= 6600263;
srom_1(14636) <= 6043549;
srom_1(14637) <= 5497832;
srom_1(14638) <= 4965671;
srom_1(14639) <= 4449561;
srom_1(14640) <= 3951923;
srom_1(14641) <= 3475090;
srom_1(14642) <= 3021298;
srom_1(14643) <= 2592675;
srom_1(14644) <= 2191231;
srom_1(14645) <= 1818849;
srom_1(14646) <= 1477275;
srom_1(14647) <= 1168110;
srom_1(14648) <= 892805;
srom_1(14649) <= 652650;
srom_1(14650) <= 448771;
srom_1(14651) <= 282126;
srom_1(14652) <= 153494;
srom_1(14653) <= 63479;
srom_1(14654) <= 12504;
srom_1(14655) <= 808;
srom_1(14656) <= 28445;
srom_1(14657) <= 95285;
srom_1(14658) <= 201015;
srom_1(14659) <= 345141;
srom_1(14660) <= 526984;
srom_1(14661) <= 745694;
srom_1(14662) <= 1000243;
srom_1(14663) <= 1289439;
srom_1(14664) <= 1611926;
srom_1(14665) <= 1966191;
srom_1(14666) <= 2350573;
srom_1(14667) <= 2763269;
srom_1(14668) <= 3202344;
srom_1(14669) <= 3665740;
srom_1(14670) <= 4151282;
srom_1(14671) <= 4656695;
srom_1(14672) <= 5179609;
srom_1(14673) <= 5717570;
srom_1(14674) <= 6268056;
srom_1(14675) <= 6828487;
srom_1(14676) <= 7396234;
srom_1(14677) <= 7968634;
srom_1(14678) <= 8543003;
srom_1(14679) <= 9116649;
srom_1(14680) <= 9686880;
srom_1(14681) <= 10251024;
srom_1(14682) <= 10806434;
srom_1(14683) <= 11350505;
srom_1(14684) <= 11880688;
srom_1(14685) <= 12394495;
srom_1(14686) <= 12889517;
srom_1(14687) <= 13363432;
srom_1(14688) <= 13814019;
srom_1(14689) <= 14239165;
srom_1(14690) <= 14636875;
srom_1(14691) <= 15005285;
srom_1(14692) <= 15342667;
srom_1(14693) <= 15647439;
srom_1(14694) <= 15918171;
srom_1(14695) <= 16153595;
srom_1(14696) <= 16352607;
srom_1(14697) <= 16514272;
srom_1(14698) <= 16637834;
srom_1(14699) <= 16722712;
srom_1(14700) <= 16768508;
srom_1(14701) <= 16775008;
srom_1(14702) <= 16742182;
srom_1(14703) <= 16670182;
srom_1(14704) <= 16559348;
srom_1(14705) <= 16410198;
srom_1(14706) <= 16223432;
srom_1(14707) <= 15999926;
srom_1(14708) <= 15740728;
srom_1(14709) <= 15447053;
srom_1(14710) <= 15120279;
srom_1(14711) <= 14761938;
srom_1(14712) <= 14373710;
srom_1(14713) <= 13957415;
srom_1(14714) <= 13515007;
srom_1(14715) <= 13048559;
srom_1(14716) <= 12560259;
srom_1(14717) <= 12052397;
srom_1(14718) <= 11527354;
srom_1(14719) <= 10987592;
srom_1(14720) <= 10435643;
srom_1(14721) <= 9874095;
srom_1(14722) <= 9305580;
srom_1(14723) <= 8732766;
srom_1(14724) <= 8158337;
srom_1(14725) <= 7584989;
srom_1(14726) <= 7015409;
srom_1(14727) <= 6452268;
srom_1(14728) <= 5898207;
srom_1(14729) <= 5355825;
srom_1(14730) <= 4827665;
srom_1(14731) <= 4316203;
srom_1(14732) <= 3823838;
srom_1(14733) <= 3352878;
srom_1(14734) <= 2905533;
srom_1(14735) <= 2483900;
srom_1(14736) <= 2089957;
srom_1(14737) <= 1725549;
srom_1(14738) <= 1392387;
srom_1(14739) <= 1092033;
srom_1(14740) <= 825895;
srom_1(14741) <= 595221;
srom_1(14742) <= 401093;
srom_1(14743) <= 244421;
srom_1(14744) <= 125940;
srom_1(14745) <= 46205;
srom_1(14746) <= 5591;
srom_1(14747) <= 4288;
srom_1(14748) <= 42302;
srom_1(14749) <= 119454;
srom_1(14750) <= 235383;
srom_1(14751) <= 389546;
srom_1(14752) <= 581218;
srom_1(14753) <= 809503;
srom_1(14754) <= 1073328;
srom_1(14755) <= 1371457;
srom_1(14756) <= 1702492;
srom_1(14757) <= 2064881;
srom_1(14758) <= 2456924;
srom_1(14759) <= 2876782;
srom_1(14760) <= 3322487;
srom_1(14761) <= 3791949;
srom_1(14762) <= 4282966;
srom_1(14763) <= 4793237;
srom_1(14764) <= 5320366;
srom_1(14765) <= 5861884;
srom_1(14766) <= 6415251;
srom_1(14767) <= 6977872;
srom_1(14768) <= 7547107;
srom_1(14769) <= 8120289;
srom_1(14770) <= 8694729;
srom_1(14771) <= 9267734;
srom_1(14772) <= 9836616;
srom_1(14773) <= 10398708;
srom_1(14774) <= 10951374;
srom_1(14775) <= 11492022;
srom_1(14776) <= 12018117;
srom_1(14777) <= 12527192;
srom_1(14778) <= 13016860;
srom_1(14779) <= 13484824;
srom_1(14780) <= 13928891;
srom_1(14781) <= 14346977;
srom_1(14782) <= 14737122;
srom_1(14783) <= 15097497;
srom_1(14784) <= 15426412;
srom_1(14785) <= 15722324;
srom_1(14786) <= 15983846;
srom_1(14787) <= 16209751;
srom_1(14788) <= 16398980;
srom_1(14789) <= 16550645;
srom_1(14790) <= 16664036;
srom_1(14791) <= 16738621;
srom_1(14792) <= 16774049;
srom_1(14793) <= 16770155;
srom_1(14794) <= 16726958;
srom_1(14795) <= 16644659;
srom_1(14796) <= 16523644;
srom_1(14797) <= 16364482;
srom_1(14798) <= 16167918;
srom_1(14799) <= 15934874;
srom_1(14800) <= 15666443;
srom_1(14801) <= 15363883;
srom_1(14802) <= 15028615;
srom_1(14803) <= 14662209;
srom_1(14804) <= 14266383;
srom_1(14805) <= 13842995;
srom_1(14806) <= 13394030;
srom_1(14807) <= 12921592;
srom_1(14808) <= 12427898;
srom_1(14809) <= 11915262;
srom_1(14810) <= 11386088;
srom_1(14811) <= 10842858;
srom_1(14812) <= 10288119;
srom_1(14813) <= 9724473;
srom_1(14814) <= 9154562;
srom_1(14815) <= 8581060;
srom_1(14816) <= 8006655;
srom_1(14817) <= 7434041;
srom_1(14818) <= 6865904;
srom_1(14819) <= 6304907;
srom_1(14820) <= 5753681;
srom_1(14821) <= 5214811;
srom_1(14822) <= 4690824;
srom_1(14823) <= 4184178;
srom_1(14824) <= 3697247;
srom_1(14825) <= 3232316;
srom_1(14826) <= 2791564;
srom_1(14827) <= 2377059;
srom_1(14828) <= 1990744;
srom_1(14829) <= 1634431;
srom_1(14830) <= 1309791;
srom_1(14831) <= 1018345;
srom_1(14832) <= 761461;
srom_1(14833) <= 540344;
srom_1(14834) <= 356030;
srom_1(14835) <= 209383;
srom_1(14836) <= 101091;
srom_1(14837) <= 31663;
srom_1(14838) <= 1423;
srom_1(14839) <= 10513;
srom_1(14840) <= 58891;
srom_1(14841) <= 146330;
srom_1(14842) <= 272420;
srom_1(14843) <= 436570;
srom_1(14844) <= 638009;
srom_1(14845) <= 875793;
srom_1(14846) <= 1148808;
srom_1(14847) <= 1455773;
srom_1(14848) <= 1795248;
srom_1(14849) <= 2165641;
srom_1(14850) <= 2565217;
srom_1(14851) <= 2992100;
srom_1(14852) <= 3444289;
srom_1(14853) <= 3919664;
srom_1(14854) <= 4415995;
srom_1(14855) <= 4930955;
srom_1(14856) <= 5462129;
srom_1(14857) <= 6007026;
srom_1(14858) <= 6563092;
srom_1(14859) <= 7127718;
srom_1(14860) <= 7698257;
srom_1(14861) <= 8272033;
srom_1(14862) <= 8846355;
srom_1(14863) <= 9418531;
srom_1(14864) <= 9985878;
srom_1(14865) <= 10545734;
srom_1(14866) <= 11095475;
srom_1(14867) <= 11632522;
srom_1(14868) <= 12154358;
srom_1(14869) <= 12658534;
srom_1(14870) <= 13142688;
srom_1(14871) <= 13604548;
srom_1(14872) <= 14041948;
srom_1(14873) <= 14452838;
srom_1(14874) <= 14835291;
srom_1(14875) <= 15187513;
srom_1(14876) <= 15507853;
srom_1(14877) <= 15794808;
srom_1(14878) <= 16047033;
srom_1(14879) <= 16263345;
srom_1(14880) <= 16442730;
srom_1(14881) <= 16584346;
srom_1(14882) <= 16687529;
srom_1(14883) <= 16751796;
srom_1(14884) <= 16776845;
srom_1(14885) <= 16762559;
srom_1(14886) <= 16709004;
srom_1(14887) <= 16616432;
srom_1(14888) <= 16485277;
srom_1(14889) <= 16316154;
srom_1(14890) <= 16109856;
srom_1(14891) <= 15867350;
srom_1(14892) <= 15589774;
srom_1(14893) <= 15278430;
srom_1(14894) <= 14934776;
srom_1(14895) <= 14560425;
srom_1(14896) <= 14157133;
srom_1(14897) <= 13726790;
srom_1(14898) <= 13271414;
srom_1(14899) <= 12793141;
srom_1(14900) <= 12294214;
srom_1(14901) <= 11776972;
srom_1(14902) <= 11243841;
srom_1(14903) <= 10697320;
srom_1(14904) <= 10139973;
srom_1(14905) <= 9574414;
srom_1(14906) <= 9003294;
srom_1(14907) <= 8429291;
srom_1(14908) <= 7855098;
srom_1(14909) <= 7283406;
srom_1(14910) <= 6716897;
srom_1(14911) <= 6158228;
srom_1(14912) <= 5610017;
srom_1(14913) <= 5074836;
srom_1(14914) <= 4555194;
srom_1(14915) <= 4053529;
srom_1(14916) <= 3572192;
srom_1(14917) <= 3113441;
srom_1(14918) <= 2679428;
srom_1(14919) <= 2272186;
srom_1(14920) <= 1893627;
srom_1(14921) <= 1545524;
srom_1(14922) <= 1229512;
srom_1(14923) <= 947070;
srom_1(14924) <= 699525;
srom_1(14925) <= 488036;
srom_1(14926) <= 313596;
srom_1(14927) <= 177022;
srom_1(14928) <= 78956;
srom_1(14929) <= 19856;
srom_1(14930) <= 0;
srom_1(14931) <= 19481;
srom_1(14932) <= 78208;
srom_1(14933) <= 175905;
srom_1(14934) <= 312114;
srom_1(14935) <= 486197;
srom_1(14936) <= 697337;
srom_1(14937) <= 944544;
srom_1(14938) <= 1226658;
srom_1(14939) <= 1542358;
srom_1(14940) <= 1890162;
srom_1(14941) <= 2268439;
srom_1(14942) <= 2675416;
srom_1(14943) <= 3109184;
srom_1(14944) <= 3567709;
srom_1(14945) <= 4048841;
srom_1(14946) <= 4550323;
srom_1(14947) <= 5069805;
srom_1(14948) <= 5604850;
srom_1(14949) <= 6152948;
srom_1(14950) <= 6711530;
srom_1(14951) <= 7277977;
srom_1(14952) <= 7849632;
srom_1(14953) <= 8423814;
srom_1(14954) <= 8997831;
srom_1(14955) <= 9568992;
srom_1(14956) <= 10134617;
srom_1(14957) <= 10692054;
srom_1(14958) <= 11238690;
srom_1(14959) <= 11771961;
srom_1(14960) <= 12289366;
srom_1(14961) <= 12788479;
srom_1(14962) <= 13266959;
srom_1(14963) <= 13722564;
srom_1(14964) <= 14153155;
srom_1(14965) <= 14556715;
srom_1(14966) <= 14931350;
srom_1(14967) <= 15275304;
srom_1(14968) <= 15586964;
srom_1(14969) <= 15864868;
srom_1(14970) <= 16107714;
srom_1(14971) <= 16314362;
srom_1(14972) <= 16483843;
srom_1(14973) <= 16615363;
srom_1(14974) <= 16708305;
srom_1(14975) <= 16762233;
srom_1(14976) <= 16776895;
srom_1(14977) <= 16752220;
srom_1(14978) <= 16688326;
srom_1(14979) <= 16585512;
srom_1(14980) <= 16444259;
srom_1(14981) <= 16265231;
srom_1(14982) <= 16049267;
srom_1(14983) <= 15797379;
srom_1(14984) <= 15510749;
srom_1(14985) <= 15190720;
srom_1(14986) <= 14838794;
srom_1(14987) <= 14456622;
srom_1(14988) <= 14045994;
srom_1(14989) <= 13608836;
srom_1(14990) <= 13147199;
srom_1(14991) <= 12663248;
srom_1(14992) <= 12159251;
srom_1(14993) <= 11637573;
srom_1(14994) <= 11100658;
srom_1(14995) <= 10551027;
srom_1(14996) <= 9991254;
srom_1(14997) <= 9423967;
srom_1(14998) <= 8851824;
srom_1(14999) <= 8277509;
srom_1(15000) <= 7703715;
srom_1(15001) <= 7133133;
srom_1(15002) <= 6568438;
srom_1(15003) <= 6012279;
srom_1(15004) <= 5467263;
srom_1(15005) <= 4935946;
srom_1(15006) <= 4420819;
srom_1(15007) <= 3924300;
srom_1(15008) <= 3448714;
srom_1(15009) <= 2996294;
srom_1(15010) <= 2569160;
srom_1(15011) <= 2169316;
srom_1(15012) <= 1798635;
srom_1(15013) <= 1458858;
srom_1(15014) <= 1151576;
srom_1(15015) <= 878232;
srom_1(15016) <= 640106;
srom_1(15017) <= 438315;
srom_1(15018) <= 273806;
srom_1(15019) <= 147351;
srom_1(15020) <= 59541;
srom_1(15021) <= 10789;
srom_1(15022) <= 1324;
srom_1(15023) <= 31189;
srom_1(15024) <= 100245;
srom_1(15025) <= 208169;
srom_1(15026) <= 354453;
srom_1(15027) <= 538412;
srom_1(15028) <= 759183;
srom_1(15029) <= 1015731;
srom_1(15030) <= 1306853;
srom_1(15031) <= 1631184;
srom_1(15032) <= 1987203;
srom_1(15033) <= 2373241;
srom_1(15034) <= 2787486;
srom_1(15035) <= 3227997;
srom_1(15036) <= 3692708;
srom_1(15037) <= 4179439;
srom_1(15038) <= 4685909;
srom_1(15039) <= 5209742;
srom_1(15040) <= 5748482;
srom_1(15041) <= 6299602;
srom_1(15042) <= 6860518;
srom_1(15043) <= 7428600;
srom_1(15044) <= 8001184;
srom_1(15045) <= 8575584;
srom_1(15046) <= 9149108;
srom_1(15047) <= 9719065;
srom_1(15048) <= 10282784;
srom_1(15049) <= 10837620;
srom_1(15050) <= 11380972;
srom_1(15051) <= 11910291;
srom_1(15052) <= 12423097;
srom_1(15053) <= 12916983;
srom_1(15054) <= 13389634;
srom_1(15055) <= 13838833;
srom_1(15056) <= 14262474;
srom_1(15057) <= 14658571;
srom_1(15058) <= 15025266;
srom_1(15059) <= 15360839;
srom_1(15060) <= 15663717;
srom_1(15061) <= 15932480;
srom_1(15062) <= 16165867;
srom_1(15063) <= 16362783;
srom_1(15064) <= 16522306;
srom_1(15065) <= 16643687;
srom_1(15066) <= 16726357;
srom_1(15067) <= 16769929;
srom_1(15068) <= 16774198;
srom_1(15069) <= 16739144;
srom_1(15070) <= 16664931;
srom_1(15071) <= 16551908;
srom_1(15072) <= 16400604;
srom_1(15073) <= 16211729;
srom_1(15074) <= 15986169;
srom_1(15075) <= 15724981;
srom_1(15076) <= 15429391;
srom_1(15077) <= 15100784;
srom_1(15078) <= 14740701;
srom_1(15079) <= 14350831;
srom_1(15080) <= 13933002;
srom_1(15081) <= 13489174;
srom_1(15082) <= 13021427;
srom_1(15083) <= 12531955;
srom_1(15084) <= 12023054;
srom_1(15085) <= 11497110;
srom_1(15086) <= 10956588;
srom_1(15087) <= 10404025;
srom_1(15088) <= 9842011;
srom_1(15089) <= 9273181;
srom_1(15090) <= 8700203;
srom_1(15091) <= 8125764;
srom_1(15092) <= 7552557;
srom_1(15093) <= 6983271;
srom_1(15094) <= 6420575;
srom_1(15095) <= 5867108;
srom_1(15096) <= 5325465;
srom_1(15097) <= 4798186;
srom_1(15098) <= 4287744;
srom_1(15099) <= 3796532;
srom_1(15100) <= 3326854;
srom_1(15101) <= 2880912;
srom_1(15102) <= 2460798;
srom_1(15103) <= 2068481;
srom_1(15104) <= 1705802;
srom_1(15105) <= 1374460;
srom_1(15106) <= 1076010;
srom_1(15107) <= 811852;
srom_1(15108) <= 583223;
srom_1(15109) <= 391197;
srom_1(15110) <= 236673;
srom_1(15111) <= 120377;
srom_1(15112) <= 42853;
srom_1(15113) <= 4465;
srom_1(15114) <= 5393;
srom_1(15115) <= 45633;
srom_1(15116) <= 124996;
srom_1(15117) <= 243110;
srom_1(15118) <= 399421;
srom_1(15119) <= 593196;
srom_1(15120) <= 823527;
srom_1(15121) <= 1089332;
srom_1(15122) <= 1389367;
srom_1(15123) <= 1722223;
srom_1(15124) <= 2086341;
srom_1(15125) <= 2480011;
srom_1(15126) <= 2901390;
srom_1(15127) <= 3348499;
srom_1(15128) <= 3819244;
srom_1(15129) <= 4311415;
srom_1(15130) <= 4822706;
srom_1(15131) <= 5350719;
srom_1(15132) <= 5892978;
srom_1(15133) <= 6446939;
srom_1(15134) <= 7010006;
srom_1(15135) <= 7579537;
srom_1(15136) <= 8152862;
srom_1(15137) <= 8727293;
srom_1(15138) <= 9300136;
srom_1(15139) <= 9868704;
srom_1(15140) <= 10430331;
srom_1(15141) <= 10982384;
srom_1(15142) <= 11522274;
srom_1(15143) <= 12047469;
srom_1(15144) <= 12555507;
srom_1(15145) <= 13044004;
srom_1(15146) <= 13510671;
srom_1(15147) <= 13953318;
srom_1(15148) <= 14369871;
srom_1(15149) <= 14758375;
srom_1(15150) <= 15117010;
srom_1(15151) <= 15444092;
srom_1(15152) <= 15738089;
srom_1(15153) <= 15997622;
srom_1(15154) <= 16221474;
srom_1(15155) <= 16408594;
srom_1(15156) <= 16558106;
srom_1(15157) <= 16669309;
srom_1(15158) <= 16741680;
srom_1(15159) <= 16774881;
srom_1(15160) <= 16768756;
srom_1(15161) <= 16723333;
srom_1(15162) <= 16638826;
srom_1(15163) <= 16515631;
srom_1(15164) <= 16354326;
srom_1(15165) <= 16155666;
srom_1(15166) <= 15920584;
srom_1(15167) <= 15650182;
srom_1(15168) <= 15345728;
srom_1(15169) <= 15008650;
srom_1(15170) <= 14640528;
srom_1(15171) <= 14243089;
srom_1(15172) <= 13818196;
srom_1(15173) <= 13367841;
srom_1(15174) <= 12894138;
srom_1(15175) <= 12399306;
srom_1(15176) <= 11885667;
srom_1(15177) <= 11355629;
srom_1(15178) <= 10811678;
srom_1(15179) <= 10256364;
srom_1(15180) <= 9692291;
srom_1(15181) <= 9122105;
srom_1(15182) <= 8548479;
srom_1(15183) <= 7974104;
srom_1(15184) <= 7401672;
srom_1(15185) <= 6833869;
srom_1(15186) <= 6273356;
srom_1(15187) <= 5722762;
srom_1(15188) <= 5184670;
srom_1(15189) <= 4661601;
srom_1(15190) <= 4156010;
srom_1(15191) <= 3670267;
srom_1(15192) <= 3206650;
srom_1(15193) <= 2767333;
srom_1(15194) <= 2354376;
srom_1(15195) <= 1969716;
srom_1(15196) <= 1615156;
srom_1(15197) <= 1292359;
srom_1(15198) <= 1002839;
srom_1(15199) <= 747953;
srom_1(15200) <= 528896;
srom_1(15201) <= 346697;
srom_1(15202) <= 202209;
srom_1(15203) <= 96110;
srom_1(15204) <= 28897;
srom_1(15205) <= 886;
srom_1(15206) <= 12207;
srom_1(15207) <= 62809;
srom_1(15208) <= 152453;
srom_1(15209) <= 280719;
srom_1(15210) <= 447006;
srom_1(15211) <= 650533;
srom_1(15212) <= 890347;
srom_1(15213) <= 1165323;
srom_1(15214) <= 1474172;
srom_1(15215) <= 1815445;
srom_1(15216) <= 2187541;
srom_1(15217) <= 2588717;
srom_1(15218) <= 3017090;
srom_1(15219) <= 3470652;
srom_1(15220) <= 3947276;
srom_1(15221) <= 4444726;
srom_1(15222) <= 4960672;
srom_1(15223) <= 5492691;
srom_1(15224) <= 6038291;
srom_1(15225) <= 6594912;
srom_1(15226) <= 7159945;
srom_1(15227) <= 7730739;
srom_1(15228) <= 8304618;
srom_1(15229) <= 8878891;
srom_1(15230) <= 9450865;
srom_1(15231) <= 10017857;
srom_1(15232) <= 10577210;
srom_1(15233) <= 11126299;
srom_1(15234) <= 11662550;
srom_1(15235) <= 12183449;
srom_1(15236) <= 12686552;
srom_1(15237) <= 13169501;
srom_1(15238) <= 13630031;
srom_1(15239) <= 14065981;
srom_1(15240) <= 14475309;
srom_1(15241) <= 14856094;
srom_1(15242) <= 15206550;
srom_1(15243) <= 15525035;
srom_1(15244) <= 15810055;
srom_1(15245) <= 16060273;
srom_1(15246) <= 16274516;
srom_1(15247) <= 16451779;
srom_1(15248) <= 16591232;
srom_1(15249) <= 16692219;
srom_1(15250) <= 16754268;
srom_1(15251) <= 16777087;
srom_1(15252) <= 16760570;
srom_1(15253) <= 16704794;
srom_1(15254) <= 16610020;
srom_1(15255) <= 16476694;
srom_1(15256) <= 16305439;
srom_1(15257) <= 16097060;
srom_1(15258) <= 15852533;
srom_1(15259) <= 15573006;
srom_1(15260) <= 15259788;
srom_1(15261) <= 14914349;
srom_1(15262) <= 14538308;
srom_1(15263) <= 14133430;
srom_1(15264) <= 13701611;
srom_1(15265) <= 13244879;
srom_1(15266) <= 12765374;
srom_1(15267) <= 12265344;
srom_1(15268) <= 11747135;
srom_1(15269) <= 11213177;
srom_1(15270) <= 10665974;
srom_1(15271) <= 10108091;
srom_1(15272) <= 9542145;
srom_1(15273) <= 8970789;
srom_1(15274) <= 8396704;
srom_1(15275) <= 7822580;
srom_1(15276) <= 7251111;
srom_1(15277) <= 6684976;
srom_1(15278) <= 6126830;
srom_1(15279) <= 5579290;
srom_1(15280) <= 5044924;
srom_1(15281) <= 4526237;
srom_1(15282) <= 4025663;
srom_1(15283) <= 3545548;
srom_1(15284) <= 3088143;
srom_1(15285) <= 2655595;
srom_1(15286) <= 2249930;
srom_1(15287) <= 1873052;
srom_1(15288) <= 1526727;
srom_1(15289) <= 1212581;
srom_1(15290) <= 932085;
srom_1(15291) <= 686555;
srom_1(15292) <= 477143;
srom_1(15293) <= 304830;
srom_1(15294) <= 170425;
srom_1(15295) <= 74558;
srom_1(15296) <= 17678;
srom_1(15297) <= 53;
srom_1(15298) <= 21764;
srom_1(15299) <= 82710;
srom_1(15300) <= 182606;
srom_1(15301) <= 320982;
srom_1(15302) <= 497190;
srom_1(15303) <= 710403;
srom_1(15304) <= 959623;
srom_1(15305) <= 1243679;
srom_1(15306) <= 1561241;
srom_1(15307) <= 1910818;
srom_1(15308) <= 2290772;
srom_1(15309) <= 2699321;
srom_1(15310) <= 3134548;
srom_1(15311) <= 3594414;
srom_1(15312) <= 4076762;
srom_1(15313) <= 4579329;
srom_1(15314) <= 5099759;
srom_1(15315) <= 5635612;
srom_1(15316) <= 6184374;
srom_1(15317) <= 6743473;
srom_1(15318) <= 7310286;
srom_1(15319) <= 7882156;
srom_1(15320) <= 8456401;
srom_1(15321) <= 9030328;
srom_1(15322) <= 9601246;
srom_1(15323) <= 10166478;
srom_1(15324) <= 10723372;
srom_1(15325) <= 11269318;
srom_1(15326) <= 11801755;
srom_1(15327) <= 12318186;
srom_1(15328) <= 12816191;
srom_1(15329) <= 13293433;
srom_1(15330) <= 13747675;
srom_1(15331) <= 14176786;
srom_1(15332) <= 14578754;
srom_1(15333) <= 14951695;
srom_1(15334) <= 15293859;
srom_1(15335) <= 15603642;
srom_1(15336) <= 15879591;
srom_1(15337) <= 16120413;
srom_1(15338) <= 16324977;
srom_1(15339) <= 16492325;
srom_1(15340) <= 16621672;
srom_1(15341) <= 16712411;
srom_1(15342) <= 16764117;
srom_1(15343) <= 16776547;
srom_1(15344) <= 16749643;
srom_1(15345) <= 16683532;
srom_1(15346) <= 16578523;
srom_1(15347) <= 16435108;
srom_1(15348) <= 16253961;
srom_1(15349) <= 16035930;
srom_1(15350) <= 15782039;
srom_1(15351) <= 15493477;
srom_1(15352) <= 15171598;
srom_1(15353) <= 14817911;
srom_1(15354) <= 14434075;
srom_1(15355) <= 14021890;
srom_1(15356) <= 13583288;
srom_1(15357) <= 13120326;
srom_1(15358) <= 12635176;
srom_1(15359) <= 12130113;
srom_1(15360) <= 11607504;
srom_1(15361) <= 11069800;
srom_1(15362) <= 10519524;
srom_1(15363) <= 9959255;
srom_1(15364) <= 9391620;
srom_1(15365) <= 8819283;
srom_1(15366) <= 8244925;
srom_1(15367) <= 7671241;
srom_1(15368) <= 7100922;
srom_1(15369) <= 6536640;
srom_1(15370) <= 5981044;
srom_1(15371) <= 5436737;
srom_1(15372) <= 4906272;
srom_1(15373) <= 4392138;
srom_1(15374) <= 3896744;
srom_1(15375) <= 3422414;
srom_1(15376) <= 2971372;
srom_1(15377) <= 2545733;
srom_1(15378) <= 2147494;
srom_1(15379) <= 1778521;
srom_1(15380) <= 1440546;
srom_1(15381) <= 1135152;
srom_1(15382) <= 863772;
srom_1(15383) <= 627679;
srom_1(15384) <= 427979;
srom_1(15385) <= 265610;
srom_1(15386) <= 141332;
srom_1(15387) <= 55728;
srom_1(15388) <= 9200;
srom_1(15389) <= 1966;
srom_1(15390) <= 34060;
srom_1(15391) <= 105331;
srom_1(15392) <= 215445;
srom_1(15393) <= 363886;
srom_1(15394) <= 549958;
srom_1(15395) <= 772787;
srom_1(15396) <= 1031330;
srom_1(15397) <= 1324374;
srom_1(15398) <= 1650545;
srom_1(15399) <= 2008312;
srom_1(15400) <= 2395999;
srom_1(15401) <= 2811787;
srom_1(15402) <= 3253727;
srom_1(15403) <= 3719746;
srom_1(15404) <= 4207659;
srom_1(15405) <= 4715178;
srom_1(15406) <= 5239923;
srom_1(15407) <= 5779433;
srom_1(15408) <= 6331179;
srom_1(15409) <= 6892572;
srom_1(15410) <= 7460981;
srom_1(15411) <= 8033740;
srom_1(15412) <= 8608163;
srom_1(15413) <= 9181556;
srom_1(15414) <= 9751231;
srom_1(15415) <= 10314516;
srom_1(15416) <= 10868770;
srom_1(15417) <= 11411393;
srom_1(15418) <= 11939842;
srom_1(15419) <= 12451637;
srom_1(15420) <= 12944380;
srom_1(15421) <= 13415759;
srom_1(15422) <= 13863564;
srom_1(15423) <= 14285695;
srom_1(15424) <= 14680173;
srom_1(15425) <= 15045147;
srom_1(15426) <= 15378907;
srom_1(15427) <= 15679886;
srom_1(15428) <= 15946675;
srom_1(15429) <= 16178021;
srom_1(15430) <= 16372839;
srom_1(15431) <= 16530217;
srom_1(15432) <= 16649416;
srom_1(15433) <= 16729877;
srom_1(15434) <= 16771224;
srom_1(15435) <= 16773261;
srom_1(15436) <= 16735979;
srom_1(15437) <= 16659554;
srom_1(15438) <= 16544344;
srom_1(15439) <= 16390889;
srom_1(15440) <= 16199908;
srom_1(15441) <= 15972297;
srom_1(15442) <= 15709124;
srom_1(15443) <= 15411622;
srom_1(15444) <= 15081187;
srom_1(15445) <= 14719368;
srom_1(15446) <= 14327863;
srom_1(15447) <= 13908505;
srom_1(15448) <= 13463264;
srom_1(15449) <= 12994225;
srom_1(15450) <= 12503589;
srom_1(15451) <= 11993656;
srom_1(15452) <= 11466818;
srom_1(15453) <= 10925546;
srom_1(15454) <= 10372377;
srom_1(15455) <= 9809905;
srom_1(15456) <= 9240768;
srom_1(15457) <= 8667635;
srom_1(15458) <= 8093194;
srom_1(15459) <= 7520138;
srom_1(15460) <= 6951154;
srom_1(15461) <= 6388912;
srom_1(15462) <= 5836046;
srom_1(15463) <= 5295150;
srom_1(15464) <= 4768761;
srom_1(15465) <= 4259346;
srom_1(15466) <= 3769295;
srom_1(15467) <= 3300905;
srom_1(15468) <= 2856374;
srom_1(15469) <= 2437785;
srom_1(15470) <= 2047101;
srom_1(15471) <= 1686155;
srom_1(15472) <= 1356639;
srom_1(15473) <= 1060098;
srom_1(15474) <= 797923;
srom_1(15475) <= 571344;
srom_1(15476) <= 381422;
srom_1(15477) <= 229049;
srom_1(15478) <= 114938;
srom_1(15479) <= 39626;
srom_1(15480) <= 3465;
srom_1(15481) <= 6625;
srom_1(15482) <= 49091;
srom_1(15483) <= 130663;
srom_1(15484) <= 250960;
srom_1(15485) <= 409417;
srom_1(15486) <= 605292;
srom_1(15487) <= 837665;
srom_1(15488) <= 1105447;
srom_1(15489) <= 1407382;
srom_1(15490) <= 1742055;
srom_1(15491) <= 2107895;
srom_1(15492) <= 2503188;
srom_1(15493) <= 2926080;
srom_1(15494) <= 3374587;
srom_1(15495) <= 3846607;
srom_1(15496) <= 4339926;
srom_1(15497) <= 4852230;
srom_1(15498) <= 5381118;
srom_1(15499) <= 5924109;
srom_1(15500) <= 6478657;
srom_1(15501) <= 7042161;
srom_1(15502) <= 7611979;
srom_1(15503) <= 8185439;
srom_1(15504) <= 8759852;
srom_1(15505) <= 9332524;
srom_1(15506) <= 9900769;
srom_1(15507) <= 10461923;
srom_1(15508) <= 11013355;
srom_1(15509) <= 11552479;
srom_1(15510) <= 12076766;
srom_1(15511) <= 12583758;
srom_1(15512) <= 13071078;
srom_1(15513) <= 13536440;
srom_1(15514) <= 13977661;
srom_1(15515) <= 14392674;
srom_1(15516) <= 14779532;
srom_1(15517) <= 15136420;
srom_1(15518) <= 15461666;
srom_1(15519) <= 15753744;
srom_1(15520) <= 16011284;
srom_1(15521) <= 16233078;
srom_1(15522) <= 16418088;
srom_1(15523) <= 16565444;
srom_1(15524) <= 16674456;
srom_1(15525) <= 16744613;
srom_1(15526) <= 16775586;
srom_1(15527) <= 16767229;
srom_1(15528) <= 16719583;
srom_1(15529) <= 16632869;
srom_1(15530) <= 16507495;
srom_1(15531) <= 16344049;
srom_1(15532) <= 16143297;
srom_1(15533) <= 15906181;
srom_1(15534) <= 15633812;
srom_1(15535) <= 15327468;
srom_1(15536) <= 14988585;
srom_1(15537) <= 14618753;
srom_1(15538) <= 14219706;
srom_1(15539) <= 13793314;
srom_1(15540) <= 13341578;
srom_1(15541) <= 12866615;
srom_1(15542) <= 12370654;
srom_1(15543) <= 11856020;
srom_1(15544) <= 11325125;
srom_1(15545) <= 10780461;
srom_1(15546) <= 10224580;
srom_1(15547) <= 9660089;
srom_1(15548) <= 9089636;
srom_1(15549) <= 8515896;
srom_1(15550) <= 7941559;
srom_1(15551) <= 7369318;
srom_1(15552) <= 6801857;
srom_1(15553) <= 6241837;
srom_1(15554) <= 5691884;
srom_1(15555) <= 5154577;
srom_1(15556) <= 4632435;
srom_1(15557) <= 4127907;
srom_1(15558) <= 3643359;
srom_1(15559) <= 3181063;
srom_1(15560) <= 2743187;
srom_1(15561) <= 2331784;
srom_1(15562) <= 1948784;
srom_1(15563) <= 1595983;
srom_1(15564) <= 1275034;
srom_1(15565) <= 987443;
srom_1(15566) <= 734559;
srom_1(15567) <= 517568;
srom_1(15568) <= 337486;
srom_1(15569) <= 195159;
srom_1(15570) <= 91254;
srom_1(15571) <= 26258;
srom_1(15572) <= 475;
srom_1(15573) <= 14028;
srom_1(15574) <= 66852;
srom_1(15575) <= 158699;
srom_1(15576) <= 289140;
srom_1(15577) <= 457561;
srom_1(15578) <= 663174;
srom_1(15579) <= 905014;
srom_1(15580) <= 1181948;
srom_1(15581) <= 1492675;
srom_1(15582) <= 1835741;
srom_1(15583) <= 2209534;
srom_1(15584) <= 2612304;
srom_1(15585) <= 3042161;
srom_1(15586) <= 3497089;
srom_1(15587) <= 3974955;
srom_1(15588) <= 4473518;
srom_1(15589) <= 4990440;
srom_1(15590) <= 5523298;
srom_1(15591) <= 6069591;
srom_1(15592) <= 6626760;
srom_1(15593) <= 7192191;
srom_1(15594) <= 7763231;
srom_1(15595) <= 8337205;
srom_1(15596) <= 8911419;
srom_1(15597) <= 9483182;
srom_1(15598) <= 10049812;
srom_1(15599) <= 10608652;
srom_1(15600) <= 11157082;
srom_1(15601) <= 11692529;
srom_1(15602) <= 12212483;
srom_1(15603) <= 12714505;
srom_1(15604) <= 13196242;
srom_1(15605) <= 13655434;
srom_1(15606) <= 14089929;
srom_1(15607) <= 14497687;
srom_1(15608) <= 14876799;
srom_1(15609) <= 15225484;
srom_1(15610) <= 15542110;
srom_1(15611) <= 15825190;
srom_1(15612) <= 16073397;
srom_1(15613) <= 16285568;
srom_1(15614) <= 16460707;
srom_1(15615) <= 16597994;
srom_1(15616) <= 16696783;
srom_1(15617) <= 16756613;
srom_1(15618) <= 16777203;
srom_1(15619) <= 16758455;
srom_1(15620) <= 16700458;
srom_1(15621) <= 16603485;
srom_1(15622) <= 16467988;
srom_1(15623) <= 16294605;
srom_1(15624) <= 16084148;
srom_1(15625) <= 15837604;
srom_1(15626) <= 15556129;
srom_1(15627) <= 15241042;
srom_1(15628) <= 14893823;
srom_1(15629) <= 14516098;
srom_1(15630) <= 14109640;
srom_1(15631) <= 13676353;
srom_1(15632) <= 13218271;
srom_1(15633) <= 12737540;
srom_1(15634) <= 12236416;
srom_1(15635) <= 11717248;
srom_1(15636) <= 11182471;
srom_1(15637) <= 10634593;
srom_1(15638) <= 10076182;
srom_1(15639) <= 9509858;
srom_1(15640) <= 8938276;
srom_1(15641) <= 8364116;
srom_1(15642) <= 7790071;
srom_1(15643) <= 7218833;
srom_1(15644) <= 6653080;
srom_1(15645) <= 6095466;
srom_1(15646) <= 5548605;
srom_1(15647) <= 5015062;
srom_1(15648) <= 4497338;
srom_1(15649) <= 3997862;
srom_1(15650) <= 3518976;
srom_1(15651) <= 3062925;
srom_1(15652) <= 2631848;
srom_1(15653) <= 2227767;
srom_1(15654) <= 1852576;
srom_1(15655) <= 1508034;
srom_1(15656) <= 1195758;
srom_1(15657) <= 917212;
srom_1(15658) <= 673701;
srom_1(15659) <= 466369;
srom_1(15660) <= 296186;
srom_1(15661) <= 163952;
srom_1(15662) <= 70285;
srom_1(15663) <= 15627;
srom_1(15664) <= 232;
srom_1(15665) <= 24173;
srom_1(15666) <= 87338;
srom_1(15667) <= 189430;
srom_1(15668) <= 329971;
srom_1(15669) <= 508302;
srom_1(15670) <= 723586;
srom_1(15671) <= 974814;
srom_1(15672) <= 1260808;
srom_1(15673) <= 1580227;
srom_1(15674) <= 1931572;
srom_1(15675) <= 2313197;
srom_1(15676) <= 2723311;
srom_1(15677) <= 3159992;
srom_1(15678) <= 3621192;
srom_1(15679) <= 4104747;
srom_1(15680) <= 4608392;
srom_1(15681) <= 5129762;
srom_1(15682) <= 5666415;
srom_1(15683) <= 6215833;
srom_1(15684) <= 6775440;
srom_1(15685) <= 7342612;
srom_1(15686) <= 7914689;
srom_1(15687) <= 8488988;
srom_1(15688) <= 9062816;
srom_1(15689) <= 9633483;
srom_1(15690) <= 10198312;
srom_1(15691) <= 10754654;
srom_1(15692) <= 11299902;
srom_1(15693) <= 11831497;
srom_1(15694) <= 12346948;
srom_1(15695) <= 12843836;
srom_1(15696) <= 13319833;
srom_1(15697) <= 13772705;
srom_1(15698) <= 14200329;
srom_1(15699) <= 14600701;
srom_1(15700) <= 14971941;
srom_1(15701) <= 15312310;
srom_1(15702) <= 15620211;
srom_1(15703) <= 15894201;
srom_1(15704) <= 16132995;
srom_1(15705) <= 16335472;
srom_1(15706) <= 16500684;
srom_1(15707) <= 16627856;
srom_1(15708) <= 16716391;
srom_1(15709) <= 16765874;
srom_1(15710) <= 16776073;
srom_1(15711) <= 16746940;
srom_1(15712) <= 16678613;
srom_1(15713) <= 16571410;
srom_1(15714) <= 16425836;
srom_1(15715) <= 16242573;
srom_1(15716) <= 16022479;
srom_1(15717) <= 15766588;
srom_1(15718) <= 15476098;
srom_1(15719) <= 15152373;
srom_1(15720) <= 14796931;
srom_1(15721) <= 14411437;
srom_1(15722) <= 13997701;
srom_1(15723) <= 13557661;
srom_1(15724) <= 13093382;
srom_1(15725) <= 12607041;
srom_1(15726) <= 12100918;
srom_1(15727) <= 11577386;
srom_1(15728) <= 11038902;
srom_1(15729) <= 10487989;
srom_1(15730) <= 9927232;
srom_1(15731) <= 9359259;
srom_1(15732) <= 8786735;
srom_1(15733) <= 8212343;
srom_1(15734) <= 7638779;
srom_1(15735) <= 7068730;
srom_1(15736) <= 6504871;
srom_1(15737) <= 5949845;
srom_1(15738) <= 5406256;
srom_1(15739) <= 4876651;
srom_1(15740) <= 4363516;
srom_1(15741) <= 3869255;
srom_1(15742) <= 3396188;
srom_1(15743) <= 2946531;
srom_1(15744) <= 2522395;
srom_1(15745) <= 2125767;
srom_1(15746) <= 1758507;
srom_1(15747) <= 1422338;
srom_1(15748) <= 1118837;
srom_1(15749) <= 849426;
srom_1(15750) <= 615369;
srom_1(15751) <= 417763;
srom_1(15752) <= 257535;
srom_1(15753) <= 135437;
srom_1(15754) <= 52041;
srom_1(15755) <= 7737;
srom_1(15756) <= 2735;
srom_1(15757) <= 37056;
srom_1(15758) <= 110541;
srom_1(15759) <= 222845;
srom_1(15760) <= 373440;
srom_1(15761) <= 561622;
srom_1(15762) <= 786507;
srom_1(15763) <= 1047041;
srom_1(15764) <= 1342002;
srom_1(15765) <= 1670007;
srom_1(15766) <= 2029517;
srom_1(15767) <= 2418848;
srom_1(15768) <= 2836173;
srom_1(15769) <= 3279535;
srom_1(15770) <= 3746855;
srom_1(15771) <= 4235943;
srom_1(15772) <= 4744503;
srom_1(15773) <= 5270152;
srom_1(15774) <= 5810424;
srom_1(15775) <= 6362787;
srom_1(15776) <= 6924649;
srom_1(15777) <= 7493376;
srom_1(15778) <= 8066301;
srom_1(15779) <= 8640737;
srom_1(15780) <= 9213992;
srom_1(15781) <= 9783375;
srom_1(15782) <= 10346219;
srom_1(15783) <= 10899882;
srom_1(15784) <= 11441769;
srom_1(15785) <= 11969338;
srom_1(15786) <= 12480117;
srom_1(15787) <= 12971709;
srom_1(15788) <= 13441809;
srom_1(15789) <= 13888213;
srom_1(15790) <= 14308827;
srom_1(15791) <= 14701680;
srom_1(15792) <= 15064928;
srom_1(15793) <= 15396869;
srom_1(15794) <= 15695945;
srom_1(15795) <= 15960755;
srom_1(15796) <= 16190057;
srom_1(15797) <= 16382775;
srom_1(15798) <= 16538005;
srom_1(15799) <= 16655020;
srom_1(15800) <= 16733272;
srom_1(15801) <= 16772392;
srom_1(15802) <= 16772197;
srom_1(15803) <= 16732689;
srom_1(15804) <= 16654053;
srom_1(15805) <= 16536657;
srom_1(15806) <= 16381053;
srom_1(15807) <= 16187969;
srom_1(15808) <= 15958311;
srom_1(15809) <= 15693156;
srom_1(15810) <= 15393748;
srom_1(15811) <= 15061490;
srom_1(15812) <= 14697940;
srom_1(15813) <= 14304804;
srom_1(15814) <= 13883925;
srom_1(15815) <= 13437277;
srom_1(15816) <= 12966953;
srom_1(15817) <= 12475160;
srom_1(15818) <= 11964204;
srom_1(15819) <= 11436481;
srom_1(15820) <= 10894465;
srom_1(15821) <= 10340698;
srom_1(15822) <= 9777777;
srom_1(15823) <= 9208342;
srom_1(15824) <= 8635063;
srom_1(15825) <= 8060628;
srom_1(15826) <= 7487732;
srom_1(15827) <= 6919059;
srom_1(15828) <= 6357278;
srom_1(15829) <= 5805023;
srom_1(15830) <= 5264883;
srom_1(15831) <= 4739391;
srom_1(15832) <= 4231011;
srom_1(15833) <= 3742128;
srom_1(15834) <= 3275034;
srom_1(15835) <= 2831919;
srom_1(15836) <= 2414861;
srom_1(15837) <= 2025817;
srom_1(15838) <= 1666609;
srom_1(15839) <= 1338923;
srom_1(15840) <= 1044296;
srom_1(15841) <= 784109;
srom_1(15842) <= 559582;
srom_1(15843) <= 371767;
srom_1(15844) <= 221547;
srom_1(15845) <= 109625;
srom_1(15846) <= 36525;
srom_1(15847) <= 2592;
srom_1(15848) <= 7983;
srom_1(15849) <= 52674;
srom_1(15850) <= 136455;
srom_1(15851) <= 258933;
srom_1(15852) <= 419534;
srom_1(15853) <= 617505;
srom_1(15854) <= 851917;
srom_1(15855) <= 1121671;
srom_1(15856) <= 1425503;
srom_1(15857) <= 1761986;
srom_1(15858) <= 2129545;
srom_1(15859) <= 2526454;
srom_1(15860) <= 2950852;
srom_1(15861) <= 3400751;
srom_1(15862) <= 3874039;
srom_1(15863) <= 4368497;
srom_1(15864) <= 4881807;
srom_1(15865) <= 5411562;
srom_1(15866) <= 5955277;
srom_1(15867) <= 6510403;
srom_1(15868) <= 7074336;
srom_1(15869) <= 7644433;
srom_1(15870) <= 8218019;
srom_1(15871) <= 8792405;
srom_1(15872) <= 9364897;
srom_1(15873) <= 9932812;
srom_1(15874) <= 10493485;
srom_1(15875) <= 11044287;
srom_1(15876) <= 11582636;
srom_1(15877) <= 12106007;
srom_1(15878) <= 12611946;
srom_1(15879) <= 13098081;
srom_1(15880) <= 13562131;
srom_1(15881) <= 14001920;
srom_1(15882) <= 14415387;
srom_1(15883) <= 14800592;
srom_1(15884) <= 15155729;
srom_1(15885) <= 15479133;
srom_1(15886) <= 15769287;
srom_1(15887) <= 16024830;
srom_1(15888) <= 16244565;
srom_1(15889) <= 16427460;
srom_1(15890) <= 16572658;
srom_1(15891) <= 16679479;
srom_1(15892) <= 16747420;
srom_1(15893) <= 16776165;
srom_1(15894) <= 16765577;
srom_1(15895) <= 16715706;
srom_1(15896) <= 16626788;
srom_1(15897) <= 16499237;
srom_1(15898) <= 16333653;
srom_1(15899) <= 16130811;
srom_1(15900) <= 15891664;
srom_1(15901) <= 15617333;
srom_1(15902) <= 15309103;
srom_1(15903) <= 14968421;
srom_1(15904) <= 14596884;
srom_1(15905) <= 14196234;
srom_1(15906) <= 13768351;
srom_1(15907) <= 13315239;
srom_1(15908) <= 12839026;
srom_1(15909) <= 12341942;
srom_1(15910) <= 11826320;
srom_1(15911) <= 11294577;
srom_1(15912) <= 10749208;
srom_1(15913) <= 10192768;
srom_1(15914) <= 9627869;
srom_1(15915) <= 9057157;
srom_1(15916) <= 8483311;
srom_1(15917) <= 7909021;
srom_1(15918) <= 7336980;
srom_1(15919) <= 6769870;
srom_1(15920) <= 6210351;
srom_1(15921) <= 5661046;
srom_1(15922) <= 5124532;
srom_1(15923) <= 4603325;
srom_1(15924) <= 4099868;
srom_1(15925) <= 3616522;
srom_1(15926) <= 3155554;
srom_1(15927) <= 2719126;
srom_1(15928) <= 2309284;
srom_1(15929) <= 1927950;
srom_1(15930) <= 1576912;
srom_1(15931) <= 1257816;
srom_1(15932) <= 972160;
srom_1(15933) <= 721281;
srom_1(15934) <= 506357;
srom_1(15935) <= 328396;
srom_1(15936) <= 188232;
srom_1(15937) <= 86523;
srom_1(15938) <= 23744;
srom_1(15939) <= 192;
srom_1(15940) <= 15975;
srom_1(15941) <= 71021;
srom_1(15942) <= 165070;
srom_1(15943) <= 297683;
srom_1(15944) <= 468237;
srom_1(15945) <= 675932;
srom_1(15946) <= 919794;
srom_1(15947) <= 1198681;
srom_1(15948) <= 1511283;
srom_1(15949) <= 1856135;
srom_1(15950) <= 2231621;
srom_1(15951) <= 2635979;
srom_1(15952) <= 3067312;
srom_1(15953) <= 3523600;
srom_1(15954) <= 4002700;
srom_1(15955) <= 4502368;
srom_1(15956) <= 5020260;
srom_1(15957) <= 5553947;
srom_1(15958) <= 6100927;
srom_1(15959) <= 6658634;
srom_1(15960) <= 7224454;
srom_1(15961) <= 7795733;
srom_1(15962) <= 8369792;
srom_1(15963) <= 8943940;
srom_1(15964) <= 9515483;
srom_1(15965) <= 10081742;
srom_1(15966) <= 10640061;
srom_1(15967) <= 11187823;
srom_1(15968) <= 11722458;
srom_1(15969) <= 12241459;
srom_1(15970) <= 12742393;
srom_1(15971) <= 13222911;
srom_1(15972) <= 13680759;
srom_1(15973) <= 14113790;
srom_1(15974) <= 14519974;
srom_1(15975) <= 14897406;
srom_1(15976) <= 15244315;
srom_1(15977) <= 15559076;
srom_1(15978) <= 15840212;
srom_1(15979) <= 16086405;
srom_1(15980) <= 16296501;
srom_1(15981) <= 16469514;
srom_1(15982) <= 16604632;
srom_1(15983) <= 16701223;
srom_1(15984) <= 16758833;
srom_1(15985) <= 16777192;
srom_1(15986) <= 16756214;
srom_1(15987) <= 16695997;
srom_1(15988) <= 16596825;
srom_1(15989) <= 16459161;
srom_1(15990) <= 16283651;
srom_1(15991) <= 16071119;
srom_1(15992) <= 15822562;
srom_1(15993) <= 15539143;
srom_1(15994) <= 15222194;
srom_1(15995) <= 14873199;
srom_1(15996) <= 14493796;
srom_1(15997) <= 14085763;
srom_1(15998) <= 13651015;
srom_1(15999) <= 13191589;
srom_1(16000) <= 12709641;
srom_1(16001) <= 12207429;
srom_1(16002) <= 11687310;
srom_1(16003) <= 11151723;
srom_1(16004) <= 10603178;
srom_1(16005) <= 10044248;
srom_1(16006) <= 9477554;
srom_1(16007) <= 8905754;
srom_1(16008) <= 8331528;
srom_1(16009) <= 7757571;
srom_1(16010) <= 7186572;
srom_1(16011) <= 6621210;
srom_1(16012) <= 6064137;
srom_1(16013) <= 5517963;
srom_1(16014) <= 4985251;
srom_1(16015) <= 4468498;
srom_1(16016) <= 3970128;
srom_1(16017) <= 3492478;
srom_1(16018) <= 3037788;
srom_1(16019) <= 2608189;
srom_1(16020) <= 2205697;
srom_1(16021) <= 1832198;
srom_1(16022) <= 1489445;
srom_1(16023) <= 1179044;
srom_1(16024) <= 902451;
srom_1(16025) <= 660964;
srom_1(16026) <= 455714;
srom_1(16027) <= 287664;
srom_1(16028) <= 157602;
srom_1(16029) <= 66139;
srom_1(16030) <= 13702;
srom_1(16031) <= 538;
srom_1(16032) <= 26708;
srom_1(16033) <= 92091;
srom_1(16034) <= 196378;
srom_1(16035) <= 339082;
srom_1(16036) <= 519532;
srom_1(16037) <= 736884;
srom_1(16038) <= 990117;
srom_1(16039) <= 1278044;
srom_1(16040) <= 1599315;
srom_1(16041) <= 1952423;
srom_1(16042) <= 2335713;
srom_1(16043) <= 2747387;
srom_1(16044) <= 3185514;
srom_1(16045) <= 3648041;
srom_1(16046) <= 4132798;
srom_1(16047) <= 4637511;
srom_1(16048) <= 5159815;
srom_1(16049) <= 5697260;
srom_1(16050) <= 6247325;
srom_1(16051) <= 6807432;
srom_1(16052) <= 7374953;
srom_1(16053) <= 7947228;
srom_1(16054) <= 8521572;
srom_1(16055) <= 9095293;
srom_1(16056) <= 9665700;
srom_1(16057) <= 10230118;
srom_1(16058) <= 10785901;
srom_1(16059) <= 11330442;
srom_1(16060) <= 11861188;
srom_1(16061) <= 12375650;
srom_1(16062) <= 12871415;
srom_1(16063) <= 13346158;
srom_1(16064) <= 13797654;
srom_1(16065) <= 14223785;
srom_1(16066) <= 14622553;
srom_1(16067) <= 14992088;
srom_1(16068) <= 15330657;
srom_1(16069) <= 15636672;
srom_1(16070) <= 15908698;
srom_1(16071) <= 16145460;
srom_1(16072) <= 16345848;
srom_1(16073) <= 16508921;
srom_1(16074) <= 16633916;
srom_1(16075) <= 16720245;
srom_1(16076) <= 16767504;
srom_1(16077) <= 16775472;
srom_1(16078) <= 16744111;
srom_1(16079) <= 16673568;
srom_1(16080) <= 16564175;
srom_1(16081) <= 16416443;
srom_1(16082) <= 16231065;
srom_1(16083) <= 16008912;
srom_1(16084) <= 15751025;
srom_1(16085) <= 15458613;
srom_1(16086) <= 15133047;
srom_1(16087) <= 14775854;
srom_1(16088) <= 14388708;
srom_1(16089) <= 13973427;
srom_1(16090) <= 13531956;
srom_1(16091) <= 13066367;
srom_1(16092) <= 12578841;
srom_1(16093) <= 12071667;
srom_1(16094) <= 11547221;
srom_1(16095) <= 11007963;
srom_1(16096) <= 10456422;
srom_1(16097) <= 9895185;
srom_1(16098) <= 9326883;
srom_1(16099) <= 8754181;
srom_1(16100) <= 8179764;
srom_1(16101) <= 7606327;
srom_1(16102) <= 7036558;
srom_1(16103) <= 6473130;
srom_1(16104) <= 5918683;
srom_1(16105) <= 5375819;
srom_1(16106) <= 4847083;
srom_1(16107) <= 4334955;
srom_1(16108) <= 3841835;
srom_1(16109) <= 3370037;
srom_1(16110) <= 2921773;
srom_1(16111) <= 2499144;
srom_1(16112) <= 2104134;
srom_1(16113) <= 1738593;
srom_1(16114) <= 1404236;
srom_1(16115) <= 1102632;
srom_1(16116) <= 835194;
srom_1(16117) <= 603176;
srom_1(16118) <= 407668;
srom_1(16119) <= 249584;
srom_1(16120) <= 129667;
srom_1(16121) <= 48479;
srom_1(16122) <= 6401;
srom_1(16123) <= 3630;
srom_1(16124) <= 40179;
srom_1(16125) <= 115877;
srom_1(16126) <= 230368;
srom_1(16127) <= 383116;
srom_1(16128) <= 573404;
srom_1(16129) <= 800341;
srom_1(16130) <= 1062862;
srom_1(16131) <= 1359735;
srom_1(16132) <= 1689570;
srom_1(16133) <= 2050818;
srom_1(16134) <= 2441787;
srom_1(16135) <= 2860642;
srom_1(16136) <= 3305420;
srom_1(16137) <= 3774035;
srom_1(16138) <= 4264288;
srom_1(16139) <= 4773883;
srom_1(16140) <= 5300428;
srom_1(16141) <= 5841454;
srom_1(16142) <= 6394425;
srom_1(16143) <= 6956747;
srom_1(16144) <= 7525784;
srom_1(16145) <= 8098867;
srom_1(16146) <= 8673309;
srom_1(16147) <= 9246415;
srom_1(16148) <= 9815499;
srom_1(16149) <= 10377892;
srom_1(16150) <= 10930956;
srom_1(16151) <= 11472098;
srom_1(16152) <= 11998781;
srom_1(16153) <= 12508535;
srom_1(16154) <= 12998968;
srom_1(16155) <= 13467782;
srom_1(16156) <= 13912779;
srom_1(16157) <= 14331870;
srom_1(16158) <= 14723091;
srom_1(16159) <= 15084608;
srom_1(16160) <= 15414725;
srom_1(16161) <= 15711894;
srom_1(16162) <= 15974722;
srom_1(16163) <= 16201976;
srom_1(16164) <= 16392590;
srom_1(16165) <= 16545671;
srom_1(16166) <= 16660500;
srom_1(16167) <= 16736540;
srom_1(16168) <= 16773433;
srom_1(16169) <= 16771007;
srom_1(16170) <= 16729273;
srom_1(16171) <= 16648427;
srom_1(16172) <= 16528848;
srom_1(16173) <= 16371096;
srom_1(16174) <= 16175912;
srom_1(16175) <= 15944210;
srom_1(16176) <= 15677078;
srom_1(16177) <= 15375767;
srom_1(16178) <= 15041691;
srom_1(16179) <= 14676417;
srom_1(16180) <= 14281657;
srom_1(16181) <= 13859262;
srom_1(16182) <= 13411214;
srom_1(16183) <= 12939613;
srom_1(16184) <= 12446670;
srom_1(16185) <= 11934698;
srom_1(16186) <= 11406097;
srom_1(16187) <= 10863346;
srom_1(16188) <= 10308990;
srom_1(16189) <= 9745629;
srom_1(16190) <= 9175904;
srom_1(16191) <= 8602488;
srom_1(16192) <= 8028068;
srom_1(16193) <= 7455339;
srom_1(16194) <= 6886987;
srom_1(16195) <= 6325676;
srom_1(16196) <= 5774039;
srom_1(16197) <= 5234662;
srom_1(16198) <= 4710076;
srom_1(16199) <= 4202739;
srom_1(16200) <= 3715031;
srom_1(16201) <= 3249239;
srom_1(16202) <= 2807548;
srom_1(16203) <= 2392028;
srom_1(16204) <= 2004628;
srom_1(16205) <= 1647165;
srom_1(16206) <= 1321315;
srom_1(16207) <= 1028605;
srom_1(16208) <= 770409;
srom_1(16209) <= 547938;
srom_1(16210) <= 362234;
srom_1(16211) <= 214169;
srom_1(16212) <= 104436;
srom_1(16213) <= 33551;
srom_1(16214) <= 1845;
srom_1(16215) <= 9468;
srom_1(16216) <= 56383;
srom_1(16217) <= 142371;
srom_1(16218) <= 267029;
srom_1(16219) <= 429771;
srom_1(16220) <= 629835;
srom_1(16221) <= 866283;
srom_1(16222) <= 1138005;
srom_1(16223) <= 1443728;
srom_1(16224) <= 1782018;
srom_1(16225) <= 2151288;
srom_1(16226) <= 2549808;
srom_1(16227) <= 2975707;
srom_1(16228) <= 3426990;
srom_1(16229) <= 3901539;
srom_1(16230) <= 4397129;
srom_1(16231) <= 4911437;
srom_1(16232) <= 5442051;
srom_1(16233) <= 5986482;
srom_1(16234) <= 6542178;
srom_1(16235) <= 7106531;
srom_1(16236) <= 7676898;
srom_1(16237) <= 8250601;
srom_1(16238) <= 8824952;
srom_1(16239) <= 9397256;
srom_1(16240) <= 9964831;
srom_1(16241) <= 10525014;
srom_1(16242) <= 11075179;
srom_1(16243) <= 11612745;
srom_1(16244) <= 12135193;
srom_1(16245) <= 12640071;
srom_1(16246) <= 13125013;
srom_1(16247) <= 13587744;
srom_1(16248) <= 14026095;
srom_1(16249) <= 14438009;
srom_1(16250) <= 14821556;
srom_1(16251) <= 15174936;
srom_1(16252) <= 15496493;
srom_1(16253) <= 15784719;
srom_1(16254) <= 16038262;
srom_1(16255) <= 16255933;
srom_1(16256) <= 16436711;
srom_1(16257) <= 16579749;
srom_1(16258) <= 16684376;
srom_1(16259) <= 16750101;
srom_1(16260) <= 16776617;
srom_1(16261) <= 16763798;
srom_1(16262) <= 16711705;
srom_1(16263) <= 16620582;
srom_1(16264) <= 16490856;
srom_1(16265) <= 16323136;
srom_1(16266) <= 16118209;
srom_1(16267) <= 15877035;
srom_1(16268) <= 15600745;
srom_1(16269) <= 15290634;
srom_1(16270) <= 14948158;
srom_1(16271) <= 14574922;
srom_1(16272) <= 14172676;
srom_1(16273) <= 13743306;
srom_1(16274) <= 13288827;
srom_1(16275) <= 12811368;
srom_1(16276) <= 12313170;
srom_1(16277) <= 11796568;
srom_1(16278) <= 11263986;
srom_1(16279) <= 10717919;
srom_1(16280) <= 10160930;
srom_1(16281) <= 9595629;
srom_1(16282) <= 9024668;
srom_1(16283) <= 8450725;
srom_1(16284) <= 7876490;
srom_1(16285) <= 7304657;
srom_1(16286) <= 6737907;
srom_1(16287) <= 6178897;
srom_1(16288) <= 5630250;
srom_1(16289) <= 5094538;
srom_1(16290) <= 4574272;
srom_1(16291) <= 4071893;
srom_1(16292) <= 3589757;
srom_1(16293) <= 3130124;
srom_1(16294) <= 2695150;
srom_1(16295) <= 2286875;
srom_1(16296) <= 1907213;
srom_1(16297) <= 1557944;
srom_1(16298) <= 1240707;
srom_1(16299) <= 956988;
srom_1(16300) <= 708119;
srom_1(16301) <= 495266;
srom_1(16302) <= 319428;
srom_1(16303) <= 181429;
srom_1(16304) <= 81917;
srom_1(16305) <= 21357;
srom_1(16306) <= 34;
srom_1(16307) <= 18048;
srom_1(16308) <= 75315;
srom_1(16309) <= 171565;
srom_1(16310) <= 306348;
srom_1(16311) <= 479032;
srom_1(16312) <= 688806;
srom_1(16313) <= 934687;
srom_1(16314) <= 1215522;
srom_1(16315) <= 1529994;
srom_1(16316) <= 1876629;
srom_1(16317) <= 2253800;
srom_1(16318) <= 2659740;
srom_1(16319) <= 3092544;
srom_1(16320) <= 3550184;
srom_1(16321) <= 4030512;
srom_1(16322) <= 4531277;
srom_1(16323) <= 5050131;
srom_1(16324) <= 5584639;
srom_1(16325) <= 6132297;
srom_1(16326) <= 6690535;
srom_1(16327) <= 7256735;
srom_1(16328) <= 7828244;
srom_1(16329) <= 8402380;
srom_1(16330) <= 8976452;
srom_1(16331) <= 9547767;
srom_1(16332) <= 10113646;
srom_1(16333) <= 10671436;
srom_1(16334) <= 11218522;
srom_1(16335) <= 11752336;
srom_1(16336) <= 12270377;
srom_1(16337) <= 12770215;
srom_1(16338) <= 13249506;
srom_1(16339) <= 13706003;
srom_1(16340) <= 14137565;
srom_1(16341) <= 14542168;
srom_1(16342) <= 14917914;
srom_1(16343) <= 15263043;
srom_1(16344) <= 15575935;
srom_1(16345) <= 15855123;
srom_1(16346) <= 16099297;
srom_1(16347) <= 16307314;
srom_1(16348) <= 16478198;
srom_1(16349) <= 16611146;
srom_1(16350) <= 16705536;
srom_1(16351) <= 16760926;
srom_1(16352) <= 16777054;
srom_1(16353) <= 16753846;
srom_1(16354) <= 16691411;
srom_1(16355) <= 16590041;
srom_1(16356) <= 16450212;
srom_1(16357) <= 16272579;
srom_1(16358) <= 16057975;
srom_1(16359) <= 15807407;
srom_1(16360) <= 15522050;
srom_1(16361) <= 15203242;
srom_1(16362) <= 14852477;
srom_1(16363) <= 14471401;
srom_1(16364) <= 14061801;
srom_1(16365) <= 13625597;
srom_1(16366) <= 13164836;
srom_1(16367) <= 12681676;
srom_1(16368) <= 12178386;
srom_1(16369) <= 11657323;
srom_1(16370) <= 11120933;
srom_1(16371) <= 10571729;
srom_1(16372) <= 10012288;
srom_1(16373) <= 9445234;
srom_1(16374) <= 8873224;
srom_1(16375) <= 8298942;
srom_1(16376) <= 7725080;
srom_1(16377) <= 7154330;
srom_1(16378) <= 6589368;
srom_1(16379) <= 6032842;
srom_1(16380) <= 5487364;
srom_1(16381) <= 4955491;
srom_1(16382) <= 4439717;
srom_1(16383) <= 3942461;
srom_1(16384) <= 3466054;
srom_1(16385) <= 3012731;
srom_1(16386) <= 2584617;
srom_1(16387) <= 2183720;
srom_1(16388) <= 1811919;
srom_1(16389) <= 1470959;
srom_1(16390) <= 1162439;
srom_1(16391) <= 887804;
srom_1(16392) <= 648343;
srom_1(16393) <= 445179;
srom_1(16394) <= 279264;
srom_1(16395) <= 151377;
srom_1(16396) <= 62117;
srom_1(16397) <= 11903;
srom_1(16398) <= 970;
srom_1(16399) <= 29370;
srom_1(16400) <= 96969;
srom_1(16401) <= 203450;
srom_1(16402) <= 348314;
srom_1(16403) <= 530882;
srom_1(16404) <= 750298;
srom_1(16405) <= 1005532;
srom_1(16406) <= 1295388;
srom_1(16407) <= 1618506;
srom_1(16408) <= 1973372;
srom_1(16409) <= 2358321;
srom_1(16410) <= 2771548;
srom_1(16411) <= 3211116;
srom_1(16412) <= 3674962;
srom_1(16413) <= 4160912;
srom_1(16414) <= 4666688;
srom_1(16415) <= 5189917;
srom_1(16416) <= 5728145;
srom_1(16417) <= 6278850;
srom_1(16418) <= 6839447;
srom_1(16419) <= 7407310;
srom_1(16420) <= 7979774;
srom_1(16421) <= 8554155;
srom_1(16422) <= 9127760;
srom_1(16423) <= 9697898;
srom_1(16424) <= 10261897;
srom_1(16425) <= 10817112;
srom_1(16426) <= 11360938;
srom_1(16427) <= 11890826;
srom_1(16428) <= 12404291;
srom_1(16429) <= 12898925;
srom_1(16430) <= 13372409;
srom_1(16431) <= 13822522;
srom_1(16432) <= 14247153;
srom_1(16433) <= 14644311;
srom_1(16434) <= 15012135;
srom_1(16435) <= 15348898;
srom_1(16436) <= 15653023;
srom_1(16437) <= 15923082;
srom_1(16438) <= 16157809;
srom_1(16439) <= 16356103;
srom_1(16440) <= 16517036;
srom_1(16441) <= 16639851;
srom_1(16442) <= 16723974;
srom_1(16443) <= 16769009;
srom_1(16444) <= 16774745;
srom_1(16445) <= 16741156;
srom_1(16446) <= 16668399;
srom_1(16447) <= 16556815;
srom_1(16448) <= 16406928;
srom_1(16449) <= 16219440;
srom_1(16450) <= 15995231;
srom_1(16451) <= 15735351;
srom_1(16452) <= 15441020;
srom_1(16453) <= 15113618;
srom_1(16454) <= 14754680;
srom_1(16455) <= 14365889;
srom_1(16456) <= 13949069;
srom_1(16457) <= 13506174;
srom_1(16458) <= 13039281;
srom_1(16459) <= 12550579;
srom_1(16460) <= 12042360;
srom_1(16461) <= 11517008;
srom_1(16462) <= 10976985;
srom_1(16463) <= 10424825;
srom_1(16464) <= 9863116;
srom_1(16465) <= 9294492;
srom_1(16466) <= 8721621;
srom_1(16467) <= 8147188;
srom_1(16468) <= 7573887;
srom_1(16469) <= 7004407;
srom_1(16470) <= 6441417;
srom_1(16471) <= 5887559;
srom_1(16472) <= 5345429;
srom_1(16473) <= 4817569;
srom_1(16474) <= 4306455;
srom_1(16475) <= 3814484;
srom_1(16476) <= 3343963;
srom_1(16477) <= 2897097;
srom_1(16478) <= 2475983;
srom_1(16479) <= 2082596;
srom_1(16480) <= 1718779;
srom_1(16481) <= 1386240;
srom_1(16482) <= 1086537;
srom_1(16483) <= 821076;
srom_1(16484) <= 591101;
srom_1(16485) <= 397692;
srom_1(16486) <= 241755;
srom_1(16487) <= 124022;
srom_1(16488) <= 45044;
srom_1(16489) <= 5192;
srom_1(16490) <= 4652;
srom_1(16491) <= 43428;
srom_1(16492) <= 121337;
srom_1(16493) <= 238014;
srom_1(16494) <= 392912;
srom_1(16495) <= 585305;
srom_1(16496) <= 814290;
srom_1(16497) <= 1078794;
srom_1(16498) <= 1377575;
srom_1(16499) <= 1709234;
srom_1(16500) <= 2072215;
srom_1(16501) <= 2464816;
srom_1(16502) <= 2885195;
srom_1(16503) <= 3331382;
srom_1(16504) <= 3801283;
srom_1(16505) <= 4292697;
srom_1(16506) <= 4803317;
srom_1(16507) <= 5330750;
srom_1(16508) <= 5872522;
srom_1(16509) <= 6426094;
srom_1(16510) <= 6988868;
srom_1(16511) <= 7558206;
srom_1(16512) <= 8131437;
srom_1(16513) <= 8705875;
srom_1(16514) <= 9278826;
srom_1(16515) <= 9847601;
srom_1(16516) <= 10409535;
srom_1(16517) <= 10961992;
srom_1(16518) <= 11502381;
srom_1(16519) <= 12028169;
srom_1(16520) <= 12536890;
srom_1(16521) <= 13026158;
srom_1(16522) <= 13493679;
srom_1(16523) <= 13937261;
srom_1(16524) <= 14354823;
srom_1(16525) <= 14744407;
srom_1(16526) <= 15104187;
srom_1(16527) <= 15432475;
srom_1(16528) <= 15727732;
srom_1(16529) <= 15988574;
srom_1(16530) <= 16213776;
srom_1(16531) <= 16402284;
srom_1(16532) <= 16553213;
srom_1(16533) <= 16665855;
srom_1(16534) <= 16739682;
srom_1(16535) <= 16774348;
srom_1(16536) <= 16769691;
srom_1(16537) <= 16725731;
srom_1(16538) <= 16642676;
srom_1(16539) <= 16520915;
srom_1(16540) <= 16361019;
srom_1(16541) <= 16163738;
srom_1(16542) <= 15929996;
srom_1(16543) <= 15660890;
srom_1(16544) <= 15357681;
srom_1(16545) <= 15021793;
srom_1(16546) <= 14654799;
srom_1(16547) <= 14258420;
srom_1(16548) <= 13834517;
srom_1(16549) <= 13385075;
srom_1(16550) <= 12912203;
srom_1(16551) <= 12418119;
srom_1(16552) <= 11905138;
srom_1(16553) <= 11375668;
srom_1(16554) <= 10832190;
srom_1(16555) <= 10277254;
srom_1(16556) <= 9713460;
srom_1(16557) <= 9143455;
srom_1(16558) <= 8569909;
srom_1(16559) <= 7995513;
srom_1(16560) <= 7422961;
srom_1(16561) <= 6854937;
srom_1(16562) <= 6294104;
srom_1(16563) <= 5743094;
srom_1(16564) <= 5204489;
srom_1(16565) <= 4680816;
srom_1(16566) <= 4174530;
srom_1(16567) <= 3688005;
srom_1(16568) <= 3223523;
srom_1(16569) <= 2783261;
srom_1(16570) <= 2369285;
srom_1(16571) <= 1983536;
srom_1(16572) <= 1627822;
srom_1(16573) <= 1303812;
srom_1(16574) <= 1013025;
srom_1(16575) <= 756825;
srom_1(16576) <= 536412;
srom_1(16577) <= 352822;
srom_1(16578) <= 206914;
srom_1(16579) <= 99372;
srom_1(16580) <= 30702;
srom_1(16581) <= 1225;
srom_1(16582) <= 11079;
srom_1(16583) <= 60218;
srom_1(16584) <= 148412;
srom_1(16585) <= 275247;
srom_1(16586) <= 440128;
srom_1(16587) <= 642282;
srom_1(16588) <= 880762;
srom_1(16589) <= 1154449;
srom_1(16590) <= 1462058;
srom_1(16591) <= 1802149;
srom_1(16592) <= 2173126;
srom_1(16593) <= 2573250;
srom_1(16594) <= 3000644;
srom_1(16595) <= 3453304;
srom_1(16596) <= 3929107;
srom_1(16597) <= 4425822;
srom_1(16598) <= 4941120;
srom_1(16599) <= 5472585;
srom_1(16600) <= 6017723;
srom_1(16601) <= 6573980;
srom_1(16602) <= 7138746;
srom_1(16603) <= 7709373;
srom_1(16604) <= 8283185;
srom_1(16605) <= 8857492;
srom_1(16606) <= 9429600;
srom_1(16607) <= 9996826;
srom_1(16608) <= 10556511;
srom_1(16609) <= 11106030;
srom_1(16610) <= 11642805;
srom_1(16611) <= 12164321;
srom_1(16612) <= 12668131;
srom_1(16613) <= 13151873;
srom_1(16614) <= 13613279;
srom_1(16615) <= 14050184;
srom_1(16616) <= 14460540;
srom_1(16617) <= 14842422;
srom_1(16618) <= 15194041;
srom_1(16619) <= 15513746;
srom_1(16620) <= 15800039;
srom_1(16621) <= 16051578;
srom_1(16622) <= 16267182;
srom_1(16623) <= 16445841;
srom_1(16624) <= 16586716;
srom_1(16625) <= 16689148;
srom_1(16626) <= 16752656;
srom_1(16627) <= 16776942;
srom_1(16628) <= 16761892;
srom_1(16629) <= 16707577;
srom_1(16630) <= 16614252;
srom_1(16631) <= 16482353;
srom_1(16632) <= 16312500;
srom_1(16633) <= 16105490;
srom_1(16634) <= 15862292;
srom_1(16635) <= 15584047;
srom_1(16636) <= 15272061;
srom_1(16637) <= 14927796;
srom_1(16638) <= 14552866;
srom_1(16639) <= 14149030;
srom_1(16640) <= 13718181;
srom_1(16641) <= 13262340;
srom_1(16642) <= 12783645;
srom_1(16643) <= 12284339;
srom_1(16644) <= 11766765;
srom_1(16645) <= 11233350;
srom_1(16646) <= 10686595;
srom_1(16647) <= 10129064;
srom_1(16648) <= 9563371;
srom_1(16649) <= 8992170;
srom_1(16650) <= 8418138;
srom_1(16651) <= 7843967;
srom_1(16652) <= 7272351;
srom_1(16653) <= 6705969;
srom_1(16654) <= 6147477;
srom_1(16655) <= 5599495;
srom_1(16656) <= 5064592;
srom_1(16657) <= 4545277;
srom_1(16658) <= 4043984;
srom_1(16659) <= 3563065;
srom_1(16660) <= 3104774;
srom_1(16661) <= 2671261;
srom_1(16662) <= 2264558;
srom_1(16663) <= 1886574;
srom_1(16664) <= 1539079;
srom_1(16665) <= 1223705;
srom_1(16666) <= 941929;
srom_1(16667) <= 695073;
srom_1(16668) <= 484294;
srom_1(16669) <= 310582;
srom_1(16670) <= 174750;
srom_1(16671) <= 77436;
srom_1(16672) <= 19096;
srom_1(16673) <= 4;
srom_1(16674) <= 20248;
srom_1(16675) <= 79735;
srom_1(16676) <= 178184;
srom_1(16677) <= 315136;
srom_1(16678) <= 489946;
srom_1(16679) <= 701796;
srom_1(16680) <= 949692;
srom_1(16681) <= 1232472;
srom_1(16682) <= 1548809;
srom_1(16683) <= 1897221;
srom_1(16684) <= 2276072;
srom_1(16685) <= 2683588;
srom_1(16686) <= 3117856;
srom_1(16687) <= 3576841;
srom_1(16688) <= 4058390;
srom_1(16689) <= 4560244;
srom_1(16690) <= 5080052;
srom_1(16691) <= 5615374;
srom_1(16692) <= 6163700;
srom_1(16693) <= 6722460;
srom_1(16694) <= 7289034;
srom_1(16695) <= 7860763;
srom_1(16696) <= 8434968;
srom_1(16697) <= 9008955;
srom_1(16698) <= 9580033;
srom_1(16699) <= 10145525;
srom_1(16700) <= 10702777;
srom_1(16701) <= 11249178;
srom_1(16702) <= 11782164;
srom_1(16703) <= 12299237;
srom_1(16704) <= 12797971;
srom_1(16705) <= 13276029;
srom_1(16706) <= 13731167;
srom_1(16707) <= 14161253;
srom_1(16708) <= 14564269;
srom_1(16709) <= 14938324;
srom_1(16710) <= 15281666;
srom_1(16711) <= 15592684;
srom_1(16712) <= 15869920;
srom_1(16713) <= 16112073;
srom_1(16714) <= 16318008;
srom_1(16715) <= 16486760;
srom_1(16716) <= 16617536;
srom_1(16717) <= 16709725;
srom_1(16718) <= 16762892;
srom_1(16719) <= 16776790;
srom_1(16720) <= 16751352;
srom_1(16721) <= 16686699;
srom_1(16722) <= 16583134;
srom_1(16723) <= 16441141;
srom_1(16724) <= 16261387;
srom_1(16725) <= 16044715;
srom_1(16726) <= 15792141;
srom_1(16727) <= 15504849;
srom_1(16728) <= 15184187;
srom_1(16729) <= 14831658;
srom_1(16730) <= 14448915;
srom_1(16731) <= 14037753;
srom_1(16732) <= 13600101;
srom_1(16733) <= 13138010;
srom_1(16734) <= 12653647;
srom_1(16735) <= 12149284;
srom_1(16736) <= 11627287;
srom_1(16737) <= 11090101;
srom_1(16738) <= 10540248;
srom_1(16739) <= 9980305;
srom_1(16740) <= 9412897;
srom_1(16741) <= 8840687;
srom_1(16742) <= 8266357;
srom_1(16743) <= 7692599;
srom_1(16744) <= 7122106;
srom_1(16745) <= 6557552;
srom_1(16746) <= 6001584;
srom_1(16747) <= 5456810;
srom_1(16748) <= 4925784;
srom_1(16749) <= 4410996;
srom_1(16750) <= 3914861;
srom_1(16751) <= 3439704;
srom_1(16752) <= 2987755;
srom_1(16753) <= 2561132;
srom_1(16754) <= 2161836;
srom_1(16755) <= 1791740;
srom_1(16756) <= 1452578;
srom_1(16757) <= 1145942;
srom_1(16758) <= 873270;
srom_1(16759) <= 635839;
srom_1(16760) <= 434764;
srom_1(16761) <= 270987;
srom_1(16762) <= 145276;
srom_1(16763) <= 58222;
srom_1(16764) <= 10231;
srom_1(16765) <= 1529;
srom_1(16766) <= 32157;
srom_1(16767) <= 101972;
srom_1(16768) <= 210645;
srom_1(16769) <= 357668;
srom_1(16770) <= 542350;
srom_1(16771) <= 763826;
srom_1(16772) <= 1021058;
srom_1(16773) <= 1312838;
srom_1(16774) <= 1637799;
srom_1(16775) <= 1994417;
srom_1(16776) <= 2381020;
srom_1(16777) <= 2795794;
srom_1(16778) <= 3236795;
srom_1(16779) <= 3701954;
srom_1(16780) <= 4189091;
srom_1(16781) <= 4695920;
srom_1(16782) <= 5220066;
srom_1(16783) <= 5759071;
srom_1(16784) <= 6310406;
srom_1(16785) <= 6871486;
srom_1(16786) <= 7439681;
srom_1(16787) <= 8012326;
srom_1(16788) <= 8586735;
srom_1(16789) <= 9160215;
srom_1(16790) <= 9730077;
srom_1(16791) <= 10293648;
srom_1(16792) <= 10848286;
srom_1(16793) <= 11391389;
srom_1(16794) <= 11920412;
srom_1(16795) <= 12432872;
srom_1(16796) <= 12926368;
srom_1(16797) <= 13398584;
srom_1(16798) <= 13847307;
srom_1(16799) <= 14270432;
srom_1(16800) <= 14665976;
srom_1(16801) <= 15032082;
srom_1(16802) <= 15367035;
srom_1(16803) <= 15669264;
srom_1(16804) <= 15937351;
srom_1(16805) <= 16170040;
srom_1(16806) <= 16366239;
srom_1(16807) <= 16525028;
srom_1(16808) <= 16645662;
srom_1(16809) <= 16727576;
srom_1(16810) <= 16770386;
srom_1(16811) <= 16773891;
srom_1(16812) <= 16738075;
srom_1(16813) <= 16663105;
srom_1(16814) <= 16549333;
srom_1(16815) <= 16397292;
srom_1(16816) <= 16207696;
srom_1(16817) <= 15981434;
srom_1(16818) <= 15719566;
srom_1(16819) <= 15423321;
srom_1(16820) <= 15094088;
srom_1(16821) <= 14733410;
srom_1(16822) <= 14342980;
srom_1(16823) <= 13924627;
srom_1(16824) <= 13480314;
srom_1(16825) <= 13012124;
srom_1(16826) <= 12522253;
srom_1(16827) <= 12012998;
srom_1(16828) <= 11486747;
srom_1(16829) <= 10945968;
srom_1(16830) <= 10393196;
srom_1(16831) <= 9831024;
srom_1(16832) <= 9262088;
srom_1(16833) <= 8689056;
srom_1(16834) <= 8114616;
srom_1(16835) <= 7541460;
srom_1(16836) <= 6972276;
srom_1(16837) <= 6409734;
srom_1(16838) <= 5856472;
srom_1(16839) <= 5315084;
srom_1(16840) <= 4788109;
srom_1(16841) <= 4278017;
srom_1(16842) <= 3787202;
srom_1(16843) <= 3317964;
srom_1(16844) <= 2872504;
srom_1(16845) <= 2452911;
srom_1(16846) <= 2061153;
srom_1(16847) <= 1699066;
srom_1(16848) <= 1368349;
srom_1(16849) <= 1070552;
srom_1(16850) <= 807072;
srom_1(16851) <= 579144;
srom_1(16852) <= 387838;
srom_1(16853) <= 234050;
srom_1(16854) <= 118501;
srom_1(16855) <= 41734;
srom_1(16856) <= 4108;
srom_1(16857) <= 5800;
srom_1(16858) <= 46802;
srom_1(16859) <= 126922;
srom_1(16860) <= 245783;
srom_1(16861) <= 402829;
srom_1(16862) <= 597323;
srom_1(16863) <= 828353;
srom_1(16864) <= 1094835;
srom_1(16865) <= 1395521;
srom_1(16866) <= 1729000;
srom_1(16867) <= 2093707;
srom_1(16868) <= 2487934;
srom_1(16869) <= 2909831;
srom_1(16870) <= 3357420;
srom_1(16871) <= 3828601;
srom_1(16872) <= 4321167;
srom_1(16873) <= 4832805;
srom_1(16874) <= 5361119;
srom_1(16875) <= 5903629;
srom_1(16876) <= 6457792;
srom_1(16877) <= 7021009;
srom_1(16878) <= 7590639;
srom_1(16879) <= 8164012;
srom_1(16880) <= 8738437;
srom_1(16881) <= 9311223;
srom_1(16882) <= 9879681;
srom_1(16883) <= 10441148;
srom_1(16884) <= 10992989;
srom_1(16885) <= 11532618;
srom_1(16886) <= 12057503;
srom_1(16887) <= 12565183;
srom_1(16888) <= 13053278;
srom_1(16889) <= 13519499;
srom_1(16890) <= 13961659;
srom_1(16891) <= 14377686;
srom_1(16892) <= 14765627;
srom_1(16893) <= 15123665;
srom_1(16894) <= 15450119;
srom_1(16895) <= 15743460;
srom_1(16896) <= 16002311;
srom_1(16897) <= 16225459;
srom_1(16898) <= 16411857;
srom_1(16899) <= 16560632;
srom_1(16900) <= 16671085;
srom_1(16901) <= 16742698;
srom_1(16902) <= 16775137;
srom_1(16903) <= 16768248;
srom_1(16904) <= 16722064;
srom_1(16905) <= 16636801;
srom_1(16906) <= 16512860;
srom_1(16907) <= 16350822;
srom_1(16908) <= 16151446;
srom_1(16909) <= 15915667;
srom_1(16910) <= 15644592;
srom_1(16911) <= 15339490;
srom_1(16912) <= 15001794;
srom_1(16913) <= 14633086;
srom_1(16914) <= 14235095;
srom_1(16915) <= 13809689;
srom_1(16916) <= 13358861;
srom_1(16917) <= 12884725;
srom_1(16918) <= 12389506;
srom_1(16919) <= 11875526;
srom_1(16920) <= 11345194;
srom_1(16921) <= 10800997;
srom_1(16922) <= 10245488;
srom_1(16923) <= 9681272;
srom_1(16924) <= 9110993;
srom_1(16925) <= 8537327;
srom_1(16926) <= 7962964;
srom_1(16927) <= 7390597;
srom_1(16928) <= 6822910;
srom_1(16929) <= 6262565;
srom_1(16930) <= 5712189;
srom_1(16931) <= 5174364;
srom_1(16932) <= 4651612;
srom_1(16933) <= 4146384;
srom_1(16934) <= 3661049;
srom_1(16935) <= 3197884;
srom_1(16936) <= 2759059;
srom_1(16937) <= 2346633;
srom_1(16938) <= 1962541;
srom_1(16939) <= 1608582;
srom_1(16940) <= 1286417;
srom_1(16941) <= 997557;
srom_1(16942) <= 743356;
srom_1(16943) <= 525006;
srom_1(16944) <= 343531;
srom_1(16945) <= 199782;
srom_1(16946) <= 94434;
srom_1(16947) <= 27979;
srom_1(16948) <= 731;
srom_1(16949) <= 12816;
srom_1(16950) <= 64178;
srom_1(16951) <= 154577;
srom_1(16952) <= 283587;
srom_1(16953) <= 450605;
srom_1(16954) <= 654847;
srom_1(16955) <= 895355;
srom_1(16956) <= 1171001;
srom_1(16957) <= 1480493;
srom_1(16958) <= 1822380;
srom_1(16959) <= 2195058;
srom_1(16960) <= 2596780;
srom_1(16961) <= 3025662;
srom_1(16962) <= 3479692;
srom_1(16963) <= 3956742;
srom_1(16964) <= 4454574;
srom_1(16965) <= 4970855;
srom_1(16966) <= 5503162;
srom_1(16967) <= 6049000;
srom_1(16968) <= 6605810;
srom_1(16969) <= 7170979;
srom_1(16970) <= 7741859;
srom_1(16971) <= 8315771;
srom_1(16972) <= 8890025;
srom_1(16973) <= 9461928;
srom_1(16974) <= 10028797;
srom_1(16975) <= 10587975;
srom_1(16976) <= 11136840;
srom_1(16977) <= 11672817;
srom_1(16978) <= 12193393;
srom_1(16979) <= 12696127;
srom_1(16980) <= 13178662;
srom_1(16981) <= 13638734;
srom_1(16982) <= 14074187;
srom_1(16983) <= 14482979;
srom_1(16984) <= 14863191;
srom_1(16985) <= 15213042;
srom_1(16986) <= 15530891;
srom_1(16987) <= 15815248;
srom_1(16988) <= 16064778;
srom_1(16989) <= 16278312;
srom_1(16990) <= 16454849;
srom_1(16991) <= 16593560;
srom_1(16992) <= 16693795;
srom_1(16993) <= 16755085;
srom_1(16994) <= 16777141;
srom_1(16995) <= 16759860;
srom_1(16996) <= 16703324;
srom_1(16997) <= 16607797;
srom_1(16998) <= 16473728;
srom_1(16999) <= 16301745;
srom_1(17000) <= 16092654;
srom_1(17001) <= 15847436;
srom_1(17002) <= 15567241;
srom_1(17003) <= 15253384;
srom_1(17004) <= 14907335;
srom_1(17005) <= 14530717;
srom_1(17006) <= 14125297;
srom_1(17007) <= 13692975;
srom_1(17008) <= 13235780;
srom_1(17009) <= 12755854;
srom_1(17010) <= 12255449;
srom_1(17011) <= 11736911;
srom_1(17012) <= 11202672;
srom_1(17013) <= 10655237;
srom_1(17014) <= 10097172;
srom_1(17015) <= 9531096;
srom_1(17016) <= 8959662;
srom_1(17017) <= 8385550;
srom_1(17018) <= 7811452;
srom_1(17019) <= 7240061;
srom_1(17020) <= 6674056;
srom_1(17021) <= 6116091;
srom_1(17022) <= 5568783;
srom_1(17023) <= 5034697;
srom_1(17024) <= 4516340;
srom_1(17025) <= 4016140;
srom_1(17026) <= 3536445;
srom_1(17027) <= 3079503;
srom_1(17028) <= 2647457;
srom_1(17029) <= 2242334;
srom_1(17030) <= 1866033;
srom_1(17031) <= 1520318;
srom_1(17032) <= 1206811;
srom_1(17033) <= 926981;
srom_1(17034) <= 682142;
srom_1(17035) <= 473442;
srom_1(17036) <= 301858;
srom_1(17037) <= 168195;
srom_1(17038) <= 73081;
srom_1(17039) <= 16962;
srom_1(17040) <= 100;
srom_1(17041) <= 22574;
srom_1(17042) <= 84280;
srom_1(17043) <= 184927;
srom_1(17044) <= 324045;
srom_1(17045) <= 500980;
srom_1(17046) <= 714902;
srom_1(17047) <= 964810;
srom_1(17048) <= 1249530;
srom_1(17049) <= 1567727;
srom_1(17050) <= 1917910;
srom_1(17051) <= 2298437;
srom_1(17052) <= 2707522;
srom_1(17053) <= 3143248;
srom_1(17054) <= 3603571;
srom_1(17055) <= 4086333;
srom_1(17056) <= 4589270;
srom_1(17057) <= 5110023;
srom_1(17058) <= 5646150;
srom_1(17059) <= 6195138;
srom_1(17060) <= 6754412;
srom_1(17061) <= 7321349;
srom_1(17062) <= 7893290;
srom_1(17063) <= 8467555;
srom_1(17064) <= 9041449;
srom_1(17065) <= 9612282;
srom_1(17066) <= 10177376;
srom_1(17067) <= 10734083;
srom_1(17068) <= 11279791;
srom_1(17069) <= 11811940;
srom_1(17070) <= 12328037;
srom_1(17071) <= 12825661;
srom_1(17072) <= 13302477;
srom_1(17073) <= 13756251;
srom_1(17074) <= 14184854;
srom_1(17075) <= 14586276;
srom_1(17076) <= 14958636;
srom_1(17077) <= 15300186;
srom_1(17078) <= 15609325;
srom_1(17079) <= 15884604;
srom_1(17080) <= 16124732;
srom_1(17081) <= 16328583;
srom_1(17082) <= 16495200;
srom_1(17083) <= 16623802;
srom_1(17084) <= 16713787;
srom_1(17085) <= 16764732;
srom_1(17086) <= 16776399;
srom_1(17087) <= 16748732;
srom_1(17088) <= 16681862;
srom_1(17089) <= 16576102;
srom_1(17090) <= 16431949;
srom_1(17091) <= 16250077;
srom_1(17092) <= 16031339;
srom_1(17093) <= 15776763;
srom_1(17094) <= 15487541;
srom_1(17095) <= 15165029;
srom_1(17096) <= 14810741;
srom_1(17097) <= 14426337;
srom_1(17098) <= 14013620;
srom_1(17099) <= 13574525;
srom_1(17100) <= 13111112;
srom_1(17101) <= 12625554;
srom_1(17102) <= 12120127;
srom_1(17103) <= 11597201;
srom_1(17104) <= 11059229;
srom_1(17105) <= 10508734;
srom_1(17106) <= 9948297;
srom_1(17107) <= 9380546;
srom_1(17108) <= 8808143;
srom_1(17109) <= 8233773;
srom_1(17110) <= 7660129;
srom_1(17111) <= 7089901;
srom_1(17112) <= 6525764;
srom_1(17113) <= 5970361;
srom_1(17114) <= 5426299;
srom_1(17115) <= 4896128;
srom_1(17116) <= 4382334;
srom_1(17117) <= 3887328;
srom_1(17118) <= 3413429;
srom_1(17119) <= 2962860;
srom_1(17120) <= 2537735;
srom_1(17121) <= 2140047;
srom_1(17122) <= 1771660;
srom_1(17123) <= 1434302;
srom_1(17124) <= 1129556;
srom_1(17125) <= 858849;
srom_1(17126) <= 623452;
srom_1(17127) <= 424469;
srom_1(17128) <= 262832;
srom_1(17129) <= 139300;
srom_1(17130) <= 54452;
srom_1(17131) <= 8685;
srom_1(17132) <= 2215;
srom_1(17133) <= 35071;
srom_1(17134) <= 107100;
srom_1(17135) <= 217964;
srom_1(17136) <= 367143;
srom_1(17137) <= 553937;
srom_1(17138) <= 777470;
srom_1(17139) <= 1036695;
srom_1(17140) <= 1330396;
srom_1(17141) <= 1657194;
srom_1(17142) <= 2015559;
srom_1(17143) <= 2403809;
srom_1(17144) <= 2820124;
srom_1(17145) <= 3262552;
srom_1(17146) <= 3729017;
srom_1(17147) <= 4217333;
srom_1(17148) <= 4725209;
srom_1(17149) <= 5250264;
srom_1(17150) <= 5790036;
srom_1(17151) <= 6341993;
srom_1(17152) <= 6903548;
srom_1(17153) <= 7472067;
srom_1(17154) <= 8044884;
srom_1(17155) <= 8619312;
srom_1(17156) <= 9192659;
srom_1(17157) <= 9762235;
srom_1(17158) <= 10325370;
srom_1(17159) <= 10879423;
srom_1(17160) <= 11421795;
srom_1(17161) <= 11949944;
srom_1(17162) <= 12461392;
srom_1(17163) <= 12953742;
srom_1(17164) <= 13424684;
srom_1(17165) <= 13872010;
srom_1(17166) <= 14293623;
srom_1(17167) <= 14687545;
srom_1(17168) <= 15051929;
srom_1(17169) <= 15385067;
srom_1(17170) <= 15685395;
srom_1(17171) <= 15951507;
srom_1(17172) <= 16182154;
srom_1(17173) <= 16376253;
srom_1(17174) <= 16532897;
srom_1(17175) <= 16651348;
srom_1(17176) <= 16731053;
srom_1(17177) <= 16771638;
srom_1(17178) <= 16772911;
srom_1(17179) <= 16734868;
srom_1(17180) <= 16657686;
srom_1(17181) <= 16541727;
srom_1(17182) <= 16387536;
srom_1(17183) <= 16195835;
srom_1(17184) <= 15967523;
srom_1(17185) <= 15703671;
srom_1(17186) <= 15405516;
srom_1(17187) <= 15074457;
srom_1(17188) <= 14712045;
srom_1(17189) <= 14319981;
srom_1(17190) <= 13900102;
srom_1(17191) <= 13454378;
srom_1(17192) <= 12984899;
srom_1(17193) <= 12493866;
srom_1(17194) <= 11983582;
srom_1(17195) <= 11456440;
srom_1(17196) <= 10914912;
srom_1(17197) <= 10361537;
srom_1(17198) <= 9798911;
srom_1(17199) <= 9229671;
srom_1(17200) <= 8656487;
srom_1(17201) <= 8082047;
srom_1(17202) <= 7509045;
srom_1(17203) <= 6940167;
srom_1(17204) <= 6378081;
srom_1(17205) <= 5825423;
srom_1(17206) <= 5284785;
srom_1(17207) <= 4758702;
srom_1(17208) <= 4249641;
srom_1(17209) <= 3759989;
srom_1(17210) <= 3292042;
srom_1(17211) <= 2847994;
srom_1(17212) <= 2429929;
srom_1(17213) <= 2039805;
srom_1(17214) <= 1679454;
srom_1(17215) <= 1350563;
srom_1(17216) <= 1054677;
srom_1(17217) <= 793182;
srom_1(17218) <= 567305;
srom_1(17219) <= 378104;
srom_1(17220) <= 226467;
srom_1(17221) <= 113105;
srom_1(17222) <= 38551;
srom_1(17223) <= 3152;
srom_1(17224) <= 7075;
srom_1(17225) <= 50303;
srom_1(17226) <= 132632;
srom_1(17227) <= 253675;
srom_1(17228) <= 412867;
srom_1(17229) <= 609459;
srom_1(17230) <= 842530;
srom_1(17231) <= 1110988;
srom_1(17232) <= 1413572;
srom_1(17233) <= 1748865;
srom_1(17234) <= 2115294;
srom_1(17235) <= 2511141;
srom_1(17236) <= 2934549;
srom_1(17237) <= 3383534;
srom_1(17238) <= 3855988;
srom_1(17239) <= 4349698;
srom_1(17240) <= 4862348;
srom_1(17241) <= 5391533;
srom_1(17242) <= 5934773;
srom_1(17243) <= 6489519;
srom_1(17244) <= 7053171;
srom_1(17245) <= 7623085;
srom_1(17246) <= 8196590;
srom_1(17247) <= 8770994;
srom_1(17248) <= 9343606;
srom_1(17249) <= 9911739;
srom_1(17250) <= 10472729;
srom_1(17251) <= 11023947;
srom_1(17252) <= 11562806;
srom_1(17253) <= 12086781;
srom_1(17254) <= 12593413;
srom_1(17255) <= 13080328;
srom_1(17256) <= 13545242;
srom_1(17257) <= 13985974;
srom_1(17258) <= 14400458;
srom_1(17259) <= 14786751;
srom_1(17260) <= 15143041;
srom_1(17261) <= 15467657;
srom_1(17262) <= 15759076;
srom_1(17263) <= 16015933;
srom_1(17264) <= 16237023;
srom_1(17265) <= 16421309;
srom_1(17266) <= 16567927;
srom_1(17267) <= 16676189;
srom_1(17268) <= 16745588;
srom_1(17269) <= 16775798;
srom_1(17270) <= 16766678;
srom_1(17271) <= 16718270;
srom_1(17272) <= 16630802;
srom_1(17273) <= 16504682;
srom_1(17274) <= 16340504;
srom_1(17275) <= 16139037;
srom_1(17276) <= 15901225;
srom_1(17277) <= 15628184;
srom_1(17278) <= 15321194;
srom_1(17279) <= 14981695;
srom_1(17280) <= 14611279;
srom_1(17281) <= 14211682;
srom_1(17282) <= 13784779;
srom_1(17283) <= 13332571;
srom_1(17284) <= 12857180;
srom_1(17285) <= 12360834;
srom_1(17286) <= 11845860;
srom_1(17287) <= 11314675;
srom_1(17288) <= 10769768;
srom_1(17289) <= 10213695;
srom_1(17290) <= 9649063;
srom_1(17291) <= 9078521;
srom_1(17292) <= 8504744;
srom_1(17293) <= 7930422;
srom_1(17294) <= 7358248;
srom_1(17295) <= 6790906;
srom_1(17296) <= 6231057;
srom_1(17297) <= 5681325;
srom_1(17298) <= 5144288;
srom_1(17299) <= 4622465;
srom_1(17300) <= 4118303;
srom_1(17301) <= 3634165;
srom_1(17302) <= 3172323;
srom_1(17303) <= 2734942;
srom_1(17304) <= 2324073;
srom_1(17305) <= 1941642;
srom_1(17306) <= 1589444;
srom_1(17307) <= 1269129;
srom_1(17308) <= 982200;
srom_1(17309) <= 730002;
srom_1(17310) <= 513717;
srom_1(17311) <= 334361;
srom_1(17312) <= 192774;
srom_1(17313) <= 89620;
srom_1(17314) <= 25383;
srom_1(17315) <= 364;
srom_1(17316) <= 14680;
srom_1(17317) <= 68265;
srom_1(17318) <= 160866;
srom_1(17319) <= 292050;
srom_1(17320) <= 461202;
srom_1(17321) <= 667528;
srom_1(17322) <= 910060;
srom_1(17323) <= 1187663;
srom_1(17324) <= 1499032;
srom_1(17325) <= 1842710;
srom_1(17326) <= 2217083;
srom_1(17327) <= 2620397;
srom_1(17328) <= 3050760;
srom_1(17329) <= 3506154;
srom_1(17330) <= 3984444;
srom_1(17331) <= 4483386;
srom_1(17332) <= 5000641;
srom_1(17333) <= 5533783;
srom_1(17334) <= 6080313;
srom_1(17335) <= 6637667;
srom_1(17336) <= 7203231;
srom_1(17337) <= 7774355;
srom_1(17338) <= 8348358;
srom_1(17339) <= 8922551;
srom_1(17340) <= 9494240;
srom_1(17341) <= 10060744;
srom_1(17342) <= 10619406;
srom_1(17343) <= 11167608;
srom_1(17344) <= 11702778;
srom_1(17345) <= 12222407;
srom_1(17346) <= 12724058;
srom_1(17347) <= 13205378;
srom_1(17348) <= 13664111;
srom_1(17349) <= 14098105;
srom_1(17350) <= 14505326;
srom_1(17351) <= 14883863;
srom_1(17352) <= 15231941;
srom_1(17353) <= 15547929;
srom_1(17354) <= 15830344;
srom_1(17355) <= 16077863;
srom_1(17356) <= 16289323;
srom_1(17357) <= 16463735;
srom_1(17358) <= 16600280;
srom_1(17359) <= 16698317;
srom_1(17360) <= 16757387;
srom_1(17361) <= 16777213;
srom_1(17362) <= 16757702;
srom_1(17363) <= 16698946;
srom_1(17364) <= 16601219;
srom_1(17365) <= 16464981;
srom_1(17366) <= 16290869;
srom_1(17367) <= 16079702;
srom_1(17368) <= 15832468;
srom_1(17369) <= 15550327;
srom_1(17370) <= 15234603;
srom_1(17371) <= 14886775;
srom_1(17372) <= 14508475;
srom_1(17373) <= 14101477;
srom_1(17374) <= 13667690;
srom_1(17375) <= 13209147;
srom_1(17376) <= 12727998;
srom_1(17377) <= 12226501;
srom_1(17378) <= 11707007;
srom_1(17379) <= 11171952;
srom_1(17380) <= 10623844;
srom_1(17381) <= 10065255;
srom_1(17382) <= 9498803;
srom_1(17383) <= 8927145;
srom_1(17384) <= 8352962;
srom_1(17385) <= 7778946;
srom_1(17386) <= 7207789;
srom_1(17387) <= 6642169;
srom_1(17388) <= 6084739;
srom_1(17389) <= 5538112;
srom_1(17390) <= 5004853;
srom_1(17391) <= 4487461;
srom_1(17392) <= 3988362;
srom_1(17393) <= 3509898;
srom_1(17394) <= 3054312;
srom_1(17395) <= 2623741;
srom_1(17396) <= 2220202;
srom_1(17397) <= 1845590;
srom_1(17398) <= 1501660;
srom_1(17399) <= 1190025;
srom_1(17400) <= 912147;
srom_1(17401) <= 669328;
srom_1(17402) <= 462708;
srom_1(17403) <= 293255;
srom_1(17404) <= 161764;
srom_1(17405) <= 68852;
srom_1(17406) <= 14954;
srom_1(17407) <= 322;
srom_1(17408) <= 25026;
srom_1(17409) <= 88950;
srom_1(17410) <= 191794;
srom_1(17411) <= 333076;
srom_1(17412) <= 512132;
srom_1(17413) <= 728124;
srom_1(17414) <= 980039;
srom_1(17415) <= 1266695;
srom_1(17416) <= 1586748;
srom_1(17417) <= 1938698;
srom_1(17418) <= 2320893;
srom_1(17419) <= 2731542;
srom_1(17420) <= 3168719;
srom_1(17421) <= 3630373;
srom_1(17422) <= 4114341;
srom_1(17423) <= 4618352;
srom_1(17424) <= 5140043;
srom_1(17425) <= 5676968;
srom_1(17426) <= 6226608;
srom_1(17427) <= 6786387;
srom_1(17428) <= 7353679;
srom_1(17429) <= 7925825;
srom_1(17430) <= 8500140;
srom_1(17431) <= 9073933;
srom_1(17432) <= 9644512;
srom_1(17433) <= 10209201;
srom_1(17434) <= 10765353;
srom_1(17435) <= 11310360;
srom_1(17436) <= 11841665;
srom_1(17437) <= 12356778;
srom_1(17438) <= 12853283;
srom_1(17439) <= 13328852;
srom_1(17440) <= 13781253;
srom_1(17441) <= 14208367;
srom_1(17442) <= 14608190;
srom_1(17443) <= 14978848;
srom_1(17444) <= 15318601;
srom_1(17445) <= 15625858;
srom_1(17446) <= 15899176;
srom_1(17447) <= 16137275;
srom_1(17448) <= 16339037;
srom_1(17449) <= 16503517;
srom_1(17450) <= 16629944;
srom_1(17451) <= 16717724;
srom_1(17452) <= 16766446;
srom_1(17453) <= 16775882;
srom_1(17454) <= 16745986;
srom_1(17455) <= 16676900;
srom_1(17456) <= 16568948;
srom_1(17457) <= 16422635;
srom_1(17458) <= 16238647;
srom_1(17459) <= 16017849;
srom_1(17460) <= 15761274;
srom_1(17461) <= 15470126;
srom_1(17462) <= 15145770;
srom_1(17463) <= 14789728;
srom_1(17464) <= 14403668;
srom_1(17465) <= 13989402;
srom_1(17466) <= 13548872;
srom_1(17467) <= 13084144;
srom_1(17468) <= 12597396;
srom_1(17469) <= 12090912;
srom_1(17470) <= 11567067;
srom_1(17471) <= 11028317;
srom_1(17472) <= 10477188;
srom_1(17473) <= 9916266;
srom_1(17474) <= 9348179;
srom_1(17475) <= 8775593;
srom_1(17476) <= 8201192;
srom_1(17477) <= 7627670;
srom_1(17478) <= 7057716;
srom_1(17479) <= 6494004;
srom_1(17480) <= 5939175;
srom_1(17481) <= 5395833;
srom_1(17482) <= 4866525;
srom_1(17483) <= 4353734;
srom_1(17484) <= 3859863;
srom_1(17485) <= 3387229;
srom_1(17486) <= 2938048;
srom_1(17487) <= 2514427;
srom_1(17488) <= 2118352;
srom_1(17489) <= 1751680;
srom_1(17490) <= 1416131;
srom_1(17491) <= 1113278;
srom_1(17492) <= 844542;
srom_1(17493) <= 611183;
srom_1(17494) <= 414294;
srom_1(17495) <= 254800;
srom_1(17496) <= 133448;
srom_1(17497) <= 50808;
srom_1(17498) <= 7266;
srom_1(17499) <= 3027;
srom_1(17500) <= 38111;
srom_1(17501) <= 112353;
srom_1(17502) <= 225406;
srom_1(17503) <= 376738;
srom_1(17504) <= 565641;
srom_1(17505) <= 791229;
srom_1(17506) <= 1052443;
srom_1(17507) <= 1348059;
srom_1(17508) <= 1676691;
srom_1(17509) <= 2036797;
srom_1(17510) <= 2426689;
srom_1(17511) <= 2844538;
srom_1(17512) <= 3288386;
srom_1(17513) <= 3756150;
srom_1(17514) <= 4245637;
srom_1(17515) <= 4754552;
srom_1(17516) <= 5280509;
srom_1(17517) <= 5821040;
srom_1(17518) <= 6373612;
srom_1(17519) <= 6935632;
srom_1(17520) <= 7504467;
srom_1(17521) <= 8077447;
srom_1(17522) <= 8651886;
srom_1(17523) <= 9225091;
srom_1(17524) <= 9794373;
srom_1(17525) <= 10357063;
srom_1(17526) <= 10910522;
srom_1(17527) <= 11452155;
srom_1(17528) <= 11979422;
srom_1(17529) <= 12489850;
srom_1(17530) <= 12981047;
srom_1(17531) <= 13450707;
srom_1(17532) <= 13896630;
srom_1(17533) <= 14316724;
srom_1(17534) <= 14709019;
srom_1(17535) <= 15071675;
srom_1(17536) <= 15402992;
srom_1(17537) <= 15701417;
srom_1(17538) <= 15965549;
srom_1(17539) <= 16194150;
srom_1(17540) <= 16386148;
srom_1(17541) <= 16540643;
srom_1(17542) <= 16656910;
srom_1(17543) <= 16734404;
srom_1(17544) <= 16772762;
srom_1(17545) <= 16771804;
srom_1(17546) <= 16731534;
srom_1(17547) <= 16652142;
srom_1(17548) <= 16533998;
srom_1(17549) <= 16377659;
srom_1(17550) <= 16183855;
srom_1(17551) <= 15953498;
srom_1(17552) <= 15687665;
srom_1(17553) <= 15387605;
srom_1(17554) <= 15054725;
srom_1(17555) <= 14690584;
srom_1(17556) <= 14296892;
srom_1(17557) <= 13875493;
srom_1(17558) <= 13428365;
srom_1(17559) <= 12957603;
srom_1(17560) <= 12465416;
srom_1(17561) <= 11954111;
srom_1(17562) <= 11426087;
srom_1(17563) <= 10883818;
srom_1(17564) <= 10329849;
srom_1(17565) <= 9766776;
srom_1(17566) <= 9197241;
srom_1(17567) <= 8623914;
srom_1(17568) <= 8049484;
srom_1(17569) <= 7476643;
srom_1(17570) <= 6908079;
srom_1(17571) <= 6346458;
srom_1(17572) <= 5794414;
srom_1(17573) <= 5254534;
srom_1(17574) <= 4729351;
srom_1(17575) <= 4221327;
srom_1(17576) <= 3732846;
srom_1(17577) <= 3266197;
srom_1(17578) <= 2823568;
srom_1(17579) <= 2407036;
srom_1(17580) <= 2018554;
srom_1(17581) <= 1659943;
srom_1(17582) <= 1332885;
srom_1(17583) <= 1038913;
srom_1(17584) <= 779407;
srom_1(17585) <= 555583;
srom_1(17586) <= 368491;
srom_1(17587) <= 219008;
srom_1(17588) <= 107835;
srom_1(17589) <= 35493;
srom_1(17590) <= 2322;
srom_1(17591) <= 8477;
srom_1(17592) <= 53929;
srom_1(17593) <= 138466;
srom_1(17594) <= 261690;
srom_1(17595) <= 423024;
srom_1(17596) <= 621712;
srom_1(17597) <= 856821;
srom_1(17598) <= 1127249;
srom_1(17599) <= 1431729;
srom_1(17600) <= 1768831;
srom_1(17601) <= 2136976;
srom_1(17602) <= 2534437;
srom_1(17603) <= 2959350;
srom_1(17604) <= 3409723;
srom_1(17605) <= 3883444;
srom_1(17606) <= 4378290;
srom_1(17607) <= 4891943;
srom_1(17608) <= 5421992;
srom_1(17609) <= 5965953;
srom_1(17610) <= 6521275;
srom_1(17611) <= 7085353;
srom_1(17612) <= 7655543;
srom_1(17613) <= 8229170;
srom_1(17614) <= 8803545;
srom_1(17615) <= 9375974;
srom_1(17616) <= 9943773;
srom_1(17617) <= 10504280;
srom_1(17618) <= 11054865;
srom_1(17619) <= 11592947;
srom_1(17620) <= 12116003;
srom_1(17621) <= 12621580;
srom_1(17622) <= 13107307;
srom_1(17623) <= 13570906;
srom_1(17624) <= 14010204;
srom_1(17625) <= 14423140;
srom_1(17626) <= 14807778;
srom_1(17627) <= 15162315;
srom_1(17628) <= 15485087;
srom_1(17629) <= 15774582;
srom_1(17630) <= 16029441;
srom_1(17631) <= 16248469;
srom_1(17632) <= 16430640;
srom_1(17633) <= 16575099;
srom_1(17634) <= 16681169;
srom_1(17635) <= 16748352;
srom_1(17636) <= 16776334;
srom_1(17637) <= 16764982;
srom_1(17638) <= 16714351;
srom_1(17639) <= 16624677;
srom_1(17640) <= 16496382;
srom_1(17641) <= 16330067;
srom_1(17642) <= 16126511;
srom_1(17643) <= 15886670;
srom_1(17644) <= 15611668;
srom_1(17645) <= 15302794;
srom_1(17646) <= 14961497;
srom_1(17647) <= 14589378;
srom_1(17648) <= 14188181;
srom_1(17649) <= 13759788;
srom_1(17650) <= 13306208;
srom_1(17651) <= 12829567;
srom_1(17652) <= 12332101;
srom_1(17653) <= 11816143;
srom_1(17654) <= 11284112;
srom_1(17655) <= 10738503;
srom_1(17656) <= 10181874;
srom_1(17657) <= 9616836;
srom_1(17658) <= 9046039;
srom_1(17659) <= 8472158;
srom_1(17660) <= 7897886;
srom_1(17661) <= 7325915;
srom_1(17662) <= 6758927;
srom_1(17663) <= 6199582;
srom_1(17664) <= 5650501;
srom_1(17665) <= 5114261;
srom_1(17666) <= 4593375;
srom_1(17667) <= 4090286;
srom_1(17668) <= 3607353;
srom_1(17669) <= 3146841;
srom_1(17670) <= 2710910;
srom_1(17671) <= 2301604;
srom_1(17672) <= 1920841;
srom_1(17673) <= 1570408;
srom_1(17674) <= 1251948;
srom_1(17675) <= 966954;
srom_1(17676) <= 716763;
srom_1(17677) <= 502548;
srom_1(17678) <= 325313;
srom_1(17679) <= 185890;
srom_1(17680) <= 84932;
srom_1(17681) <= 22913;
srom_1(17682) <= 123;
srom_1(17683) <= 16670;
srom_1(17684) <= 72476;
srom_1(17685) <= 167279;
srom_1(17686) <= 300635;
srom_1(17687) <= 471918;
srom_1(17688) <= 680325;
srom_1(17689) <= 924879;
srom_1(17690) <= 1204433;
srom_1(17691) <= 1517676;
srom_1(17692) <= 1863139;
srom_1(17693) <= 2239202;
srom_1(17694) <= 2644102;
srom_1(17695) <= 3075939;
srom_1(17696) <= 3532690;
srom_1(17697) <= 4012212;
srom_1(17698) <= 4512256;
srom_1(17699) <= 5030478;
srom_1(17700) <= 5564447;
srom_1(17701) <= 6111660;
srom_1(17702) <= 6669550;
srom_1(17703) <= 7235501;
srom_1(17704) <= 7806860;
srom_1(17705) <= 8380946;
srom_1(17706) <= 8955069;
srom_1(17707) <= 9526535;
srom_1(17708) <= 10092665;
srom_1(17709) <= 10650804;
srom_1(17710) <= 11198335;
srom_1(17711) <= 11732690;
srom_1(17712) <= 12251363;
srom_1(17713) <= 12751923;
srom_1(17714) <= 13232022;
srom_1(17715) <= 13689408;
srom_1(17716) <= 14121937;
srom_1(17717) <= 14527580;
srom_1(17718) <= 14904436;
srom_1(17719) <= 15250737;
srom_1(17720) <= 15564858;
srom_1(17721) <= 15845328;
srom_1(17722) <= 16090831;
srom_1(17723) <= 16300215;
srom_1(17724) <= 16472500;
srom_1(17725) <= 16606876;
srom_1(17726) <= 16702713;
srom_1(17727) <= 16759563;
srom_1(17728) <= 16777159;
srom_1(17729) <= 16755418;
srom_1(17730) <= 16694442;
srom_1(17731) <= 16594517;
srom_1(17732) <= 16456112;
srom_1(17733) <= 16279875;
srom_1(17734) <= 16066634;
srom_1(17735) <= 15817387;
srom_1(17736) <= 15533305;
srom_1(17737) <= 15215719;
srom_1(17738) <= 14866118;
srom_1(17739) <= 14486141;
srom_1(17740) <= 14077572;
srom_1(17741) <= 13642324;
srom_1(17742) <= 13182441;
srom_1(17743) <= 12700077;
srom_1(17744) <= 12197495;
srom_1(17745) <= 11677052;
srom_1(17746) <= 11141189;
srom_1(17747) <= 10592418;
srom_1(17748) <= 10033312;
srom_1(17749) <= 9466494;
srom_1(17750) <= 8894621;
srom_1(17751) <= 8320375;
srom_1(17752) <= 7746449;
srom_1(17753) <= 7175535;
srom_1(17754) <= 6610309;
srom_1(17755) <= 6053422;
srom_1(17756) <= 5507485;
srom_1(17757) <= 4975059;
srom_1(17758) <= 4458641;
srom_1(17759) <= 3960651;
srom_1(17760) <= 3483426;
srom_1(17761) <= 3029202;
srom_1(17762) <= 2600111;
srom_1(17763) <= 2198164;
srom_1(17764) <= 1825246;
srom_1(17765) <= 1483106;
srom_1(17766) <= 1173348;
srom_1(17767) <= 897425;
srom_1(17768) <= 656631;
srom_1(17769) <= 452095;
srom_1(17770) <= 284775;
srom_1(17771) <= 155458;
srom_1(17772) <= 64748;
srom_1(17773) <= 13072;
srom_1(17774) <= 671;
srom_1(17775) <= 27605;
srom_1(17776) <= 93746;
srom_1(17777) <= 198785;
srom_1(17778) <= 342228;
srom_1(17779) <= 523404;
srom_1(17780) <= 741462;
srom_1(17781) <= 995380;
srom_1(17782) <= 1283968;
srom_1(17783) <= 1605872;
srom_1(17784) <= 1959582;
srom_1(17785) <= 2343441;
srom_1(17786) <= 2755647;
srom_1(17787) <= 3194268;
srom_1(17788) <= 3657247;
srom_1(17789) <= 4142413;
srom_1(17790) <= 4647491;
srom_1(17791) <= 5170112;
srom_1(17792) <= 5707826;
srom_1(17793) <= 6258111;
srom_1(17794) <= 6818387;
srom_1(17795) <= 7386026;
srom_1(17796) <= 7958366;
srom_1(17797) <= 8532724;
srom_1(17798) <= 9106407;
srom_1(17799) <= 9676723;
srom_1(17800) <= 10240998;
srom_1(17801) <= 10796588;
srom_1(17802) <= 11340885;
srom_1(17803) <= 11871338;
srom_1(17804) <= 12385459;
srom_1(17805) <= 12880838;
srom_1(17806) <= 13355151;
srom_1(17807) <= 13806175;
srom_1(17808) <= 14231793;
srom_1(17809) <= 14630011;
srom_1(17810) <= 14998960;
srom_1(17811) <= 15336912;
srom_1(17812) <= 15642280;
srom_1(17813) <= 15913634;
srom_1(17814) <= 16149700;
srom_1(17815) <= 16349372;
srom_1(17816) <= 16511712;
srom_1(17817) <= 16635961;
srom_1(17818) <= 16721535;
srom_1(17819) <= 16768034;
srom_1(17820) <= 16775238;
srom_1(17821) <= 16743114;
srom_1(17822) <= 16671813;
srom_1(17823) <= 16561670;
srom_1(17824) <= 16413200;
srom_1(17825) <= 16227100;
srom_1(17826) <= 16004242;
srom_1(17827) <= 15745673;
srom_1(17828) <= 15452603;
srom_1(17829) <= 15126408;
srom_1(17830) <= 14768617;
srom_1(17831) <= 14380908;
srom_1(17832) <= 13965100;
srom_1(17833) <= 13523141;
srom_1(17834) <= 13057104;
srom_1(17835) <= 12569175;
srom_1(17836) <= 12061642;
srom_1(17837) <= 11536885;
srom_1(17838) <= 10997365;
srom_1(17839) <= 10445611;
srom_1(17840) <= 9884211;
srom_1(17841) <= 9315798;
srom_1(17842) <= 8743037;
srom_1(17843) <= 8168614;
srom_1(17844) <= 7595222;
srom_1(17845) <= 7025551;
srom_1(17846) <= 6462272;
srom_1(17847) <= 5908026;
srom_1(17848) <= 5365413;
srom_1(17849) <= 4836976;
srom_1(17850) <= 4325194;
srom_1(17851) <= 3832466;
srom_1(17852) <= 3361104;
srom_1(17853) <= 2913318;
srom_1(17854) <= 2491207;
srom_1(17855) <= 2096751;
srom_1(17856) <= 1731800;
srom_1(17857) <= 1398065;
srom_1(17858) <= 1097111;
srom_1(17859) <= 830349;
srom_1(17860) <= 599030;
srom_1(17861) <= 404240;
srom_1(17862) <= 246891;
srom_1(17863) <= 127721;
srom_1(17864) <= 47289;
srom_1(17865) <= 5973;
srom_1(17866) <= 3966;
srom_1(17867) <= 41277;
srom_1(17868) <= 117731;
srom_1(17869) <= 232971;
srom_1(17870) <= 386455;
srom_1(17871) <= 577464;
srom_1(17872) <= 805102;
srom_1(17873) <= 1068302;
srom_1(17874) <= 1365830;
srom_1(17875) <= 1696289;
srom_1(17876) <= 2058131;
srom_1(17877) <= 2449659;
srom_1(17878) <= 2869036;
srom_1(17879) <= 3314297;
srom_1(17880) <= 3783353;
srom_1(17881) <= 4274005;
srom_1(17882) <= 4783951;
srom_1(17883) <= 5310801;
srom_1(17884) <= 5852083;
srom_1(17885) <= 6405261;
srom_1(17886) <= 6967739;
srom_1(17887) <= 7536879;
srom_1(17888) <= 8110014;
srom_1(17889) <= 8684456;
srom_1(17890) <= 9257510;
srom_1(17891) <= 9826489;
srom_1(17892) <= 10388726;
srom_1(17893) <= 10941583;
srom_1(17894) <= 11482469;
srom_1(17895) <= 12008846;
srom_1(17896) <= 12518247;
srom_1(17897) <= 13008282;
srom_1(17898) <= 13476655;
srom_1(17899) <= 13921167;
srom_1(17900) <= 14339736;
srom_1(17901) <= 14730398;
srom_1(17902) <= 15091321;
srom_1(17903) <= 15420812;
srom_1(17904) <= 15717328;
srom_1(17905) <= 15979476;
srom_1(17906) <= 16206028;
srom_1(17907) <= 16395921;
srom_1(17908) <= 16548266;
srom_1(17909) <= 16662347;
srom_1(17910) <= 16737629;
srom_1(17911) <= 16773761;
srom_1(17912) <= 16770571;
srom_1(17913) <= 16728075;
srom_1(17914) <= 16646473;
srom_1(17915) <= 16526147;
srom_1(17916) <= 16367661;
srom_1(17917) <= 16171758;
srom_1(17918) <= 15939358;
srom_1(17919) <= 15671549;
srom_1(17920) <= 15369589;
srom_1(17921) <= 15034892;
srom_1(17922) <= 14669028;
srom_1(17923) <= 14273714;
srom_1(17924) <= 13850802;
srom_1(17925) <= 13402276;
srom_1(17926) <= 12930239;
srom_1(17927) <= 12436905;
srom_1(17928) <= 11924587;
srom_1(17929) <= 11395687;
srom_1(17930) <= 10852687;
srom_1(17931) <= 10298131;
srom_1(17932) <= 9734621;
srom_1(17933) <= 9164799;
srom_1(17934) <= 8591337;
srom_1(17935) <= 8016925;
srom_1(17936) <= 7444256;
srom_1(17937) <= 6876014;
srom_1(17938) <= 6314866;
srom_1(17939) <= 5763443;
srom_1(17940) <= 5224330;
srom_1(17941) <= 4700055;
srom_1(17942) <= 4193077;
srom_1(17943) <= 3705773;
srom_1(17944) <= 3240429;
srom_1(17945) <= 2799226;
srom_1(17946) <= 2384234;
srom_1(17947) <= 1997398;
srom_1(17948) <= 1640533;
srom_1(17949) <= 1315312;
srom_1(17950) <= 1023260;
srom_1(17951) <= 765747;
srom_1(17952) <= 543980;
srom_1(17953) <= 358999;
srom_1(17954) <= 211672;
srom_1(17955) <= 102689;
srom_1(17956) <= 32561;
srom_1(17957) <= 1618;
srom_1(17958) <= 10005;
srom_1(17959) <= 57681;
srom_1(17960) <= 144425;
srom_1(17961) <= 269828;
srom_1(17962) <= 433302;
srom_1(17963) <= 634082;
srom_1(17964) <= 871226;
srom_1(17965) <= 1143621;
srom_1(17966) <= 1449990;
srom_1(17967) <= 1788897;
srom_1(17968) <= 2158752;
srom_1(17969) <= 2557821;
srom_1(17970) <= 2984233;
srom_1(17971) <= 3435988;
srom_1(17972) <= 3910967;
srom_1(17973) <= 4406943;
srom_1(17974) <= 4921591;
srom_1(17975) <= 5452497;
srom_1(17976) <= 5997171;
srom_1(17977) <= 6553059;
srom_1(17978) <= 7117555;
srom_1(17979) <= 7688012;
srom_1(17980) <= 8261753;
srom_1(17981) <= 8836090;
srom_1(17982) <= 9408328;
srom_1(17983) <= 9975784;
srom_1(17984) <= 10535798;
srom_1(17985) <= 11085742;
srom_1(17986) <= 11623039;
srom_1(17987) <= 12145169;
srom_1(17988) <= 12649682;
srom_1(17989) <= 13134214;
srom_1(17990) <= 13596492;
srom_1(17991) <= 14034349;
srom_1(17992) <= 14445731;
srom_1(17993) <= 14828709;
srom_1(17994) <= 15181487;
srom_1(17995) <= 15502411;
srom_1(17996) <= 15789975;
srom_1(17997) <= 16042833;
srom_1(17998) <= 16259796;
srom_1(17999) <= 16439850;
srom_1(18000) <= 16582148;
srom_1(18001) <= 16686024;
srom_1(18002) <= 16750990;
srom_1(18003) <= 16776742;
srom_1(18004) <= 16763160;
srom_1(18005) <= 16710306;
srom_1(18006) <= 16618429;
srom_1(18007) <= 16487960;
srom_1(18008) <= 16319509;
srom_1(18009) <= 16113869;
srom_1(18010) <= 15872001;
srom_1(18011) <= 15595042;
srom_1(18012) <= 15284289;
srom_1(18013) <= 14941200;
srom_1(18014) <= 14567383;
srom_1(18015) <= 14164592;
srom_1(18016) <= 13734716;
srom_1(18017) <= 13279770;
srom_1(18018) <= 12801887;
srom_1(18019) <= 12303309;
srom_1(18020) <= 11786374;
srom_1(18021) <= 11253505;
srom_1(18022) <= 10707202;
srom_1(18023) <= 10150026;
srom_1(18024) <= 9584590;
srom_1(18025) <= 9013546;
srom_1(18026) <= 8439571;
srom_1(18027) <= 7865358;
srom_1(18028) <= 7293598;
srom_1(18029) <= 6726973;
srom_1(18030) <= 6168140;
srom_1(18031) <= 5619719;
srom_1(18032) <= 5084283;
srom_1(18033) <= 4564341;
srom_1(18034) <= 4062333;
srom_1(18035) <= 3580613;
srom_1(18036) <= 3121439;
srom_1(18037) <= 2686964;
srom_1(18038) <= 2279226;
srom_1(18039) <= 1900138;
srom_1(18040) <= 1551476;
srom_1(18041) <= 1234875;
srom_1(18042) <= 951821;
srom_1(18043) <= 703641;
srom_1(18044) <= 491498;
srom_1(18045) <= 316387;
srom_1(18046) <= 179129;
srom_1(18047) <= 80369;
srom_1(18048) <= 20569;
srom_1(18049) <= 10;
srom_1(18050) <= 18787;
srom_1(18051) <= 76814;
srom_1(18052) <= 173817;
srom_1(18053) <= 309342;
srom_1(18054) <= 482754;
srom_1(18055) <= 693239;
srom_1(18056) <= 939810;
srom_1(18057) <= 1221311;
srom_1(18058) <= 1536422;
srom_1(18059) <= 1883666;
srom_1(18060) <= 2261413;
srom_1(18061) <= 2667893;
srom_1(18062) <= 3101199;
srom_1(18063) <= 3559300;
srom_1(18064) <= 4040046;
srom_1(18065) <= 4541185;
srom_1(18066) <= 5060366;
srom_1(18067) <= 5595154;
srom_1(18068) <= 6143041;
srom_1(18069) <= 6701459;
srom_1(18070) <= 7267788;
srom_1(18071) <= 7839373;
srom_1(18072) <= 8413534;
srom_1(18073) <= 8987578;
srom_1(18074) <= 9558813;
srom_1(18075) <= 10124560;
srom_1(18076) <= 10682167;
srom_1(18077) <= 11229019;
srom_1(18078) <= 11762551;
srom_1(18079) <= 12280261;
srom_1(18080) <= 12779723;
srom_1(18081) <= 13258592;
srom_1(18082) <= 13714625;
srom_1(18083) <= 14145682;
srom_1(18084) <= 14549742;
srom_1(18085) <= 14924911;
srom_1(18086) <= 15269429;
srom_1(18087) <= 15581680;
srom_1(18088) <= 15860200;
srom_1(18089) <= 16103683;
srom_1(18090) <= 16310988;
srom_1(18091) <= 16481142;
srom_1(18092) <= 16613347;
srom_1(18093) <= 16706984;
srom_1(18094) <= 16761613;
srom_1(18095) <= 16776978;
srom_1(18096) <= 16753007;
srom_1(18097) <= 16689812;
srom_1(18098) <= 16587691;
srom_1(18099) <= 16447121;
srom_1(18100) <= 16268762;
srom_1(18101) <= 16053450;
srom_1(18102) <= 15802195;
srom_1(18103) <= 15516175;
srom_1(18104) <= 15196731;
srom_1(18105) <= 14845362;
srom_1(18106) <= 14463715;
srom_1(18107) <= 14053580;
srom_1(18108) <= 13616880;
srom_1(18109) <= 13155662;
srom_1(18110) <= 12672090;
srom_1(18111) <= 12168432;
srom_1(18112) <= 11647048;
srom_1(18113) <= 11110385;
srom_1(18114) <= 10560958;
srom_1(18115) <= 10001344;
srom_1(18116) <= 9434168;
srom_1(18117) <= 8862088;
srom_1(18118) <= 8287789;
srom_1(18119) <= 7713962;
srom_1(18120) <= 7143299;
srom_1(18121) <= 6578475;
srom_1(18122) <= 6022140;
srom_1(18123) <= 5476902;
srom_1(18124) <= 4945317;
srom_1(18125) <= 4429880;
srom_1(18126) <= 3933007;
srom_1(18127) <= 3457027;
srom_1(18128) <= 3004173;
srom_1(18129) <= 2576569;
srom_1(18130) <= 2176219;
srom_1(18131) <= 1805001;
srom_1(18132) <= 1464656;
srom_1(18133) <= 1156780;
srom_1(18134) <= 882817;
srom_1(18135) <= 644050;
srom_1(18136) <= 441601;
srom_1(18137) <= 276418;
srom_1(18138) <= 149275;
srom_1(18139) <= 60770;
srom_1(18140) <= 11317;
srom_1(18141) <= 1147;
srom_1(18142) <= 30310;
srom_1(18143) <= 98667;
srom_1(18144) <= 205899;
srom_1(18145) <= 351502;
srom_1(18146) <= 534794;
srom_1(18147) <= 754915;
srom_1(18148) <= 1010833;
srom_1(18149) <= 1301348;
srom_1(18150) <= 1625098;
srom_1(18151) <= 1980564;
srom_1(18152) <= 2366080;
srom_1(18153) <= 2779837;
srom_1(18154) <= 3219896;
srom_1(18155) <= 3684193;
srom_1(18156) <= 4170550;
srom_1(18157) <= 4676687;
srom_1(18158) <= 5200231;
srom_1(18159) <= 5738726;
srom_1(18160) <= 6289647;
srom_1(18161) <= 6850411;
srom_1(18162) <= 7418388;
srom_1(18163) <= 7990915;
srom_1(18164) <= 8565306;
srom_1(18165) <= 9138869;
srom_1(18166) <= 9708914;
srom_1(18167) <= 10272768;
srom_1(18168) <= 10827786;
srom_1(18169) <= 11371366;
srom_1(18170) <= 11900958;
srom_1(18171) <= 12414080;
srom_1(18172) <= 12908325;
srom_1(18173) <= 13381376;
srom_1(18174) <= 13831014;
srom_1(18175) <= 14255131;
srom_1(18176) <= 14651737;
srom_1(18177) <= 15018973;
srom_1(18178) <= 15355118;
srom_1(18179) <= 15658594;
srom_1(18180) <= 15927978;
srom_1(18181) <= 16162008;
srom_1(18182) <= 16359586;
srom_1(18183) <= 16519785;
srom_1(18184) <= 16641854;
srom_1(18185) <= 16725221;
srom_1(18186) <= 16769494;
srom_1(18187) <= 16774467;
srom_1(18188) <= 16740116;
srom_1(18189) <= 16666601;
srom_1(18190) <= 16554268;
srom_1(18191) <= 16403644;
srom_1(18192) <= 16215434;
srom_1(18193) <= 15990521;
srom_1(18194) <= 15729961;
srom_1(18195) <= 15434974;
srom_1(18196) <= 15106945;
srom_1(18197) <= 14747411;
srom_1(18198) <= 14358058;
srom_1(18199) <= 13940713;
srom_1(18200) <= 13497332;
srom_1(18201) <= 13029994;
srom_1(18202) <= 12540891;
srom_1(18203) <= 12032317;
srom_1(18204) <= 11506656;
srom_1(18205) <= 10966373;
srom_1(18206) <= 10414003;
srom_1(18207) <= 9852134;
srom_1(18208) <= 9283403;
srom_1(18209) <= 8710476;
srom_1(18210) <= 8136039;
srom_1(18211) <= 7562787;
srom_1(18212) <= 6993407;
srom_1(18213) <= 6430570;
srom_1(18214) <= 5876915;
srom_1(18215) <= 5335037;
srom_1(18216) <= 4807480;
srom_1(18217) <= 4296715;
srom_1(18218) <= 3805138;
srom_1(18219) <= 3335055;
srom_1(18220) <= 2888670;
srom_1(18221) <= 2468076;
srom_1(18222) <= 2075246;
srom_1(18223) <= 1712020;
srom_1(18224) <= 1380104;
srom_1(18225) <= 1081053;
srom_1(18226) <= 816270;
srom_1(18227) <= 586996;
srom_1(18228) <= 394306;
srom_1(18229) <= 239104;
srom_1(18230) <= 122118;
srom_1(18231) <= 43897;
srom_1(18232) <= 4807;
srom_1(18233) <= 5031;
srom_1(18234) <= 44569;
srom_1(18235) <= 123234;
srom_1(18236) <= 240659;
srom_1(18237) <= 396293;
srom_1(18238) <= 589405;
srom_1(18239) <= 819090;
srom_1(18240) <= 1084272;
srom_1(18241) <= 1383706;
srom_1(18242) <= 1715988;
srom_1(18243) <= 2079560;
srom_1(18244) <= 2472718;
srom_1(18245) <= 2893618;
srom_1(18246) <= 3340285;
srom_1(18247) <= 3810626;
srom_1(18248) <= 4302434;
srom_1(18249) <= 4813404;
srom_1(18250) <= 5341139;
srom_1(18251) <= 5883165;
srom_1(18252) <= 6436940;
srom_1(18253) <= 6999866;
srom_1(18254) <= 7569305;
srom_1(18255) <= 8142586;
srom_1(18256) <= 8717021;
srom_1(18257) <= 9289915;
srom_1(18258) <= 9858584;
srom_1(18259) <= 10420358;
srom_1(18260) <= 10972606;
srom_1(18261) <= 11512736;
srom_1(18262) <= 12038215;
srom_1(18263) <= 12546581;
srom_1(18264) <= 13035448;
srom_1(18265) <= 13502525;
srom_1(18266) <= 13945621;
srom_1(18267) <= 14362658;
srom_1(18268) <= 14751681;
srom_1(18269) <= 15110865;
srom_1(18270) <= 15438526;
srom_1(18271) <= 15733128;
srom_1(18272) <= 15993288;
srom_1(18273) <= 16217788;
srom_1(18274) <= 16405574;
srom_1(18275) <= 16555766;
srom_1(18276) <= 16667659;
srom_1(18277) <= 16740728;
srom_1(18278) <= 16774632;
srom_1(18279) <= 16769211;
srom_1(18280) <= 16724490;
srom_1(18281) <= 16640680;
srom_1(18282) <= 16518172;
srom_1(18283) <= 16357543;
srom_1(18284) <= 16159544;
srom_1(18285) <= 15925104;
srom_1(18286) <= 15655324;
srom_1(18287) <= 15351467;
srom_1(18288) <= 15014959;
srom_1(18289) <= 14647378;
srom_1(18290) <= 14250447;
srom_1(18291) <= 13826028;
srom_1(18292) <= 13376111;
srom_1(18293) <= 12902806;
srom_1(18294) <= 12408332;
srom_1(18295) <= 11895009;
srom_1(18296) <= 11365243;
srom_1(18297) <= 10821518;
srom_1(18298) <= 10266385;
srom_1(18299) <= 9702445;
srom_1(18300) <= 9132345;
srom_1(18301) <= 8558758;
srom_1(18302) <= 7984372;
srom_1(18303) <= 7411882;
srom_1(18304) <= 6843972;
srom_1(18305) <= 6283306;
srom_1(18306) <= 5732512;
srom_1(18307) <= 5194173;
srom_1(18308) <= 4670814;
srom_1(18309) <= 4164889;
srom_1(18310) <= 3678771;
srom_1(18311) <= 3214739;
srom_1(18312) <= 2774968;
srom_1(18313) <= 2361522;
srom_1(18314) <= 1976339;
srom_1(18315) <= 1621225;
srom_1(18316) <= 1297846;
srom_1(18317) <= 1007718;
srom_1(18318) <= 752202;
srom_1(18319) <= 532495;
srom_1(18320) <= 349628;
srom_1(18321) <= 204459;
srom_1(18322) <= 97668;
srom_1(18323) <= 29756;
srom_1(18324) <= 1041;
srom_1(18325) <= 11659;
srom_1(18326) <= 61559;
srom_1(18327) <= 150508;
srom_1(18328) <= 278088;
srom_1(18329) <= 443700;
srom_1(18330) <= 646570;
srom_1(18331) <= 885744;
srom_1(18332) <= 1160102;
srom_1(18333) <= 1468356;
srom_1(18334) <= 1809062;
srom_1(18335) <= 2180622;
srom_1(18336) <= 2581294;
srom_1(18337) <= 3009197;
srom_1(18338) <= 3462327;
srom_1(18339) <= 3938558;
srom_1(18340) <= 4435656;
srom_1(18341) <= 4951291;
srom_1(18342) <= 5483045;
srom_1(18343) <= 6028424;
srom_1(18344) <= 6584871;
srom_1(18345) <= 7149776;
srom_1(18346) <= 7720491;
srom_1(18347) <= 8294338;
srom_1(18348) <= 8868628;
srom_1(18349) <= 9440666;
srom_1(18350) <= 10007772;
srom_1(18351) <= 10567284;
srom_1(18352) <= 11116579;
srom_1(18353) <= 11653083;
srom_1(18354) <= 12174278;
srom_1(18355) <= 12677721;
srom_1(18356) <= 13161050;
srom_1(18357) <= 13622000;
srom_1(18358) <= 14058409;
srom_1(18359) <= 14468230;
srom_1(18360) <= 14849542;
srom_1(18361) <= 15200556;
srom_1(18362) <= 15519627;
srom_1(18363) <= 15805257;
srom_1(18364) <= 16056109;
srom_1(18365) <= 16271005;
srom_1(18366) <= 16448938;
srom_1(18367) <= 16589073;
srom_1(18368) <= 16690753;
srom_1(18369) <= 16753502;
srom_1(18370) <= 16777024;
srom_1(18371) <= 16761211;
srom_1(18372) <= 16706136;
srom_1(18373) <= 16612056;
srom_1(18374) <= 16479415;
srom_1(18375) <= 16308832;
srom_1(18376) <= 16101109;
srom_1(18377) <= 15857220;
srom_1(18378) <= 15578307;
srom_1(18379) <= 15265680;
srom_1(18380) <= 14920804;
srom_1(18381) <= 14545295;
srom_1(18382) <= 14140917;
srom_1(18383) <= 13709563;
srom_1(18384) <= 13253258;
srom_1(18385) <= 12774140;
srom_1(18386) <= 12274458;
srom_1(18387) <= 11756553;
srom_1(18388) <= 11222855;
srom_1(18389) <= 10675866;
srom_1(18390) <= 10118151;
srom_1(18391) <= 9552326;
srom_1(18392) <= 8981044;
srom_1(18393) <= 8406984;
srom_1(18394) <= 7832837;
srom_1(18395) <= 7261297;
srom_1(18396) <= 6695043;
srom_1(18397) <= 6136731;
srom_1(18398) <= 5588979;
srom_1(18399) <= 5054355;
srom_1(18400) <= 4535366;
srom_1(18401) <= 4034447;
srom_1(18402) <= 3553945;
srom_1(18403) <= 3096115;
srom_1(18404) <= 2663104;
srom_1(18405) <= 2256941;
srom_1(18406) <= 1879532;
srom_1(18407) <= 1532646;
srom_1(18408) <= 1217910;
srom_1(18409) <= 936800;
srom_1(18410) <= 690634;
srom_1(18411) <= 480566;
srom_1(18412) <= 307582;
srom_1(18413) <= 172493;
srom_1(18414) <= 75932;
srom_1(18415) <= 18352;
srom_1(18416) <= 22;
srom_1(18417) <= 21030;
srom_1(18418) <= 81276;
srom_1(18419) <= 180478;
srom_1(18420) <= 318171;
srom_1(18421) <= 493709;
srom_1(18422) <= 706269;
srom_1(18423) <= 954854;
srom_1(18424) <= 1238298;
srom_1(18425) <= 1555273;
srom_1(18426) <= 1904291;
srom_1(18427) <= 2283717;
srom_1(18428) <= 2691770;
srom_1(18429) <= 3126538;
srom_1(18430) <= 3585982;
srom_1(18431) <= 4067946;
srom_1(18432) <= 4570172;
srom_1(18433) <= 5090304;
srom_1(18434) <= 5625903;
srom_1(18435) <= 6174457;
srom_1(18436) <= 6733393;
srom_1(18437) <= 7300092;
srom_1(18438) <= 7871895;
srom_1(18439) <= 8446121;
srom_1(18440) <= 9020078;
srom_1(18441) <= 9591073;
srom_1(18442) <= 10156429;
srom_1(18443) <= 10713496;
srom_1(18444) <= 11259660;
srom_1(18445) <= 11792361;
srom_1(18446) <= 12309101;
srom_1(18447) <= 12807456;
srom_1(18448) <= 13285089;
srom_1(18449) <= 13739762;
srom_1(18450) <= 14169341;
srom_1(18451) <= 14571812;
srom_1(18452) <= 14945287;
srom_1(18453) <= 15288017;
srom_1(18454) <= 15598392;
srom_1(18455) <= 15874959;
srom_1(18456) <= 16116419;
srom_1(18457) <= 16321641;
srom_1(18458) <= 16489662;
srom_1(18459) <= 16619695;
srom_1(18460) <= 16711129;
srom_1(18461) <= 16763536;
srom_1(18462) <= 16776670;
srom_1(18463) <= 16750470;
srom_1(18464) <= 16685058;
srom_1(18465) <= 16580741;
srom_1(18466) <= 16438008;
srom_1(18467) <= 16257529;
srom_1(18468) <= 16040150;
srom_1(18469) <= 15786890;
srom_1(18470) <= 15498937;
srom_1(18471) <= 15177641;
srom_1(18472) <= 14824510;
srom_1(18473) <= 14441198;
srom_1(18474) <= 14029503;
srom_1(18475) <= 13591356;
srom_1(18476) <= 13128812;
srom_1(18477) <= 12644039;
srom_1(18478) <= 12139311;
srom_1(18479) <= 11616995;
srom_1(18480) <= 11079539;
srom_1(18481) <= 10529465;
srom_1(18482) <= 9969352;
srom_1(18483) <= 9401826;
srom_1(18484) <= 8829549;
srom_1(18485) <= 8255204;
srom_1(18486) <= 7681485;
srom_1(18487) <= 7111081;
srom_1(18488) <= 6546669;
srom_1(18489) <= 5990893;
srom_1(18490) <= 5446362;
srom_1(18491) <= 4915628;
srom_1(18492) <= 4401179;
srom_1(18493) <= 3905429;
srom_1(18494) <= 3430703;
srom_1(18495) <= 2979225;
srom_1(18496) <= 2553114;
srom_1(18497) <= 2154368;
srom_1(18498) <= 1784856;
srom_1(18499) <= 1446311;
srom_1(18500) <= 1140321;
srom_1(18501) <= 868321;
srom_1(18502) <= 631586;
srom_1(18503) <= 431227;
srom_1(18504) <= 268182;
srom_1(18505) <= 143217;
srom_1(18506) <= 56917;
srom_1(18507) <= 9688;
srom_1(18508) <= 1750;
srom_1(18509) <= 33140;
srom_1(18510) <= 103713;
srom_1(18511) <= 213136;
srom_1(18512) <= 360897;
srom_1(18513) <= 546303;
srom_1(18514) <= 768483;
srom_1(18515) <= 1026397;
srom_1(18516) <= 1318835;
srom_1(18517) <= 1644426;
srom_1(18518) <= 2001643;
srom_1(18519) <= 2388810;
srom_1(18520) <= 2804112;
srom_1(18521) <= 3245602;
srom_1(18522) <= 3711209;
srom_1(18523) <= 4198750;
srom_1(18524) <= 4705939;
srom_1(18525) <= 5230397;
srom_1(18526) <= 5769665;
srom_1(18527) <= 6321214;
srom_1(18528) <= 6882458;
srom_1(18529) <= 7450764;
srom_1(18530) <= 8023469;
srom_1(18531) <= 8597885;
srom_1(18532) <= 9171321;
srom_1(18533) <= 9741086;
srom_1(18534) <= 10304509;
srom_1(18535) <= 10858947;
srom_1(18536) <= 11401801;
srom_1(18537) <= 11930525;
srom_1(18538) <= 12442640;
srom_1(18539) <= 12935745;
srom_1(18540) <= 13407526;
srom_1(18541) <= 13855771;
srom_1(18542) <= 14278380;
srom_1(18543) <= 14673369;
srom_1(18544) <= 15038886;
srom_1(18545) <= 15373219;
srom_1(18546) <= 15674798;
srom_1(18547) <= 15942209;
srom_1(18548) <= 16174199;
srom_1(18549) <= 16369680;
srom_1(18550) <= 16527735;
srom_1(18551) <= 16647622;
srom_1(18552) <= 16728781;
srom_1(18553) <= 16770829;
srom_1(18554) <= 16773570;
srom_1(18555) <= 16736991;
srom_1(18556) <= 16661264;
srom_1(18557) <= 16546743;
srom_1(18558) <= 16393967;
srom_1(18559) <= 16203650;
srom_1(18560) <= 15976686;
srom_1(18561) <= 15714138;
srom_1(18562) <= 15417239;
srom_1(18563) <= 15087380;
srom_1(18564) <= 14726109;
srom_1(18565) <= 14335118;
srom_1(18566) <= 13916242;
srom_1(18567) <= 13471446;
srom_1(18568) <= 13002814;
srom_1(18569) <= 12512544;
srom_1(18570) <= 12002936;
srom_1(18571) <= 11476379;
srom_1(18572) <= 10935343;
srom_1(18573) <= 10382364;
srom_1(18574) <= 9820035;
srom_1(18575) <= 9250995;
srom_1(18576) <= 8677910;
srom_1(18577) <= 8103468;
srom_1(18578) <= 7530364;
srom_1(18579) <= 6961284;
srom_1(18580) <= 6398897;
srom_1(18581) <= 5845841;
srom_1(18582) <= 5304709;
srom_1(18583) <= 4778038;
srom_1(18584) <= 4268298;
srom_1(18585) <= 3777880;
srom_1(18586) <= 3309083;
srom_1(18587) <= 2864106;
srom_1(18588) <= 2445035;
srom_1(18589) <= 2053835;
srom_1(18590) <= 1692342;
srom_1(18591) <= 1362249;
srom_1(18592) <= 1065106;
srom_1(18593) <= 802305;
srom_1(18594) <= 575079;
srom_1(18595) <= 384493;
srom_1(18596) <= 231441;
srom_1(18597) <= 116640;
srom_1(18598) <= 40630;
srom_1(18599) <= 3767;
srom_1(18600) <= 6223;
srom_1(18601) <= 47986;
srom_1(18602) <= 128862;
srom_1(18603) <= 248471;
srom_1(18604) <= 406251;
srom_1(18605) <= 601463;
srom_1(18606) <= 833192;
srom_1(18607) <= 1100351;
srom_1(18608) <= 1401687;
srom_1(18609) <= 1735788;
srom_1(18610) <= 2101085;
srom_1(18611) <= 2495867;
srom_1(18612) <= 2918282;
srom_1(18613) <= 3366349;
srom_1(18614) <= 3837967;
srom_1(18615) <= 4330925;
srom_1(18616) <= 4842911;
srom_1(18617) <= 5371523;
srom_1(18618) <= 5914284;
srom_1(18619) <= 6468648;
srom_1(18620) <= 7032015;
srom_1(18621) <= 7601743;
srom_1(18622) <= 8175162;
srom_1(18623) <= 8749581;
srom_1(18624) <= 9322308;
srom_1(18625) <= 9890656;
srom_1(18626) <= 10451960;
srom_1(18627) <= 11003589;
srom_1(18628) <= 11542955;
srom_1(18629) <= 12067530;
srom_1(18630) <= 12574853;
srom_1(18631) <= 13062544;
srom_1(18632) <= 13528319;
srom_1(18633) <= 13969991;
srom_1(18634) <= 14385490;
srom_1(18635) <= 14772868;
srom_1(18636) <= 15130308;
srom_1(18637) <= 15456134;
srom_1(18638) <= 15748817;
srom_1(18639) <= 16006986;
srom_1(18640) <= 16229430;
srom_1(18641) <= 16415106;
srom_1(18642) <= 16563142;
srom_1(18643) <= 16672846;
srom_1(18644) <= 16743701;
srom_1(18645) <= 16775377;
srom_1(18646) <= 16767725;
srom_1(18647) <= 16720779;
srom_1(18648) <= 16634762;
srom_1(18649) <= 16510075;
srom_1(18650) <= 16347304;
srom_1(18651) <= 16147212;
srom_1(18652) <= 15910737;
srom_1(18653) <= 15638988;
srom_1(18654) <= 15333240;
srom_1(18655) <= 14994926;
srom_1(18656) <= 14625633;
srom_1(18657) <= 14227092;
srom_1(18658) <= 13801172;
srom_1(18659) <= 13349871;
srom_1(18660) <= 12875305;
srom_1(18661) <= 12379699;
srom_1(18662) <= 11865378;
srom_1(18663) <= 11334753;
srom_1(18664) <= 10790313;
srom_1(18665) <= 10234610;
srom_1(18666) <= 9670250;
srom_1(18667) <= 9099880;
srom_1(18668) <= 8526175;
srom_1(18669) <= 7951825;
srom_1(18670) <= 7379523;
srom_1(18671) <= 6811953;
srom_1(18672) <= 6251777;
srom_1(18673) <= 5701621;
srom_1(18674) <= 5164065;
srom_1(18675) <= 4641630;
srom_1(18676) <= 4136766;
srom_1(18677) <= 3651840;
srom_1(18678) <= 3189126;
srom_1(18679) <= 2750795;
srom_1(18680) <= 2338901;
srom_1(18681) <= 1955377;
srom_1(18682) <= 1602020;
srom_1(18683) <= 1280488;
srom_1(18684) <= 992288;
srom_1(18685) <= 738772;
srom_1(18686) <= 521129;
srom_1(18687) <= 340379;
srom_1(18688) <= 197370;
srom_1(18689) <= 92772;
srom_1(18690) <= 27077;
srom_1(18691) <= 591;
srom_1(18692) <= 13440;
srom_1(18693) <= 65563;
srom_1(18694) <= 156715;
srom_1(18695) <= 286470;
srom_1(18696) <= 454218;
srom_1(18697) <= 659174;
srom_1(18698) <= 900375;
srom_1(18699) <= 1176692;
srom_1(18700) <= 1486827;
srom_1(18701) <= 1829327;
srom_1(18702) <= 2202586;
srom_1(18703) <= 2604854;
srom_1(18704) <= 3034243;
srom_1(18705) <= 3488741;
srom_1(18706) <= 3966216;
srom_1(18707) <= 4464429;
srom_1(18708) <= 4981044;
srom_1(18709) <= 5513638;
srom_1(18710) <= 6059713;
srom_1(18711) <= 6616710;
srom_1(18712) <= 7182016;
srom_1(18713) <= 7752980;
srom_1(18714) <= 8326925;
srom_1(18715) <= 8901159;
srom_1(18716) <= 9472989;
srom_1(18717) <= 10039734;
srom_1(18718) <= 10598737;
srom_1(18719) <= 11147375;
srom_1(18720) <= 11683077;
srom_1(18721) <= 12203330;
srom_1(18722) <= 12705694;
srom_1(18723) <= 13187814;
srom_1(18724) <= 13647429;
srom_1(18725) <= 14082383;
srom_1(18726) <= 14490638;
srom_1(18727) <= 14870277;
srom_1(18728) <= 15219522;
srom_1(18729) <= 15536735;
srom_1(18730) <= 15820427;
srom_1(18731) <= 16069270;
srom_1(18732) <= 16282094;
srom_1(18733) <= 16457904;
srom_1(18734) <= 16595874;
srom_1(18735) <= 16695357;
srom_1(18736) <= 16755887;
srom_1(18737) <= 16777180;
srom_1(18738) <= 16759136;
srom_1(18739) <= 16701840;
srom_1(18740) <= 16605560;
srom_1(18741) <= 16470748;
srom_1(18742) <= 16298036;
srom_1(18743) <= 16088234;
srom_1(18744) <= 15842326;
srom_1(18745) <= 15561464;
srom_1(18746) <= 15246967;
srom_1(18747) <= 14900309;
srom_1(18748) <= 14523115;
srom_1(18749) <= 14117154;
srom_1(18750) <= 13684330;
srom_1(18751) <= 13226672;
srom_1(18752) <= 12746328;
srom_1(18753) <= 12245548;
srom_1(18754) <= 11726682;
srom_1(18755) <= 11192162;
srom_1(18756) <= 10644496;
srom_1(18757) <= 10086251;
srom_1(18758) <= 9520045;
srom_1(18759) <= 8948533;
srom_1(18760) <= 8374396;
srom_1(18761) <= 7800325;
srom_1(18762) <= 7229014;
srom_1(18763) <= 6663139;
srom_1(18764) <= 6105356;
srom_1(18765) <= 5558280;
srom_1(18766) <= 5024477;
srom_1(18767) <= 4506449;
srom_1(18768) <= 4006625;
srom_1(18769) <= 3527351;
srom_1(18770) <= 3070872;
srom_1(18771) <= 2639330;
srom_1(18772) <= 2234749;
srom_1(18773) <= 1859025;
srom_1(18774) <= 1513920;
srom_1(18775) <= 1201053;
srom_1(18776) <= 921891;
srom_1(18777) <= 677744;
srom_1(18778) <= 469755;
srom_1(18779) <= 298900;
srom_1(18780) <= 165980;
srom_1(18781) <= 71620;
srom_1(18782) <= 16260;
srom_1(18783) <= 162;
srom_1(18784) <= 23399;
srom_1(18785) <= 85864;
srom_1(18786) <= 187264;
srom_1(18787) <= 327122;
srom_1(18788) <= 504783;
srom_1(18789) <= 719415;
srom_1(18790) <= 970010;
srom_1(18791) <= 1255393;
srom_1(18792) <= 1574226;
srom_1(18793) <= 1925014;
srom_1(18794) <= 2306112;
srom_1(18795) <= 2715734;
srom_1(18796) <= 3151957;
srom_1(18797) <= 3612736;
srom_1(18798) <= 4095912;
srom_1(18799) <= 4599217;
srom_1(18800) <= 5120292;
srom_1(18801) <= 5656693;
srom_1(18802) <= 6205905;
srom_1(18803) <= 6765353;
srom_1(18804) <= 7332413;
srom_1(18805) <= 7904425;
srom_1(18806) <= 8478708;
srom_1(18807) <= 9052568;
srom_1(18808) <= 9623315;
srom_1(18809) <= 10188272;
srom_1(18810) <= 10744790;
srom_1(18811) <= 11290258;
srom_1(18812) <= 11822120;
srom_1(18813) <= 12337881;
srom_1(18814) <= 12835122;
srom_1(18815) <= 13311513;
srom_1(18816) <= 13764818;
srom_1(18817) <= 14192912;
srom_1(18818) <= 14593787;
srom_1(18819) <= 14965565;
srom_1(18820) <= 15306501;
srom_1(18821) <= 15614996;
srom_1(18822) <= 15889605;
srom_1(18823) <= 16129038;
srom_1(18824) <= 16332174;
srom_1(18825) <= 16498060;
srom_1(18826) <= 16625918;
srom_1(18827) <= 16715149;
srom_1(18828) <= 16765333;
srom_1(18829) <= 16776236;
srom_1(18830) <= 16747807;
srom_1(18831) <= 16680178;
srom_1(18832) <= 16573668;
srom_1(18833) <= 16428774;
srom_1(18834) <= 16246178;
srom_1(18835) <= 16026735;
srom_1(18836) <= 15771474;
srom_1(18837) <= 15481592;
srom_1(18838) <= 15158449;
srom_1(18839) <= 14803560;
srom_1(18840) <= 14418588;
srom_1(18841) <= 14005341;
srom_1(18842) <= 13565754;
srom_1(18843) <= 13101890;
srom_1(18844) <= 12615923;
srom_1(18845) <= 12110134;
srom_1(18846) <= 11586893;
srom_1(18847) <= 11048654;
srom_1(18848) <= 10497941;
srom_1(18849) <= 9937336;
srom_1(18850) <= 9369470;
srom_1(18851) <= 8797003;
srom_1(18852) <= 8222622;
srom_1(18853) <= 7649018;
srom_1(18854) <= 7078883;
srom_1(18855) <= 6514890;
srom_1(18856) <= 5959683;
srom_1(18857) <= 5415867;
srom_1(18858) <= 4885990;
srom_1(18859) <= 4372539;
srom_1(18860) <= 3877920;
srom_1(18861) <= 3404453;
srom_1(18862) <= 2954359;
srom_1(18863) <= 2529748;
srom_1(18864) <= 2132611;
srom_1(18865) <= 1764810;
srom_1(18866) <= 1428071;
srom_1(18867) <= 1123972;
srom_1(18868) <= 853940;
srom_1(18869) <= 619240;
srom_1(18870) <= 420973;
srom_1(18871) <= 260069;
srom_1(18872) <= 137283;
srom_1(18873) <= 53190;
srom_1(18874) <= 8185;
srom_1(18875) <= 2478;
srom_1(18876) <= 36097;
srom_1(18877) <= 108884;
srom_1(18878) <= 220497;
srom_1(18879) <= 370413;
srom_1(18880) <= 557930;
srom_1(18881) <= 782167;
srom_1(18882) <= 1042073;
srom_1(18883) <= 1336429;
srom_1(18884) <= 1663856;
srom_1(18885) <= 2022817;
srom_1(18886) <= 2411630;
srom_1(18887) <= 2828471;
srom_1(18888) <= 3271385;
srom_1(18889) <= 3738296;
srom_1(18890) <= 4227013;
srom_1(18891) <= 4735246;
srom_1(18892) <= 5260611;
srom_1(18893) <= 5800643;
srom_1(18894) <= 6352812;
srom_1(18895) <= 6914527;
srom_1(18896) <= 7483155;
srom_1(18897) <= 8056028;
srom_1(18898) <= 8630462;
srom_1(18899) <= 9203761;
srom_1(18900) <= 9773237;
srom_1(18901) <= 10336221;
srom_1(18902) <= 10890071;
srom_1(18903) <= 11432191;
srom_1(18904) <= 11960039;
srom_1(18905) <= 12471139;
srom_1(18906) <= 12963095;
srom_1(18907) <= 13433599;
srom_1(18908) <= 13880446;
srom_1(18909) <= 14301540;
srom_1(18910) <= 14694905;
srom_1(18911) <= 15058699;
srom_1(18912) <= 15391214;
srom_1(18913) <= 15690891;
srom_1(18914) <= 15956326;
srom_1(18915) <= 16186273;
srom_1(18916) <= 16379654;
srom_1(18917) <= 16535562;
srom_1(18918) <= 16653266;
srom_1(18919) <= 16732214;
srom_1(18920) <= 16772037;
srom_1(18921) <= 16772546;
srom_1(18922) <= 16733741;
srom_1(18923) <= 16655802;
srom_1(18924) <= 16539096;
srom_1(18925) <= 16384169;
srom_1(18926) <= 16191748;
srom_1(18927) <= 15962735;
srom_1(18928) <= 15698205;
srom_1(18929) <= 15399398;
srom_1(18930) <= 15067714;
srom_1(18931) <= 14704710;
srom_1(18932) <= 14312088;
srom_1(18933) <= 13891688;
srom_1(18934) <= 13445483;
srom_1(18935) <= 12975564;
srom_1(18936) <= 12484135;
srom_1(18937) <= 11973501;
srom_1(18938) <= 11446056;
srom_1(18939) <= 10904274;
srom_1(18940) <= 10350695;
srom_1(18941) <= 9787915;
srom_1(18942) <= 9218573;
srom_1(18943) <= 8645339;
srom_1(18944) <= 8070901;
srom_1(18945) <= 7497953;
srom_1(18946) <= 6929182;
srom_1(18947) <= 6367254;
srom_1(18948) <= 5814805;
srom_1(18949) <= 5274426;
srom_1(18950) <= 4748650;
srom_1(18951) <= 4239943;
srom_1(18952) <= 3750691;
srom_1(18953) <= 3283187;
srom_1(18954) <= 2839625;
srom_1(18955) <= 2422083;
srom_1(18956) <= 2032521;
srom_1(18957) <= 1672764;
srom_1(18958) <= 1344501;
srom_1(18959) <= 1049269;
srom_1(18960) <= 788454;
srom_1(18961) <= 563279;
srom_1(18962) <= 374800;
srom_1(18963) <= 223900;
srom_1(18964) <= 111287;
srom_1(18965) <= 37490;
srom_1(18966) <= 2854;
srom_1(18967) <= 7541;
srom_1(18968) <= 51530;
srom_1(18969) <= 134614;
srom_1(18970) <= 256405;
srom_1(18971) <= 416330;
srom_1(18972) <= 613639;
srom_1(18973) <= 847409;
srom_1(18974) <= 1116541;
srom_1(18975) <= 1419775;
srom_1(18976) <= 1755688;
srom_1(18977) <= 2122705;
srom_1(18978) <= 2519105;
srom_1(18979) <= 2943029;
srom_1(18980) <= 3392489;
srom_1(18981) <= 3865378;
srom_1(18982) <= 4359477;
srom_1(18983) <= 4872471;
srom_1(18984) <= 5401953;
srom_1(18985) <= 5945441;
srom_1(18986) <= 6500385;
srom_1(18987) <= 7064184;
srom_1(18988) <= 7634193;
srom_1(18989) <= 8207741;
srom_1(18990) <= 8782136;
srom_1(18991) <= 9354686;
srom_1(18992) <= 9922706;
srom_1(18993) <= 10483531;
srom_1(18994) <= 11034533;
srom_1(18995) <= 11573128;
srom_1(18996) <= 12096789;
srom_1(18997) <= 12603061;
srom_1(18998) <= 13089570;
srom_1(18999) <= 13554034;
srom_1(19000) <= 13994277;
srom_1(19001) <= 14408232;
srom_1(19002) <= 14793959;
srom_1(19003) <= 15149649;
srom_1(19004) <= 15473635;
srom_1(19005) <= 15764396;
srom_1(19006) <= 16020569;
srom_1(19007) <= 16240954;
srom_1(19008) <= 16424517;
srom_1(19009) <= 16570396;
srom_1(19010) <= 16677908;
srom_1(19011) <= 16746548;
srom_1(19012) <= 16775996;
srom_1(19013) <= 16766112;
srom_1(19014) <= 16716943;
srom_1(19015) <= 16628719;
srom_1(19016) <= 16501855;
srom_1(19017) <= 16336945;
srom_1(19018) <= 16134763;
srom_1(19019) <= 15896256;
srom_1(19020) <= 15622543;
srom_1(19021) <= 15314908;
srom_1(19022) <= 14974793;
srom_1(19023) <= 14603793;
srom_1(19024) <= 14203648;
srom_1(19025) <= 13776235;
srom_1(19026) <= 13323556;
srom_1(19027) <= 12847737;
srom_1(19028) <= 12351006;
srom_1(19029) <= 11835695;
srom_1(19030) <= 11304219;
srom_1(19031) <= 10759071;
srom_1(19032) <= 10202807;
srom_1(19033) <= 9638035;
srom_1(19034) <= 9067405;
srom_1(19035) <= 8493591;
srom_1(19036) <= 7919285;
srom_1(19037) <= 7347180;
srom_1(19038) <= 6779958;
srom_1(19039) <= 6220280;
srom_1(19040) <= 5670770;
srom_1(19041) <= 5134005;
srom_1(19042) <= 4612502;
srom_1(19043) <= 4108706;
srom_1(19044) <= 3624980;
srom_1(19045) <= 3163593;
srom_1(19046) <= 2726707;
srom_1(19047) <= 2316372;
srom_1(19048) <= 1934512;
srom_1(19049) <= 1582917;
srom_1(19050) <= 1263236;
srom_1(19051) <= 976969;
srom_1(19052) <= 725458;
srom_1(19053) <= 509881;
srom_1(19054) <= 331251;
srom_1(19055) <= 190404;
srom_1(19056) <= 88002;
srom_1(19057) <= 24523;
srom_1(19058) <= 267;
srom_1(19059) <= 15347;
srom_1(19060) <= 69692;
srom_1(19061) <= 163047;
srom_1(19062) <= 294975;
srom_1(19063) <= 464856;
srom_1(19064) <= 671895;
srom_1(19065) <= 915120;
srom_1(19066) <= 1193390;
srom_1(19067) <= 1505402;
srom_1(19068) <= 1849691;
srom_1(19069) <= 2224643;
srom_1(19070) <= 2628501;
srom_1(19071) <= 3059369;
srom_1(19072) <= 3515228;
srom_1(19073) <= 3993940;
srom_1(19074) <= 4493260;
srom_1(19075) <= 5010847;
srom_1(19076) <= 5544273;
srom_1(19077) <= 6091038;
srom_1(19078) <= 6648576;
srom_1(19079) <= 7214274;
srom_1(19080) <= 7785479;
srom_1(19081) <= 8359512;
srom_1(19082) <= 8933682;
srom_1(19083) <= 9505295;
srom_1(19084) <= 10071672;
srom_1(19085) <= 10630157;
srom_1(19086) <= 11178130;
srom_1(19087) <= 11713022;
srom_1(19088) <= 12232324;
srom_1(19089) <= 12733603;
srom_1(19090) <= 13214506;
srom_1(19091) <= 13672778;
srom_1(19092) <= 14106272;
srom_1(19093) <= 14512953;
srom_1(19094) <= 14890915;
srom_1(19095) <= 15238386;
srom_1(19096) <= 15553736;
srom_1(19097) <= 15835485;
srom_1(19098) <= 16082314;
srom_1(19099) <= 16293065;
srom_1(19100) <= 16466749;
srom_1(19101) <= 16602551;
srom_1(19102) <= 16699836;
srom_1(19103) <= 16758146;
srom_1(19104) <= 16777209;
srom_1(19105) <= 16756935;
srom_1(19106) <= 16697418;
srom_1(19107) <= 16598939;
srom_1(19108) <= 16461959;
srom_1(19109) <= 16287120;
srom_1(19110) <= 16075242;
srom_1(19111) <= 15827319;
srom_1(19112) <= 15544513;
srom_1(19113) <= 15228151;
srom_1(19114) <= 14879716;
srom_1(19115) <= 14500841;
srom_1(19116) <= 14093305;
srom_1(19117) <= 13659017;
srom_1(19118) <= 13200014;
srom_1(19119) <= 12718449;
srom_1(19120) <= 12216580;
srom_1(19121) <= 11696760;
srom_1(19122) <= 11161427;
srom_1(19123) <= 10613092;
srom_1(19124) <= 10054325;
srom_1(19125) <= 9487746;
srom_1(19126) <= 8916014;
srom_1(19127) <= 8341809;
srom_1(19128) <= 7767822;
srom_1(19129) <= 7196747;
srom_1(19130) <= 6631261;
srom_1(19131) <= 6074016;
srom_1(19132) <= 5527625;
srom_1(19133) <= 4994650;
srom_1(19134) <= 4477590;
srom_1(19135) <= 3978870;
srom_1(19136) <= 3500829;
srom_1(19137) <= 3045709;
srom_1(19138) <= 2615643;
srom_1(19139) <= 2212649;
srom_1(19140) <= 1838616;
srom_1(19141) <= 1495298;
srom_1(19142) <= 1184305;
srom_1(19143) <= 907096;
srom_1(19144) <= 664969;
srom_1(19145) <= 459062;
srom_1(19146) <= 290339;
srom_1(19147) <= 159592;
srom_1(19148) <= 67433;
srom_1(19149) <= 14295;
srom_1(19150) <= 428;
srom_1(19151) <= 25895;
srom_1(19152) <= 90578;
srom_1(19153) <= 194173;
srom_1(19154) <= 336194;
srom_1(19155) <= 515977;
srom_1(19156) <= 732676;
srom_1(19157) <= 985277;
srom_1(19158) <= 1272595;
srom_1(19159) <= 1593282;
srom_1(19160) <= 1945835;
srom_1(19161) <= 2328600;
srom_1(19162) <= 2739783;
srom_1(19163) <= 3177454;
srom_1(19164) <= 3639563;
srom_1(19165) <= 4123942;
srom_1(19166) <= 4628319;
srom_1(19167) <= 5150329;
srom_1(19168) <= 5687525;
srom_1(19169) <= 6237387;
srom_1(19170) <= 6797337;
srom_1(19171) <= 7364749;
srom_1(19172) <= 7936962;
srom_1(19173) <= 8511293;
srom_1(19174) <= 9085049;
srom_1(19175) <= 9655539;
srom_1(19176) <= 10220087;
srom_1(19177) <= 10776048;
srom_1(19178) <= 11320812;
srom_1(19179) <= 11851827;
srom_1(19180) <= 12366602;
srom_1(19181) <= 12862722;
srom_1(19182) <= 13337861;
srom_1(19183) <= 13789792;
srom_1(19184) <= 14216395;
srom_1(19185) <= 14615669;
srom_1(19186) <= 14985743;
srom_1(19187) <= 15324880;
srom_1(19188) <= 15631491;
srom_1(19189) <= 15904137;
srom_1(19190) <= 16141541;
srom_1(19191) <= 16342588;
srom_1(19192) <= 16506336;
srom_1(19193) <= 16632017;
srom_1(19194) <= 16719043;
srom_1(19195) <= 16767004;
srom_1(19196) <= 16775675;
srom_1(19197) <= 16745017;
srom_1(19198) <= 16675173;
srom_1(19199) <= 16566471;
srom_1(19200) <= 16419419;
srom_1(19201) <= 16234708;
srom_1(19202) <= 16013205;
srom_1(19203) <= 15755946;
srom_1(19204) <= 15464140;
srom_1(19205) <= 15139154;
srom_1(19206) <= 14782513;
srom_1(19207) <= 14395888;
srom_1(19208) <= 13981094;
srom_1(19209) <= 13540074;
srom_1(19210) <= 13074897;
srom_1(19211) <= 12587744;
srom_1(19212) <= 12080900;
srom_1(19213) <= 11556742;
srom_1(19214) <= 11017728;
srom_1(19215) <= 10466384;
srom_1(19216) <= 9905297;
srom_1(19217) <= 9337098;
srom_1(19218) <= 8764451;
srom_1(19219) <= 8190041;
srom_1(19220) <= 7616563;
srom_1(19221) <= 7046705;
srom_1(19222) <= 6483140;
srom_1(19223) <= 5928510;
srom_1(19224) <= 5385416;
srom_1(19225) <= 4856405;
srom_1(19226) <= 4343958;
srom_1(19227) <= 3850478;
srom_1(19228) <= 3378279;
srom_1(19229) <= 2929574;
srom_1(19230) <= 2506469;
srom_1(19231) <= 2110948;
srom_1(19232) <= 1744864;
srom_1(19233) <= 1409936;
srom_1(19234) <= 1107732;
srom_1(19235) <= 839671;
srom_1(19236) <= 607010;
srom_1(19237) <= 410839;
srom_1(19238) <= 252079;
srom_1(19239) <= 131474;
srom_1(19240) <= 49589;
srom_1(19241) <= 6809;
srom_1(19242) <= 3334;
srom_1(19243) <= 39180;
srom_1(19244) <= 114180;
srom_1(19245) <= 227981;
srom_1(19246) <= 380051;
srom_1(19247) <= 569675;
srom_1(19248) <= 795965;
srom_1(19249) <= 1057859;
srom_1(19250) <= 1354130;
srom_1(19251) <= 1683387;
srom_1(19252) <= 2044088;
srom_1(19253) <= 2434541;
srom_1(19254) <= 2852914;
srom_1(19255) <= 3297246;
srom_1(19256) <= 3765453;
srom_1(19257) <= 4255340;
srom_1(19258) <= 4764608;
srom_1(19259) <= 5290872;
srom_1(19260) <= 5831661;
srom_1(19261) <= 6384441;
srom_1(19262) <= 6946619;
srom_1(19263) <= 7515559;
srom_1(19264) <= 8088593;
srom_1(19265) <= 8663034;
srom_1(19266) <= 9236188;
srom_1(19267) <= 9805367;
srom_1(19268) <= 10367903;
srom_1(19269) <= 10921157;
srom_1(19270) <= 11462535;
srom_1(19271) <= 11989499;
srom_1(19272) <= 12499576;
srom_1(19273) <= 12990376;
srom_1(19274) <= 13459597;
srom_1(19275) <= 13905038;
srom_1(19276) <= 14324610;
srom_1(19277) <= 14716347;
srom_1(19278) <= 15078411;
srom_1(19279) <= 15409103;
srom_1(19280) <= 15706875;
srom_1(19281) <= 15970328;
srom_1(19282) <= 16198228;
srom_1(19283) <= 16389507;
srom_1(19284) <= 16543266;
srom_1(19285) <= 16658785;
srom_1(19286) <= 16735522;
srom_1(19287) <= 16773118;
srom_1(19288) <= 16771396;
srom_1(19289) <= 16730365;
srom_1(19290) <= 16650215;
srom_1(19291) <= 16531325;
srom_1(19292) <= 16374250;
srom_1(19293) <= 16179728;
srom_1(19294) <= 15948671;
srom_1(19295) <= 15682162;
srom_1(19296) <= 15381451;
srom_1(19297) <= 15047948;
srom_1(19298) <= 14683217;
srom_1(19299) <= 14288969;
srom_1(19300) <= 13867051;
srom_1(19301) <= 13419444;
srom_1(19302) <= 12948245;
srom_1(19303) <= 12455664;
srom_1(19304) <= 11944012;
srom_1(19305) <= 11415687;
srom_1(19306) <= 10873167;
srom_1(19307) <= 10318996;
srom_1(19308) <= 9755773;
srom_1(19309) <= 9186139;
srom_1(19310) <= 8612765;
srom_1(19311) <= 8038339;
srom_1(19312) <= 7465556;
srom_1(19313) <= 6897102;
srom_1(19314) <= 6335642;
srom_1(19315) <= 5783809;
srom_1(19316) <= 5244191;
srom_1(19317) <= 4719318;
srom_1(19318) <= 4211651;
srom_1(19319) <= 3723572;
srom_1(19320) <= 3257368;
srom_1(19321) <= 2815227;
srom_1(19322) <= 2399221;
srom_1(19323) <= 2011302;
srom_1(19324) <= 1653288;
srom_1(19325) <= 1326858;
srom_1(19326) <= 1033543;
srom_1(19327) <= 774719;
srom_1(19328) <= 551598;
srom_1(19329) <= 365228;
srom_1(19330) <= 216483;
srom_1(19331) <= 106059;
srom_1(19332) <= 34475;
srom_1(19333) <= 2067;
srom_1(19334) <= 8986;
srom_1(19335) <= 55199;
srom_1(19336) <= 140491;
srom_1(19337) <= 264462;
srom_1(19338) <= 426529;
srom_1(19339) <= 625933;
srom_1(19340) <= 861739;
srom_1(19341) <= 1132840;
srom_1(19342) <= 1437967;
srom_1(19343) <= 1775688;
srom_1(19344) <= 2144419;
srom_1(19345) <= 2542431;
srom_1(19346) <= 2967858;
srom_1(19347) <= 3418704;
srom_1(19348) <= 3892856;
srom_1(19349) <= 4388090;
srom_1(19350) <= 4902084;
srom_1(19351) <= 5432428;
srom_1(19352) <= 5976634;
srom_1(19353) <= 6532151;
srom_1(19354) <= 7096373;
srom_1(19355) <= 7666655;
srom_1(19356) <= 8240322;
srom_1(19357) <= 8814685;
srom_1(19358) <= 9387050;
srom_1(19359) <= 9954732;
srom_1(19360) <= 10515071;
srom_1(19361) <= 11065438;
srom_1(19362) <= 11603252;
srom_1(19363) <= 12125992;
srom_1(19364) <= 12631205;
srom_1(19365) <= 13116524;
srom_1(19366) <= 13579672;
srom_1(19367) <= 14018478;
srom_1(19368) <= 14430882;
srom_1(19369) <= 14814953;
srom_1(19370) <= 15168888;
srom_1(19371) <= 15491028;
srom_1(19372) <= 15779863;
srom_1(19373) <= 16034037;
srom_1(19374) <= 16252359;
srom_1(19375) <= 16433806;
srom_1(19376) <= 16577526;
srom_1(19377) <= 16682845;
srom_1(19378) <= 16749269;
srom_1(19379) <= 16776488;
srom_1(19380) <= 16764373;
srom_1(19381) <= 16712981;
srom_1(19382) <= 16622553;
srom_1(19383) <= 16493513;
srom_1(19384) <= 16326467;
srom_1(19385) <= 16122197;
srom_1(19386) <= 15881662;
srom_1(19387) <= 15605989;
srom_1(19388) <= 15296472;
srom_1(19389) <= 14954561;
srom_1(19390) <= 14581860;
srom_1(19391) <= 14180117;
srom_1(19392) <= 13751216;
srom_1(19393) <= 13297167;
srom_1(19394) <= 12820101;
srom_1(19395) <= 12322253;
srom_1(19396) <= 11805960;
srom_1(19397) <= 11273641;
srom_1(19398) <= 10727793;
srom_1(19399) <= 10170976;
srom_1(19400) <= 9605801;
srom_1(19401) <= 9034919;
srom_1(19402) <= 8461005;
srom_1(19403) <= 7886752;
srom_1(19404) <= 7314852;
srom_1(19405) <= 6747988;
srom_1(19406) <= 6188816;
srom_1(19407) <= 5639961;
srom_1(19408) <= 5103995;
srom_1(19409) <= 4583431;
srom_1(19410) <= 4080711;
srom_1(19411) <= 3598193;
srom_1(19412) <= 3138138;
srom_1(19413) <= 2702705;
srom_1(19414) <= 2293934;
srom_1(19415) <= 1913744;
srom_1(19416) <= 1563917;
srom_1(19417) <= 1246093;
srom_1(19418) <= 961762;
srom_1(19419) <= 712259;
srom_1(19420) <= 498752;
srom_1(19421) <= 322244;
srom_1(19422) <= 183562;
srom_1(19423) <= 83356;
srom_1(19424) <= 22097;
srom_1(19425) <= 70;
srom_1(19426) <= 17381;
srom_1(19427) <= 73947;
srom_1(19428) <= 169503;
srom_1(19429) <= 303602;
srom_1(19430) <= 475613;
srom_1(19431) <= 684732;
srom_1(19432) <= 929977;
srom_1(19433) <= 1210198;
srom_1(19434) <= 1524080;
srom_1(19435) <= 1870153;
srom_1(19436) <= 2246794;
srom_1(19437) <= 2652235;
srom_1(19438) <= 3084576;
srom_1(19439) <= 3541789;
srom_1(19440) <= 4021731;
srom_1(19441) <= 4522151;
srom_1(19442) <= 5040702;
srom_1(19443) <= 5574952;
srom_1(19444) <= 6122397;
srom_1(19445) <= 6680468;
srom_1(19446) <= 7246550;
srom_1(19447) <= 7817987;
srom_1(19448) <= 8392100;
srom_1(19449) <= 8966196;
srom_1(19450) <= 9537584;
srom_1(19451) <= 10103584;
srom_1(19452) <= 10661542;
srom_1(19453) <= 11208842;
srom_1(19454) <= 11742916;
srom_1(19455) <= 12261261;
srom_1(19456) <= 12761445;
srom_1(19457) <= 13241124;
srom_1(19458) <= 13698048;
srom_1(19459) <= 14130074;
srom_1(19460) <= 14535176;
srom_1(19461) <= 14911455;
srom_1(19462) <= 15257146;
srom_1(19463) <= 15570628;
srom_1(19464) <= 15850431;
srom_1(19465) <= 16095243;
srom_1(19466) <= 16303916;
srom_1(19467) <= 16475471;
srom_1(19468) <= 16609105;
srom_1(19469) <= 16704189;
srom_1(19470) <= 16760279;
srom_1(19471) <= 16777111;
srom_1(19472) <= 16754607;
srom_1(19473) <= 16692871;
srom_1(19474) <= 16592194;
srom_1(19475) <= 16453048;
srom_1(19476) <= 16276085;
srom_1(19477) <= 16062134;
srom_1(19478) <= 15812200;
srom_1(19479) <= 15527454;
srom_1(19480) <= 15209231;
srom_1(19481) <= 14859025;
srom_1(19482) <= 14478476;
srom_1(19483) <= 14069370;
srom_1(19484) <= 13633624;
srom_1(19485) <= 13173283;
srom_1(19486) <= 12690505;
srom_1(19487) <= 12187554;
srom_1(19488) <= 11666788;
srom_1(19489) <= 11130650;
srom_1(19490) <= 10581654;
srom_1(19491) <= 10022373;
srom_1(19492) <= 9455431;
srom_1(19493) <= 8883487;
srom_1(19494) <= 8309222;
srom_1(19495) <= 7735329;
srom_1(19496) <= 7164499;
srom_1(19497) <= 6599410;
srom_1(19498) <= 6042711;
srom_1(19499) <= 5497013;
srom_1(19500) <= 4964874;
srom_1(19501) <= 4448790;
srom_1(19502) <= 3951182;
srom_1(19503) <= 3474382;
srom_1(19504) <= 3020627;
srom_1(19505) <= 2592043;
srom_1(19506) <= 2190642;
srom_1(19507) <= 1818306;
srom_1(19508) <= 1476780;
srom_1(19509) <= 1167665;
srom_1(19510) <= 892413;
srom_1(19511) <= 652312;
srom_1(19512) <= 448490;
srom_1(19513) <= 281901;
srom_1(19514) <= 153328;
srom_1(19515) <= 63372;
srom_1(19516) <= 12457;
srom_1(19517) <= 820;
srom_1(19518) <= 28516;
srom_1(19519) <= 95416;
srom_1(19520) <= 201206;
srom_1(19521) <= 345388;
srom_1(19522) <= 527289;
srom_1(19523) <= 746054;
srom_1(19524) <= 1000657;
srom_1(19525) <= 1289905;
srom_1(19526) <= 1612441;
srom_1(19527) <= 1966753;
srom_1(19528) <= 2351179;
srom_1(19529) <= 2763917;
srom_1(19530) <= 3203031;
srom_1(19531) <= 3666462;
srom_1(19532) <= 4152036;
srom_1(19533) <= 4657478;
srom_1(19534) <= 5180415;
srom_1(19535) <= 5718398;
srom_1(19536) <= 6268901;
srom_1(19537) <= 6829345;
srom_1(19538) <= 7397101;
srom_1(19539) <= 7969506;
srom_1(19540) <= 8543876;
srom_1(19541) <= 9117519;
srom_1(19542) <= 9687743;
srom_1(19543) <= 10251875;
srom_1(19544) <= 10807270;
srom_1(19545) <= 11351322;
srom_1(19546) <= 11881482;
srom_1(19547) <= 12395262;
srom_1(19548) <= 12890254;
srom_1(19549) <= 13364136;
srom_1(19550) <= 13814686;
srom_1(19551) <= 14239791;
srom_1(19552) <= 14637458;
srom_1(19553) <= 15005821;
srom_1(19554) <= 15343155;
srom_1(19555) <= 15647876;
srom_1(19556) <= 15918556;
srom_1(19557) <= 16153926;
srom_1(19558) <= 16352881;
srom_1(19559) <= 16514489;
srom_1(19560) <= 16637992;
srom_1(19561) <= 16722811;
srom_1(19562) <= 16768548;
srom_1(19563) <= 16774988;
srom_1(19564) <= 16742102;
srom_1(19565) <= 16670043;
srom_1(19566) <= 16559150;
srom_1(19567) <= 16409943;
srom_1(19568) <= 16223120;
srom_1(19569) <= 15999559;
srom_1(19570) <= 15740308;
srom_1(19571) <= 15446581;
srom_1(19572) <= 15119758;
srom_1(19573) <= 14761370;
srom_1(19574) <= 14373098;
srom_1(19575) <= 13956762;
srom_1(19576) <= 13514316;
srom_1(19577) <= 13047833;
srom_1(19578) <= 12559502;
srom_1(19579) <= 12051611;
srom_1(19580) <= 11526544;
srom_1(19581) <= 10986762;
srom_1(19582) <= 10434796;
srom_1(19583) <= 9873235;
srom_1(19584) <= 9304712;
srom_1(19585) <= 8731893;
srom_1(19586) <= 8157464;
srom_1(19587) <= 7584119;
srom_1(19588) <= 7014547;
srom_1(19589) <= 6451418;
srom_1(19590) <= 5897374;
srom_1(19591) <= 5355011;
srom_1(19592) <= 4826874;
srom_1(19593) <= 4315439;
srom_1(19594) <= 3823105;
srom_1(19595) <= 3352180;
srom_1(19596) <= 2904873;
srom_1(19597) <= 2483280;
srom_1(19598) <= 2089380;
srom_1(19599) <= 1725019;
srom_1(19600) <= 1391906;
srom_1(19601) <= 1091602;
srom_1(19602) <= 825517;
srom_1(19603) <= 594898;
srom_1(19604) <= 400826;
srom_1(19605) <= 244212;
srom_1(19606) <= 125789;
srom_1(19607) <= 46114;
srom_1(19608) <= 5559;
srom_1(19609) <= 4316;
srom_1(19610) <= 42389;
srom_1(19611) <= 119601;
srom_1(19612) <= 235589;
srom_1(19613) <= 389809;
srom_1(19614) <= 581538;
srom_1(19615) <= 809877;
srom_1(19616) <= 1073756;
srom_1(19617) <= 1371936;
srom_1(19618) <= 1703020;
srom_1(19619) <= 2065455;
srom_1(19620) <= 2457541;
srom_1(19621) <= 2877440;
srom_1(19622) <= 3323183;
srom_1(19623) <= 3792680;
srom_1(19624) <= 4283728;
srom_1(19625) <= 4794026;
srom_1(19626) <= 5321179;
srom_1(19627) <= 5862717;
srom_1(19628) <= 6416100;
srom_1(19629) <= 6978732;
srom_1(19630) <= 7547976;
srom_1(19631) <= 8121162;
srom_1(19632) <= 8695602;
srom_1(19633) <= 9268602;
srom_1(19634) <= 9837476;
srom_1(19635) <= 10399556;
srom_1(19636) <= 10952205;
srom_1(19637) <= 11492833;
srom_1(19638) <= 12018904;
srom_1(19639) <= 12527952;
srom_1(19640) <= 13017588;
srom_1(19641) <= 13485518;
srom_1(19642) <= 13929547;
srom_1(19643) <= 14347592;
srom_1(19644) <= 14737693;
srom_1(19645) <= 15098022;
srom_1(19646) <= 15426887;
srom_1(19647) <= 15722748;
srom_1(19648) <= 15984216;
srom_1(19649) <= 16210066;
srom_1(19650) <= 16399239;
srom_1(19651) <= 16550847;
srom_1(19652) <= 16664179;
srom_1(19653) <= 16738704;
srom_1(19654) <= 16774073;
srom_1(19655) <= 16770120;
srom_1(19656) <= 16726862;
srom_1(19657) <= 16644504;
srom_1(19658) <= 16523431;
srom_1(19659) <= 16364211;
srom_1(19660) <= 16167591;
srom_1(19661) <= 15934492;
srom_1(19662) <= 15666008;
srom_1(19663) <= 15363398;
srom_1(19664) <= 15028081;
srom_1(19665) <= 14661629;
srom_1(19666) <= 14265760;
srom_1(19667) <= 13842332;
srom_1(19668) <= 13393329;
srom_1(19669) <= 12920857;
srom_1(19670) <= 12427132;
srom_1(19671) <= 11914469;
srom_1(19672) <= 11385272;
srom_1(19673) <= 10842023;
srom_1(19674) <= 10287269;
srom_1(19675) <= 9723611;
srom_1(19676) <= 9153693;
srom_1(19677) <= 8580187;
srom_1(19678) <= 8005783;
srom_1(19679) <= 7433174;
srom_1(19680) <= 6865045;
srom_1(19681) <= 6304061;
srom_1(19682) <= 5752852;
srom_1(19683) <= 5214003;
srom_1(19684) <= 4690040;
srom_1(19685) <= 4183422;
srom_1(19686) <= 3696523;
srom_1(19687) <= 3231627;
srom_1(19688) <= 2790914;
srom_1(19689) <= 2376450;
srom_1(19690) <= 1990180;
srom_1(19691) <= 1633913;
srom_1(19692) <= 1309322;
srom_1(19693) <= 1017928;
srom_1(19694) <= 761098;
srom_1(19695) <= 540036;
srom_1(19696) <= 355778;
srom_1(19697) <= 209189;
srom_1(19698) <= 100956;
srom_1(19699) <= 31587;
srom_1(19700) <= 1407;
srom_1(19701) <= 10557;
srom_1(19702) <= 58995;
srom_1(19703) <= 146493;
srom_1(19704) <= 272641;
srom_1(19705) <= 436848;
srom_1(19706) <= 638343;
srom_1(19707) <= 876182;
srom_1(19708) <= 1149249;
srom_1(19709) <= 1456265;
srom_1(19710) <= 1795788;
srom_1(19711) <= 2166227;
srom_1(19712) <= 2565845;
srom_1(19713) <= 2992768;
srom_1(19714) <= 3444994;
srom_1(19715) <= 3920403;
srom_1(19716) <= 4416764;
srom_1(19717) <= 4931750;
srom_1(19718) <= 5462947;
srom_1(19719) <= 6007864;
srom_1(19720) <= 6563944;
srom_1(19721) <= 7128581;
srom_1(19722) <= 7699127;
srom_1(19723) <= 8272906;
srom_1(19724) <= 8847227;
srom_1(19725) <= 9419398;
srom_1(19726) <= 9986735;
srom_1(19727) <= 10546578;
srom_1(19728) <= 11096302;
srom_1(19729) <= 11633328;
srom_1(19730) <= 12155138;
srom_1(19731) <= 12659286;
srom_1(19732) <= 13143407;
srom_1(19733) <= 13605232;
srom_1(19734) <= 14042594;
srom_1(19735) <= 14453442;
srom_1(19736) <= 14835850;
srom_1(19737) <= 15188025;
srom_1(19738) <= 15508315;
srom_1(19739) <= 15795218;
srom_1(19740) <= 16047390;
srom_1(19741) <= 16263646;
srom_1(19742) <= 16442974;
srom_1(19743) <= 16584532;
srom_1(19744) <= 16687656;
srom_1(19745) <= 16751864;
srom_1(19746) <= 16776853;
srom_1(19747) <= 16762507;
srom_1(19748) <= 16708893;
srom_1(19749) <= 16616262;
srom_1(19750) <= 16485049;
srom_1(19751) <= 16315869;
srom_1(19752) <= 16109515;
srom_1(19753) <= 15866955;
srom_1(19754) <= 15589326;
srom_1(19755) <= 15277931;
srom_1(19756) <= 14934230;
srom_1(19757) <= 14559834;
srom_1(19758) <= 14156499;
srom_1(19759) <= 13726116;
srom_1(19760) <= 13270704;
srom_1(19761) <= 12792398;
srom_1(19762) <= 12293441;
srom_1(19763) <= 11776173;
srom_1(19764) <= 11243019;
srom_1(19765) <= 10696481;
srom_1(19766) <= 10139119;
srom_1(19767) <= 9573549;
srom_1(19768) <= 9002423;
srom_1(19769) <= 8428418;
srom_1(19770) <= 7854226;
srom_1(19771) <= 7282541;
srom_1(19772) <= 6716041;
srom_1(19773) <= 6157386;
srom_1(19774) <= 5609193;
srom_1(19775) <= 5074034;
srom_1(19776) <= 4554418;
srom_1(19777) <= 4052781;
srom_1(19778) <= 3571477;
srom_1(19779) <= 3112762;
srom_1(19780) <= 2678788;
srom_1(19781) <= 2271588;
srom_1(19782) <= 1893074;
srom_1(19783) <= 1545019;
srom_1(19784) <= 1229056;
srom_1(19785) <= 946667;
srom_1(19786) <= 699176;
srom_1(19787) <= 487743;
srom_1(19788) <= 313360;
srom_1(19789) <= 176844;
srom_1(19790) <= 78836;
srom_1(19791) <= 19796;
srom_1(19792) <= 0;
srom_1(19793) <= 19541;
srom_1(19794) <= 78327;
srom_1(19795) <= 176083;
srom_1(19796) <= 312350;
srom_1(19797) <= 486490;
srom_1(19798) <= 697686;
srom_1(19799) <= 944946;
srom_1(19800) <= 1227113;
srom_1(19801) <= 1542863;
srom_1(19802) <= 1890714;
srom_1(19803) <= 2269036;
srom_1(19804) <= 2676056;
srom_1(19805) <= 3109863;
srom_1(19806) <= 3568424;
srom_1(19807) <= 4049588;
srom_1(19808) <= 4551100;
srom_1(19809) <= 5070607;
srom_1(19810) <= 5605673;
srom_1(19811) <= 6153790;
srom_1(19812) <= 6712386;
srom_1(19813) <= 7278843;
srom_1(19814) <= 7850503;
srom_1(19815) <= 8424688;
srom_1(19816) <= 8998702;
srom_1(19817) <= 9569856;
srom_1(19818) <= 10135471;
srom_1(19819) <= 10692894;
srom_1(19820) <= 11239511;
srom_1(19821) <= 11772760;
srom_1(19822) <= 12290139;
srom_1(19823) <= 12789222;
srom_1(19824) <= 13267670;
srom_1(19825) <= 13723238;
srom_1(19826) <= 14153789;
srom_1(19827) <= 14557306;
srom_1(19828) <= 14931896;
srom_1(19829) <= 15275802;
srom_1(19830) <= 15587412;
srom_1(19831) <= 15865264;
srom_1(19832) <= 16108055;
srom_1(19833) <= 16314648;
srom_1(19834) <= 16484072;
srom_1(19835) <= 16615534;
srom_1(19836) <= 16708417;
srom_1(19837) <= 16762285;
srom_1(19838) <= 16776887;
srom_1(19839) <= 16752153;
srom_1(19840) <= 16688199;
srom_1(19841) <= 16585326;
srom_1(19842) <= 16444016;
srom_1(19843) <= 16264931;
srom_1(19844) <= 16048911;
srom_1(19845) <= 15796969;
srom_1(19846) <= 15510287;
srom_1(19847) <= 15190209;
srom_1(19848) <= 14838236;
srom_1(19849) <= 14456018;
srom_1(19850) <= 14045349;
srom_1(19851) <= 13608153;
srom_1(19852) <= 13146480;
srom_1(19853) <= 12662496;
srom_1(19854) <= 12158471;
srom_1(19855) <= 11636767;
srom_1(19856) <= 11099832;
srom_1(19857) <= 10550183;
srom_1(19858) <= 9990397;
srom_1(19859) <= 9423100;
srom_1(19860) <= 8850952;
srom_1(19861) <= 8276636;
srom_1(19862) <= 7702845;
srom_1(19863) <= 7132270;
srom_1(19864) <= 6567586;
srom_1(19865) <= 6011441;
srom_1(19866) <= 5466444;
srom_1(19867) <= 4935150;
srom_1(19868) <= 4420050;
srom_1(19869) <= 3923560;
srom_1(19870) <= 3448009;
srom_1(19871) <= 2995625;
srom_1(19872) <= 2568531;
srom_1(19873) <= 2168730;
srom_1(19874) <= 1798095;
srom_1(19875) <= 1458366;
srom_1(19876) <= 1151135;
srom_1(19877) <= 877843;
srom_1(19878) <= 639771;
srom_1(19879) <= 438037;
srom_1(19880) <= 273585;
srom_1(19881) <= 147188;
srom_1(19882) <= 59437;
srom_1(19883) <= 10745;
srom_1(19884) <= 1339;
srom_1(19885) <= 31264;
srom_1(19886) <= 100380;
srom_1(19887) <= 208362;
srom_1(19888) <= 354704;
srom_1(19889) <= 538720;
srom_1(19890) <= 759546;
srom_1(19891) <= 1016148;
srom_1(19892) <= 1307322;
srom_1(19893) <= 1631702;
srom_1(19894) <= 1987768;
srom_1(19895) <= 2373849;
srom_1(19896) <= 2788136;
srom_1(19897) <= 3228685;
srom_1(19898) <= 3693431;
srom_1(19899) <= 4180195;
srom_1(19900) <= 4686693;
srom_1(19901) <= 5210550;
srom_1(19902) <= 5749310;
srom_1(19903) <= 6300448;
srom_1(19904) <= 6861377;
srom_1(19905) <= 7429468;
srom_1(19906) <= 8002056;
srom_1(19907) <= 8576457;
srom_1(19908) <= 9149978;
srom_1(19909) <= 9719928;
srom_1(19910) <= 10283635;
srom_1(19911) <= 10838455;
srom_1(19912) <= 11381788;
srom_1(19913) <= 11911084;
srom_1(19914) <= 12423862;
srom_1(19915) <= 12917718;
srom_1(19916) <= 13390335;
srom_1(19917) <= 13839497;
srom_1(19918) <= 14263098;
srom_1(19919) <= 14659151;
srom_1(19920) <= 15025800;
srom_1(19921) <= 15361325;
srom_1(19922) <= 15664152;
srom_1(19923) <= 15932862;
srom_1(19924) <= 16166194;
srom_1(19925) <= 16363054;
srom_1(19926) <= 16522520;
srom_1(19927) <= 16643842;
srom_1(19928) <= 16726453;
srom_1(19929) <= 16769965;
srom_1(19930) <= 16774174;
srom_1(19931) <= 16739060;
srom_1(19932) <= 16664788;
srom_1(19933) <= 16551707;
srom_1(19934) <= 16400345;
srom_1(19935) <= 16211414;
srom_1(19936) <= 15985799;
srom_1(19937) <= 15724558;
srom_1(19938) <= 15428916;
srom_1(19939) <= 15100260;
srom_1(19940) <= 14740131;
srom_1(19941) <= 14350217;
srom_1(19942) <= 13932347;
srom_1(19943) <= 13488480;
srom_1(19944) <= 13020699;
srom_1(19945) <= 12531196;
srom_1(19946) <= 12022267;
srom_1(19947) <= 11496298;
srom_1(19948) <= 10955757;
srom_1(19949) <= 10403177;
srom_1(19950) <= 9841150;
srom_1(19951) <= 9272312;
srom_1(19952) <= 8699330;
srom_1(19953) <= 8124891;
srom_1(19954) <= 7551688;
srom_1(19955) <= 6982410;
srom_1(19956) <= 6419726;
srom_1(19957) <= 5866275;
srom_1(19958) <= 5324652;
srom_1(19959) <= 4797397;
srom_1(19960) <= 4286982;
srom_1(19961) <= 3795801;
srom_1(19962) <= 3326157;
srom_1(19963) <= 2880253;
srom_1(19964) <= 2460180;
srom_1(19965) <= 2067907;
srom_1(19966) <= 1705274;
srom_1(19967) <= 1373981;
srom_1(19968) <= 1075582;
srom_1(19969) <= 811477;
srom_1(19970) <= 582903;
srom_1(19971) <= 390933;
srom_1(19972) <= 236467;
srom_1(19973) <= 120229;
srom_1(19974) <= 42765;
srom_1(19975) <= 4436;
srom_1(19976) <= 5425;
srom_1(19977) <= 45724;
srom_1(19978) <= 125147;
srom_1(19979) <= 243319;
srom_1(19980) <= 399688;
srom_1(19981) <= 593519;
srom_1(19982) <= 823904;
srom_1(19983) <= 1089763;
srom_1(19984) <= 1389848;
srom_1(19985) <= 1722753;
srom_1(19986) <= 2086917;
srom_1(19987) <= 2480631;
srom_1(19988) <= 2902050;
srom_1(19989) <= 3349197;
srom_1(19990) <= 3819976;
srom_1(19991) <= 4312179;
srom_1(19992) <= 4823497;
srom_1(19993) <= 5351533;
srom_1(19994) <= 5893812;
srom_1(19995) <= 6447789;
srom_1(19996) <= 7010867;
srom_1(19997) <= 7580406;
srom_1(19998) <= 8153735;
srom_1(19999) <= 8728166;
srom_1(20000) <= 9301004;
srom_1(20001) <= 9869563;
srom_1(20002) <= 10431178;
srom_1(20003) <= 10983215;
srom_1(20004) <= 11523084;
srom_1(20005) <= 12048255;
srom_1(20006) <= 12556265;
srom_1(20007) <= 13044730;
srom_1(20008) <= 13511362;
srom_1(20009) <= 13953972;
srom_1(20010) <= 14370483;
srom_1(20011) <= 14758943;
srom_1(20012) <= 15117531;
srom_1(20013) <= 15444565;
srom_1(20014) <= 15738510;
srom_1(20015) <= 15997990;
srom_1(20016) <= 16221786;
srom_1(20017) <= 16408850;
srom_1(20018) <= 16558304;
srom_1(20019) <= 16669448;
srom_1(20020) <= 16741760;
srom_1(20021) <= 16774901;
srom_1(20022) <= 16768716;
srom_1(20023) <= 16723234;
srom_1(20024) <= 16638668;
srom_1(20025) <= 16515415;
srom_1(20026) <= 16354052;
srom_1(20027) <= 16155336;
srom_1(20028) <= 15920200;
srom_1(20029) <= 15649745;
srom_1(20030) <= 15345240;
srom_1(20031) <= 15008114;
srom_1(20032) <= 14639946;
srom_1(20033) <= 14242463;
srom_1(20034) <= 13817530;
srom_1(20035) <= 13367139;
srom_1(20036) <= 12893401;
srom_1(20037) <= 12398539;
srom_1(20038) <= 11884873;
srom_1(20039) <= 11354812;
srom_1(20040) <= 10810842;
srom_1(20041) <= 10255512;
srom_1(20042) <= 9691428;
srom_1(20043) <= 9121235;
srom_1(20044) <= 8547606;
srom_1(20045) <= 7973232;
srom_1(20046) <= 7400805;
srom_1(20047) <= 6833011;
srom_1(20048) <= 6272511;
srom_1(20049) <= 5721934;
srom_1(20050) <= 5183863;
srom_1(20051) <= 4660819;
srom_1(20052) <= 4155256;
srom_1(20053) <= 3669545;
srom_1(20054) <= 3205964;
srom_1(20055) <= 2766685;
srom_1(20056) <= 2353770;
srom_1(20057) <= 1969154;
srom_1(20058) <= 1614641;
srom_1(20059) <= 1291893;
srom_1(20060) <= 1002424;
srom_1(20061) <= 747592;
srom_1(20062) <= 528591;
srom_1(20063) <= 346449;
srom_1(20064) <= 202019;
srom_1(20065) <= 95978;
srom_1(20066) <= 28825;
srom_1(20067) <= 873;
srom_1(20068) <= 12254;
srom_1(20069) <= 62915;
srom_1(20070) <= 152618;
srom_1(20071) <= 280943;
srom_1(20072) <= 447287;
srom_1(20073) <= 650870;
srom_1(20074) <= 890739;
srom_1(20075) <= 1165768;
srom_1(20076) <= 1474666;
srom_1(20077) <= 1815987;
srom_1(20078) <= 2188129;
srom_1(20079) <= 2589348;
srom_1(20080) <= 3017760;
srom_1(20081) <= 3471359;
srom_1(20082) <= 3948016;
srom_1(20083) <= 4445497;
srom_1(20084) <= 4961469;
srom_1(20085) <= 5493511;
srom_1(20086) <= 6039130;
srom_1(20087) <= 6595766;
srom_1(20088) <= 7160809;
srom_1(20089) <= 7731610;
srom_1(20090) <= 8305491;
srom_1(20091) <= 8879763;
srom_1(20092) <= 9451731;
srom_1(20093) <= 10018714;
srom_1(20094) <= 10578053;
srom_1(20095) <= 11127125;
srom_1(20096) <= 11663354;
srom_1(20097) <= 12184228;
srom_1(20098) <= 12687302;
srom_1(20099) <= 13170219;
srom_1(20100) <= 13630712;
srom_1(20101) <= 14066624;
srom_1(20102) <= 14475910;
srom_1(20103) <= 14856650;
srom_1(20104) <= 15207059;
srom_1(20105) <= 15525494;
srom_1(20106) <= 15810462;
srom_1(20107) <= 16060626;
srom_1(20108) <= 16274814;
srom_1(20109) <= 16452020;
srom_1(20110) <= 16591414;
srom_1(20111) <= 16692343;
srom_1(20112) <= 16754332;
srom_1(20113) <= 16777092;
srom_1(20114) <= 16760515;
srom_1(20115) <= 16704679;
srom_1(20116) <= 16609847;
srom_1(20117) <= 16476462;
srom_1(20118) <= 16305151;
srom_1(20119) <= 16096716;
srom_1(20120) <= 15852135;
srom_1(20121) <= 15572555;
srom_1(20122) <= 15259287;
srom_1(20123) <= 14913800;
srom_1(20124) <= 14537714;
srom_1(20125) <= 14132793;
srom_1(20126) <= 13700936;
srom_1(20127) <= 13244167;
srom_1(20128) <= 12764628;
srom_1(20129) <= 12264570;
srom_1(20130) <= 11746335;
srom_1(20131) <= 11212355;
srom_1(20132) <= 10665133;
srom_1(20133) <= 10107236;
srom_1(20134) <= 9541280;
srom_1(20135) <= 8969918;
srom_1(20136) <= 8395830;
srom_1(20137) <= 7821709;
srom_1(20138) <= 7250246;
srom_1(20139) <= 6684121;
srom_1(20140) <= 6125989;
srom_1(20141) <= 5578467;
srom_1(20142) <= 5044123;
srom_1(20143) <= 4525462;
srom_1(20144) <= 4024917;
srom_1(20145) <= 3544835;
srom_1(20146) <= 3087467;
srom_1(20147) <= 2654957;
srom_1(20148) <= 2249335;
srom_1(20149) <= 1872502;
srom_1(20150) <= 1526225;
srom_1(20151) <= 1212128;
srom_1(20152) <= 931685;
srom_1(20153) <= 686209;
srom_1(20154) <= 476852;
srom_1(20155) <= 304597;
srom_1(20156) <= 170250;
srom_1(20157) <= 74442;
srom_1(20158) <= 17622;
srom_1(20159) <= 56;
srom_1(20160) <= 21827;
srom_1(20161) <= 82832;
srom_1(20162) <= 182787;
srom_1(20163) <= 321221;
srom_1(20164) <= 497486;
srom_1(20165) <= 710755;
srom_1(20166) <= 960028;
srom_1(20167) <= 1244137;
srom_1(20168) <= 1561748;
srom_1(20169) <= 1911373;
srom_1(20170) <= 2291372;
srom_1(20171) <= 2699962;
srom_1(20172) <= 3135229;
srom_1(20173) <= 3595131;
srom_1(20174) <= 4077511;
srom_1(20175) <= 4580107;
srom_1(20176) <= 5100562;
srom_1(20177) <= 5636437;
srom_1(20178) <= 6185217;
srom_1(20179) <= 6744329;
srom_1(20180) <= 7311152;
srom_1(20181) <= 7883028;
srom_1(20182) <= 8457275;
srom_1(20183) <= 9031199;
srom_1(20184) <= 9602110;
srom_1(20185) <= 10167331;
srom_1(20186) <= 10724211;
srom_1(20187) <= 11270138;
srom_1(20188) <= 11802553;
srom_1(20189) <= 12318958;
srom_1(20190) <= 12816933;
srom_1(20191) <= 13294142;
srom_1(20192) <= 13748347;
srom_1(20193) <= 14177418;
srom_1(20194) <= 14579344;
srom_1(20195) <= 14952239;
srom_1(20196) <= 15294355;
srom_1(20197) <= 15604087;
srom_1(20198) <= 15879984;
srom_1(20199) <= 16120751;
srom_1(20200) <= 16325260;
srom_1(20201) <= 16492550;
srom_1(20202) <= 16621839;
srom_1(20203) <= 16712519;
srom_1(20204) <= 16764165;
srom_1(20205) <= 16776536;
srom_1(20206) <= 16749573;
srom_1(20207) <= 16683402;
srom_1(20208) <= 16578334;
srom_1(20209) <= 16434862;
srom_1(20210) <= 16253657;
srom_1(20211) <= 16035572;
srom_1(20212) <= 15781626;
srom_1(20213) <= 15493013;
srom_1(20214) <= 15171084;
srom_1(20215) <= 14817350;
srom_1(20216) <= 14433469;
srom_1(20217) <= 14021242;
srom_1(20218) <= 13582602;
srom_1(20219) <= 13119605;
srom_1(20220) <= 12634423;
srom_1(20221) <= 12129331;
srom_1(20222) <= 11606697;
srom_1(20223) <= 11068973;
srom_1(20224) <= 10518679;
srom_1(20225) <= 9958397;
srom_1(20226) <= 9390753;
srom_1(20227) <= 8818410;
srom_1(20228) <= 8244052;
srom_1(20229) <= 7670371;
srom_1(20230) <= 7100059;
srom_1(20231) <= 6535789;
srom_1(20232) <= 5980207;
srom_1(20233) <= 5435919;
srom_1(20234) <= 4905478;
srom_1(20235) <= 4391370;
srom_1(20236) <= 3896006;
srom_1(20237) <= 3421710;
srom_1(20238) <= 2970705;
srom_1(20239) <= 2545107;
srom_1(20240) <= 2146910;
srom_1(20241) <= 1777984;
srom_1(20242) <= 1440056;
srom_1(20243) <= 1134713;
srom_1(20244) <= 863386;
srom_1(20245) <= 627347;
srom_1(20246) <= 427704;
srom_1(20247) <= 265392;
srom_1(20248) <= 141172;
srom_1(20249) <= 55627;
srom_1(20250) <= 9159;
srom_1(20251) <= 1985;
srom_1(20252) <= 34138;
srom_1(20253) <= 105469;
srom_1(20254) <= 215642;
srom_1(20255) <= 364140;
srom_1(20256) <= 550269;
srom_1(20257) <= 773154;
srom_1(20258) <= 1031750;
srom_1(20259) <= 1324845;
srom_1(20260) <= 1651065;
srom_1(20261) <= 2008879;
srom_1(20262) <= 2396610;
srom_1(20263) <= 2812440;
srom_1(20264) <= 3254418;
srom_1(20265) <= 3720472;
srom_1(20266) <= 4208416;
srom_1(20267) <= 4715963;
srom_1(20268) <= 5240733;
srom_1(20269) <= 5780263;
srom_1(20270) <= 6332025;
srom_1(20271) <= 6893431;
srom_1(20272) <= 7461849;
srom_1(20273) <= 8034612;
srom_1(20274) <= 8609036;
srom_1(20275) <= 9182425;
srom_1(20276) <= 9752092;
srom_1(20277) <= 10315366;
srom_1(20278) <= 10869604;
srom_1(20279) <= 11412208;
srom_1(20280) <= 11940633;
srom_1(20281) <= 12452401;
srom_1(20282) <= 12945113;
srom_1(20283) <= 13416458;
srom_1(20284) <= 13864226;
srom_1(20285) <= 14286316;
srom_1(20286) <= 14680751;
srom_1(20287) <= 15045679;
srom_1(20288) <= 15379390;
srom_1(20289) <= 15680318;
srom_1(20290) <= 15947054;
srom_1(20291) <= 16178345;
srom_1(20292) <= 16373107;
srom_1(20293) <= 16530427;
srom_1(20294) <= 16649568;
srom_1(20295) <= 16729970;
srom_1(20296) <= 16771257;
srom_1(20297) <= 16773234;
srom_1(20298) <= 16735893;
srom_1(20299) <= 16659409;
srom_1(20300) <= 16544140;
srom_1(20301) <= 16390627;
srom_1(20302) <= 16199589;
srom_1(20303) <= 15971924;
srom_1(20304) <= 15708697;
srom_1(20305) <= 15411145;
srom_1(20306) <= 15080661;
srom_1(20307) <= 14718795;
srom_1(20308) <= 14327246;
srom_1(20309) <= 13907848;
srom_1(20310) <= 13462568;
srom_1(20311) <= 12993495;
srom_1(20312) <= 12502828;
srom_1(20313) <= 11992868;
srom_1(20314) <= 11466006;
srom_1(20315) <= 10924713;
srom_1(20316) <= 10371528;
srom_1(20317) <= 9809044;
srom_1(20318) <= 9239899;
srom_1(20319) <= 8666762;
srom_1(20320) <= 8092321;
srom_1(20321) <= 7519269;
srom_1(20322) <= 6950294;
srom_1(20323) <= 6388063;
srom_1(20324) <= 5835214;
srom_1(20325) <= 5294339;
srom_1(20326) <= 4767973;
srom_1(20327) <= 4258586;
srom_1(20328) <= 3768566;
srom_1(20329) <= 3300211;
srom_1(20330) <= 2855717;
srom_1(20331) <= 2437169;
srom_1(20332) <= 2046529;
srom_1(20333) <= 1685630;
srom_1(20334) <= 1356163;
srom_1(20335) <= 1059673;
srom_1(20336) <= 797551;
srom_1(20337) <= 571027;
srom_1(20338) <= 381162;
srom_1(20339) <= 228846;
srom_1(20340) <= 114794;
srom_1(20341) <= 39541;
srom_1(20342) <= 3440;
srom_1(20343) <= 6660;
srom_1(20344) <= 49185;
srom_1(20345) <= 130817;
srom_1(20346) <= 251172;
srom_1(20347) <= 409687;
srom_1(20348) <= 605618;
srom_1(20349) <= 838045;
srom_1(20350) <= 1105880;
srom_1(20351) <= 1407866;
srom_1(20352) <= 1742587;
srom_1(20353) <= 2108474;
srom_1(20354) <= 2503810;
srom_1(20355) <= 2926743;
srom_1(20356) <= 3375287;
srom_1(20357) <= 3847341;
srom_1(20358) <= 4340691;
srom_1(20359) <= 4853022;
srom_1(20360) <= 5381933;
srom_1(20361) <= 5924944;
srom_1(20362) <= 6479507;
srom_1(20363) <= 7043023;
srom_1(20364) <= 7612849;
srom_1(20365) <= 8186312;
srom_1(20366) <= 8760724;
srom_1(20367) <= 9333391;
srom_1(20368) <= 9901628;
srom_1(20369) <= 10462770;
srom_1(20370) <= 11014185;
srom_1(20371) <= 11553288;
srom_1(20372) <= 12077550;
srom_1(20373) <= 12584514;
srom_1(20374) <= 13071802;
srom_1(20375) <= 13537129;
srom_1(20376) <= 13978313;
srom_1(20377) <= 14393284;
srom_1(20378) <= 14780098;
srom_1(20379) <= 15136939;
srom_1(20380) <= 15462136;
srom_1(20381) <= 15754162;
srom_1(20382) <= 16011648;
srom_1(20383) <= 16233388;
srom_1(20384) <= 16418340;
srom_1(20385) <= 16565639;
srom_1(20386) <= 16674592;
srom_1(20387) <= 16744690;
srom_1(20388) <= 16775603;
srom_1(20389) <= 16767187;
srom_1(20390) <= 16719480;
srom_1(20391) <= 16632708;
srom_1(20392) <= 16507276;
srom_1(20393) <= 16343772;
srom_1(20394) <= 16142964;
srom_1(20395) <= 15905793;
srom_1(20396) <= 15633372;
srom_1(20397) <= 15326977;
srom_1(20398) <= 14988046;
srom_1(20399) <= 14618168;
srom_1(20400) <= 14219078;
srom_1(20401) <= 13792646;
srom_1(20402) <= 13340873;
srom_1(20403) <= 12865877;
srom_1(20404) <= 12369886;
srom_1(20405) <= 11855224;
srom_1(20406) <= 11324307;
srom_1(20407) <= 10779624;
srom_1(20408) <= 10223728;
srom_1(20409) <= 9659226;
srom_1(20410) <= 9088766;
srom_1(20411) <= 8515023;
srom_1(20412) <= 7940687;
srom_1(20413) <= 7368452;
srom_1(20414) <= 6801000;
srom_1(20415) <= 6240993;
srom_1(20416) <= 5691057;
srom_1(20417) <= 5153771;
srom_1(20418) <= 4631654;
srom_1(20419) <= 4127155;
srom_1(20420) <= 3642639;
srom_1(20421) <= 3180378;
srom_1(20422) <= 2742541;
srom_1(20423) <= 2331180;
srom_1(20424) <= 1948225;
srom_1(20425) <= 1595470;
srom_1(20426) <= 1274571;
srom_1(20427) <= 987032;
srom_1(20428) <= 734202;
srom_1(20429) <= 517266;
srom_1(20430) <= 337241;
srom_1(20431) <= 194972;
srom_1(20432) <= 91125;
srom_1(20433) <= 26188;
srom_1(20434) <= 466;
srom_1(20435) <= 14079;
srom_1(20436) <= 66962;
srom_1(20437) <= 158869;
srom_1(20438) <= 289367;
srom_1(20439) <= 457846;
srom_1(20440) <= 663515;
srom_1(20441) <= 905409;
srom_1(20442) <= 1182395;
srom_1(20443) <= 1493173;
srom_1(20444) <= 1836286;
srom_1(20445) <= 2210125;
srom_1(20446) <= 2612937;
srom_1(20447) <= 3042834;
srom_1(20448) <= 3497798;
srom_1(20449) <= 3975697;
srom_1(20450) <= 4474290;
srom_1(20451) <= 4991239;
srom_1(20452) <= 5524118;
srom_1(20453) <= 6070431;
srom_1(20454) <= 6627614;
srom_1(20455) <= 7193055;
srom_1(20456) <= 7764102;
srom_1(20457) <= 8338078;
srom_1(20458) <= 8912291;
srom_1(20459) <= 9484048;
srom_1(20460) <= 10050668;
srom_1(20461) <= 10609495;
srom_1(20462) <= 11157906;
srom_1(20463) <= 11693332;
srom_1(20464) <= 12213260;
srom_1(20465) <= 12715254;
srom_1(20466) <= 13196958;
srom_1(20467) <= 13656114;
srom_1(20468) <= 14090569;
srom_1(20469) <= 14498286;
srom_1(20470) <= 14877352;
srom_1(20471) <= 15225990;
srom_1(20472) <= 15542566;
srom_1(20473) <= 15825594;
srom_1(20474) <= 16073747;
srom_1(20475) <= 16285863;
srom_1(20476) <= 16460945;
srom_1(20477) <= 16598173;
srom_1(20478) <= 16696904;
srom_1(20479) <= 16756674;
srom_1(20480) <= 16777204;
srom_1(20481) <= 16758397;
srom_1(20482) <= 16700340;
srom_1(20483) <= 16603308;
srom_1(20484) <= 16467753;
srom_1(20485) <= 16294313;
srom_1(20486) <= 16083800;
srom_1(20487) <= 15837202;
srom_1(20488) <= 15555675;
srom_1(20489) <= 15240539;
srom_1(20490) <= 14893272;
srom_1(20491) <= 14515502;
srom_1(20492) <= 14109001;
srom_1(20493) <= 13675675;
srom_1(20494) <= 13217556;
srom_1(20495) <= 12736793;
srom_1(20496) <= 12235640;
srom_1(20497) <= 11716446;
srom_1(20498) <= 11181647;
srom_1(20499) <= 10633751;
srom_1(20500) <= 10075326;
srom_1(20501) <= 9508992;
srom_1(20502) <= 8937404;
srom_1(20503) <= 8363242;
srom_1(20504) <= 7789200;
srom_1(20505) <= 7217968;
srom_1(20506) <= 6652226;
srom_1(20507) <= 6094626;
srom_1(20508) <= 5547783;
srom_1(20509) <= 5014262;
srom_1(20510) <= 4496565;
srom_1(20511) <= 3997118;
srom_1(20512) <= 3518265;
srom_1(20513) <= 3062251;
srom_1(20514) <= 2631213;
srom_1(20515) <= 2227174;
srom_1(20516) <= 1852028;
srom_1(20517) <= 1507535;
srom_1(20518) <= 1195309;
srom_1(20519) <= 916815;
srom_1(20520) <= 673358;
srom_1(20521) <= 466081;
srom_1(20522) <= 295956;
srom_1(20523) <= 163780;
srom_1(20524) <= 70173;
srom_1(20525) <= 15574;
srom_1(20526) <= 238;
srom_1(20527) <= 24239;
srom_1(20528) <= 87463;
srom_1(20529) <= 189615;
srom_1(20530) <= 330214;
srom_1(20531) <= 508601;
srom_1(20532) <= 723941;
srom_1(20533) <= 975223;
srom_1(20534) <= 1261268;
srom_1(20535) <= 1580737;
srom_1(20536) <= 1932129;
srom_1(20537) <= 2313799;
srom_1(20538) <= 2723955;
srom_1(20539) <= 3160675;
srom_1(20540) <= 3621910;
srom_1(20541) <= 4105498;
srom_1(20542) <= 4609171;
srom_1(20543) <= 5130567;
srom_1(20544) <= 5667241;
srom_1(20545) <= 6216677;
srom_1(20546) <= 6776297;
srom_1(20547) <= 7343478;
srom_1(20548) <= 7915561;
srom_1(20549) <= 8489861;
srom_1(20550) <= 9063686;
srom_1(20551) <= 9634346;
srom_1(20552) <= 10199164;
srom_1(20553) <= 10755492;
srom_1(20554) <= 11300721;
srom_1(20555) <= 11832294;
srom_1(20556) <= 12347718;
srom_1(20557) <= 12844576;
srom_1(20558) <= 13320539;
srom_1(20559) <= 13773375;
srom_1(20560) <= 14200959;
srom_1(20561) <= 14601287;
srom_1(20562) <= 14972482;
srom_1(20563) <= 15312803;
srom_1(20564) <= 15620654;
srom_1(20565) <= 15894591;
srom_1(20566) <= 16133330;
srom_1(20567) <= 16335752;
srom_1(20568) <= 16500907;
srom_1(20569) <= 16628020;
srom_1(20570) <= 16716496;
srom_1(20571) <= 16765919;
srom_1(20572) <= 16776059;
srom_1(20573) <= 16746866;
srom_1(20574) <= 16678479;
srom_1(20575) <= 16571218;
srom_1(20576) <= 16425586;
srom_1(20577) <= 16242266;
srom_1(20578) <= 16022117;
srom_1(20579) <= 15766172;
srom_1(20580) <= 15475631;
srom_1(20581) <= 15151857;
srom_1(20582) <= 14796367;
srom_1(20583) <= 14410829;
srom_1(20584) <= 13997051;
srom_1(20585) <= 13556973;
srom_1(20586) <= 13092659;
srom_1(20587) <= 12606286;
srom_1(20588) <= 12100135;
srom_1(20589) <= 11576579;
srom_1(20590) <= 11038073;
srom_1(20591) <= 10487143;
srom_1(20592) <= 9926373;
srom_1(20593) <= 9358391;
srom_1(20594) <= 8785862;
srom_1(20595) <= 8211470;
srom_1(20596) <= 7637909;
srom_1(20597) <= 7067868;
srom_1(20598) <= 6504020;
srom_1(20599) <= 5949010;
srom_1(20600) <= 5405439;
srom_1(20601) <= 4875858;
srom_1(20602) <= 4362750;
srom_1(20603) <= 3868520;
srom_1(20604) <= 3395486;
srom_1(20605) <= 2945867;
srom_1(20606) <= 2521770;
srom_1(20607) <= 2125186;
srom_1(20608) <= 1757972;
srom_1(20609) <= 1421852;
srom_1(20610) <= 1118401;
srom_1(20611) <= 849043;
srom_1(20612) <= 615041;
srom_1(20613) <= 417491;
srom_1(20614) <= 257321;
srom_1(20615) <= 135281;
srom_1(20616) <= 51944;
srom_1(20617) <= 7700;
srom_1(20618) <= 2757;
srom_1(20619) <= 37138;
srom_1(20620) <= 110683;
srom_1(20621) <= 223045;
srom_1(20622) <= 373698;
srom_1(20623) <= 561936;
srom_1(20624) <= 786876;
srom_1(20625) <= 1047463;
srom_1(20626) <= 1342476;
srom_1(20627) <= 1670530;
srom_1(20628) <= 2030087;
srom_1(20629) <= 2419462;
srom_1(20630) <= 2836828;
srom_1(20631) <= 3280228;
srom_1(20632) <= 3747583;
srom_1(20633) <= 4236701;
srom_1(20634) <= 4745290;
srom_1(20635) <= 5270963;
srom_1(20636) <= 5811255;
srom_1(20637) <= 6363634;
srom_1(20638) <= 6925509;
srom_1(20639) <= 7494244;
srom_1(20640) <= 8067174;
srom_1(20641) <= 8641610;
srom_1(20642) <= 9214861;
srom_1(20643) <= 9784237;
srom_1(20644) <= 10347068;
srom_1(20645) <= 10900715;
srom_1(20646) <= 11442582;
srom_1(20647) <= 11970128;
srom_1(20648) <= 12480879;
srom_1(20649) <= 12972440;
srom_1(20650) <= 13442506;
srom_1(20651) <= 13888872;
srom_1(20652) <= 14309446;
srom_1(20653) <= 14702255;
srom_1(20654) <= 15065457;
srom_1(20655) <= 15397349;
srom_1(20656) <= 15696374;
srom_1(20657) <= 15961131;
srom_1(20658) <= 16190378;
srom_1(20659) <= 16383039;
srom_1(20660) <= 16538212;
srom_1(20661) <= 16655169;
srom_1(20662) <= 16733361;
srom_1(20663) <= 16772421;
srom_1(20664) <= 16772167;
srom_1(20665) <= 16732599;
srom_1(20666) <= 16653904;
srom_1(20667) <= 16536450;
srom_1(20668) <= 16380788;
srom_1(20669) <= 16187647;
srom_1(20670) <= 15957934;
srom_1(20671) <= 15692727;
srom_1(20672) <= 15393267;
srom_1(20673) <= 15060960;
srom_1(20674) <= 14697365;
srom_1(20675) <= 14304185;
srom_1(20676) <= 13883265;
srom_1(20677) <= 13436579;
srom_1(20678) <= 12966221;
srom_1(20679) <= 12474398;
srom_1(20680) <= 11963414;
srom_1(20681) <= 11435667;
srom_1(20682) <= 10893631;
srom_1(20683) <= 10339849;
srom_1(20684) <= 9776916;
srom_1(20685) <= 9207473;
srom_1(20686) <= 8634190;
srom_1(20687) <= 8059756;
srom_1(20688) <= 7486863;
srom_1(20689) <= 6918200;
srom_1(20690) <= 6356431;
srom_1(20691) <= 5804192;
srom_1(20692) <= 5264072;
srom_1(20693) <= 4738604;
srom_1(20694) <= 4230253;
srom_1(20695) <= 3741401;
srom_1(20696) <= 3274342;
srom_1(20697) <= 2831265;
srom_1(20698) <= 2414248;
srom_1(20699) <= 2025247;
srom_1(20700) <= 1666087;
srom_1(20701) <= 1338450;
srom_1(20702) <= 1043874;
srom_1(20703) <= 783740;
srom_1(20704) <= 559268;
srom_1(20705) <= 371510;
srom_1(20706) <= 221348;
srom_1(20707) <= 109484;
srom_1(20708) <= 36444;
srom_1(20709) <= 2570;
srom_1(20710) <= 8021;
srom_1(20711) <= 52772;
srom_1(20712) <= 136612;
srom_1(20713) <= 259148;
srom_1(20714) <= 419807;
srom_1(20715) <= 617834;
srom_1(20716) <= 852300;
srom_1(20717) <= 1122107;
srom_1(20718) <= 1425990;
srom_1(20719) <= 1762522;
srom_1(20720) <= 2130126;
srom_1(20721) <= 2527078;
srom_1(20722) <= 2951518;
srom_1(20723) <= 3401453;
srom_1(20724) <= 3874775;
srom_1(20725) <= 4369264;
srom_1(20726) <= 4882601;
srom_1(20727) <= 5412379;
srom_1(20728) <= 5956113;
srom_1(20729) <= 6511254;
srom_1(20730) <= 7075199;
srom_1(20731) <= 7645303;
srom_1(20732) <= 8218892;
srom_1(20733) <= 8793277;
srom_1(20734) <= 9365765;
srom_1(20735) <= 9933670;
srom_1(20736) <= 10494330;
srom_1(20737) <= 11045115;
srom_1(20738) <= 11583444;
srom_1(20739) <= 12106790;
srom_1(20740) <= 12612701;
srom_1(20741) <= 13098803;
srom_1(20742) <= 13562818;
srom_1(20743) <= 14002569;
srom_1(20744) <= 14415995;
srom_1(20745) <= 14801155;
srom_1(20746) <= 15156246;
srom_1(20747) <= 15479600;
srom_1(20748) <= 15769702;
srom_1(20749) <= 16025192;
srom_1(20750) <= 16244871;
srom_1(20751) <= 16427710;
srom_1(20752) <= 16572850;
srom_1(20753) <= 16679612;
srom_1(20754) <= 16747494;
srom_1(20755) <= 16776178;
srom_1(20756) <= 16765531;
srom_1(20757) <= 16715601;
srom_1(20758) <= 16626623;
srom_1(20759) <= 16499014;
srom_1(20760) <= 16333372;
srom_1(20761) <= 16130475;
srom_1(20762) <= 15891274;
srom_1(20763) <= 15616890;
srom_1(20764) <= 15308610;
srom_1(20765) <= 14967880;
srom_1(20766) <= 14596297;
srom_1(20767) <= 14195604;
srom_1(20768) <= 13767681;
srom_1(20769) <= 13314533;
srom_1(20770) <= 12838285;
srom_1(20771) <= 12341172;
srom_1(20772) <= 11825523;
srom_1(20773) <= 11293758;
srom_1(20774) <= 10748370;
srom_1(20775) <= 10191915;
srom_1(20776) <= 9627005;
srom_1(20777) <= 9056287;
srom_1(20778) <= 8482438;
srom_1(20779) <= 7908149;
srom_1(20780) <= 7336113;
srom_1(20781) <= 6769013;
srom_1(20782) <= 6209508;
srom_1(20783) <= 5660221;
srom_1(20784) <= 5123728;
srom_1(20785) <= 4602545;
srom_1(20786) <= 4099117;
srom_1(20787) <= 3615804;
srom_1(20788) <= 3154872;
srom_1(20789) <= 2718482;
srom_1(20790) <= 2308682;
srom_1(20791) <= 1927393;
srom_1(20792) <= 1576402;
srom_1(20793) <= 1257356;
srom_1(20794) <= 971752;
srom_1(20795) <= 720927;
srom_1(20796) <= 506059;
srom_1(20797) <= 328154;
srom_1(20798) <= 188048;
srom_1(20799) <= 86397;
srom_1(20800) <= 23679;
srom_1(20801) <= 186;
srom_1(20802) <= 16029;
srom_1(20803) <= 71134;
srom_1(20804) <= 165243;
srom_1(20805) <= 297914;
srom_1(20806) <= 468525;
srom_1(20807) <= 676275;
srom_1(20808) <= 920192;
srom_1(20809) <= 1199131;
srom_1(20810) <= 1511783;
srom_1(20811) <= 1856683;
srom_1(20812) <= 2232214;
srom_1(20813) <= 2636614;
srom_1(20814) <= 3067988;
srom_1(20815) <= 3524311;
srom_1(20816) <= 4003445;
srom_1(20817) <= 4503142;
srom_1(20818) <= 5021060;
srom_1(20819) <= 5554769;
srom_1(20820) <= 6101767;
srom_1(20821) <= 6659489;
srom_1(20822) <= 7225319;
srom_1(20823) <= 7796604;
srom_1(20824) <= 8370666;
srom_1(20825) <= 8944811;
srom_1(20826) <= 9516349;
srom_1(20827) <= 10082597;
srom_1(20828) <= 10640903;
srom_1(20829) <= 11188646;
srom_1(20830) <= 11723259;
srom_1(20831) <= 12242235;
srom_1(20832) <= 12743140;
srom_1(20833) <= 13223625;
srom_1(20834) <= 13681436;
srom_1(20835) <= 14114428;
srom_1(20836) <= 14520570;
srom_1(20837) <= 14897956;
srom_1(20838) <= 15244819;
srom_1(20839) <= 15559529;
srom_1(20840) <= 15840613;
srom_1(20841) <= 16086753;
srom_1(20842) <= 16296792;
srom_1(20843) <= 16469748;
srom_1(20844) <= 16604808;
srom_1(20845) <= 16701340;
srom_1(20846) <= 16758890;
srom_1(20847) <= 16777190;
srom_1(20848) <= 16756152;
srom_1(20849) <= 16695876;
srom_1(20850) <= 16596645;
srom_1(20851) <= 16458923;
srom_1(20852) <= 16283356;
srom_1(20853) <= 16070769;
srom_1(20854) <= 15822157;
srom_1(20855) <= 15538687;
srom_1(20856) <= 15221687;
srom_1(20857) <= 14872645;
srom_1(20858) <= 14493197;
srom_1(20859) <= 14085122;
srom_1(20860) <= 13650335;
srom_1(20861) <= 13190873;
srom_1(20862) <= 12708892;
srom_1(20863) <= 12206652;
srom_1(20864) <= 11686507;
srom_1(20865) <= 11150898;
srom_1(20866) <= 10602335;
srom_1(20867) <= 10043392;
srom_1(20868) <= 9476688;
srom_1(20869) <= 8904882;
srom_1(20870) <= 8330655;
srom_1(20871) <= 7756700;
srom_1(20872) <= 7185708;
srom_1(20873) <= 6620357;
srom_1(20874) <= 6063297;
srom_1(20875) <= 5517142;
srom_1(20876) <= 4984453;
srom_1(20877) <= 4467726;
srom_1(20878) <= 3969386;
srom_1(20879) <= 3491769;
srom_1(20880) <= 3037115;
srom_1(20881) <= 2607556;
srom_1(20882) <= 2205106;
srom_1(20883) <= 1831653;
srom_1(20884) <= 1488948;
srom_1(20885) <= 1178598;
srom_1(20886) <= 902057;
srom_1(20887) <= 660624;
srom_1(20888) <= 455430;
srom_1(20889) <= 287437;
srom_1(20890) <= 157434;
srom_1(20891) <= 66029;
srom_1(20892) <= 13652;
srom_1(20893) <= 548;
srom_1(20894) <= 26778;
srom_1(20895) <= 92220;
srom_1(20896) <= 196566;
srom_1(20897) <= 339328;
srom_1(20898) <= 519835;
srom_1(20899) <= 737242;
srom_1(20900) <= 990529;
srom_1(20901) <= 1278508;
srom_1(20902) <= 1599828;
srom_1(20903) <= 1952984;
srom_1(20904) <= 2336318;
srom_1(20905) <= 2748033;
srom_1(20906) <= 3186200;
srom_1(20907) <= 3648762;
srom_1(20908) <= 4133550;
srom_1(20909) <= 4638293;
srom_1(20910) <= 5160621;
srom_1(20911) <= 5698087;
srom_1(20912) <= 6248170;
srom_1(20913) <= 6808290;
srom_1(20914) <= 7375820;
srom_1(20915) <= 7948100;
srom_1(20916) <= 8522445;
srom_1(20917) <= 9096163;
srom_1(20918) <= 9666563;
srom_1(20919) <= 10230970;
srom_1(20920) <= 10786738;
srom_1(20921) <= 11331260;
srom_1(20922) <= 11861983;
srom_1(20923) <= 12376418;
srom_1(20924) <= 12872153;
srom_1(20925) <= 13346863;
srom_1(20926) <= 13798322;
srom_1(20927) <= 14224413;
srom_1(20928) <= 14623137;
srom_1(20929) <= 14992626;
srom_1(20930) <= 15331147;
srom_1(20931) <= 15637111;
srom_1(20932) <= 15909085;
srom_1(20933) <= 16145793;
srom_1(20934) <= 16346124;
srom_1(20935) <= 16509140;
srom_1(20936) <= 16634076;
srom_1(20937) <= 16720347;
srom_1(20938) <= 16767546;
srom_1(20939) <= 16775455;
srom_1(20940) <= 16744034;
srom_1(20941) <= 16673432;
srom_1(20942) <= 16563979;
srom_1(20943) <= 16416189;
srom_1(20944) <= 16230755;
srom_1(20945) <= 16008547;
srom_1(20946) <= 15750606;
srom_1(20947) <= 15458142;
srom_1(20948) <= 15132527;
srom_1(20949) <= 14775287;
srom_1(20950) <= 14388098;
srom_1(20951) <= 13972775;
srom_1(20952) <= 13531266;
srom_1(20953) <= 13065642;
srom_1(20954) <= 12578085;
srom_1(20955) <= 12070882;
srom_1(20956) <= 11546412;
srom_1(20957) <= 11007133;
srom_1(20958) <= 10455576;
srom_1(20959) <= 9894326;
srom_1(20960) <= 9326015;
srom_1(20961) <= 8753308;
srom_1(20962) <= 8178891;
srom_1(20963) <= 7605457;
srom_1(20964) <= 7035696;
srom_1(20965) <= 6472279;
srom_1(20966) <= 5917849;
srom_1(20967) <= 5375004;
srom_1(20968) <= 4846292;
srom_1(20969) <= 4334190;
srom_1(20970) <= 3841102;
srom_1(20971) <= 3369338;
srom_1(20972) <= 2921111;
srom_1(20973) <= 2498523;
srom_1(20974) <= 2103555;
srom_1(20975) <= 1738061;
srom_1(20976) <= 1403753;
srom_1(20977) <= 1102199;
srom_1(20978) <= 834814;
srom_1(20979) <= 602851;
srom_1(20980) <= 407399;
srom_1(20981) <= 249373;
srom_1(20982) <= 129514;
srom_1(20983) <= 48386;
srom_1(20984) <= 6367;
srom_1(20985) <= 3656;
srom_1(20986) <= 40264;
srom_1(20987) <= 116021;
srom_1(20988) <= 230571;
srom_1(20989) <= 383377;
srom_1(20990) <= 573722;
srom_1(20991) <= 800713;
srom_1(20992) <= 1063287;
srom_1(20993) <= 1360212;
srom_1(20994) <= 1690096;
srom_1(20995) <= 2051391;
srom_1(20996) <= 2442403;
srom_1(20997) <= 2861299;
srom_1(20998) <= 3306115;
srom_1(20999) <= 3774764;
srom_1(21000) <= 4265049;
srom_1(21001) <= 4774671;
srom_1(21002) <= 5301240;
srom_1(21003) <= 5842286;
srom_1(21004) <= 6395273;
srom_1(21005) <= 6957608;
srom_1(21006) <= 7526653;
srom_1(21007) <= 8099740;
srom_1(21008) <= 8674181;
srom_1(21009) <= 9247284;
srom_1(21010) <= 9816360;
srom_1(21011) <= 10378740;
srom_1(21012) <= 10931788;
srom_1(21013) <= 11472911;
srom_1(21014) <= 11999570;
srom_1(21015) <= 12509295;
srom_1(21016) <= 12999698;
srom_1(21017) <= 13468478;
srom_1(21018) <= 13913436;
srom_1(21019) <= 14332486;
srom_1(21020) <= 14723664;
srom_1(21021) <= 15085134;
srom_1(21022) <= 15415202;
srom_1(21023) <= 15712320;
srom_1(21024) <= 15975095;
srom_1(21025) <= 16202293;
srom_1(21026) <= 16392851;
srom_1(21027) <= 16545874;
srom_1(21028) <= 16660645;
srom_1(21029) <= 16736626;
srom_1(21030) <= 16773459;
srom_1(21031) <= 16770974;
srom_1(21032) <= 16729180;
srom_1(21033) <= 16648275;
srom_1(21034) <= 16528637;
srom_1(21035) <= 16370828;
srom_1(21036) <= 16175587;
srom_1(21037) <= 15943831;
srom_1(21038) <= 15676645;
srom_1(21039) <= 15375284;
srom_1(21040) <= 15041159;
srom_1(21041) <= 14675839;
srom_1(21042) <= 14281035;
srom_1(21043) <= 13858600;
srom_1(21044) <= 13410514;
srom_1(21045) <= 12938879;
srom_1(21046) <= 12445906;
srom_1(21047) <= 11933907;
srom_1(21048) <= 11405282;
srom_1(21049) <= 10862512;
srom_1(21050) <= 10308140;
srom_1(21051) <= 9744767;
srom_1(21052) <= 9175035;
srom_1(21053) <= 8601615;
srom_1(21054) <= 8027196;
srom_1(21055) <= 7454471;
srom_1(21056) <= 6886127;
srom_1(21057) <= 6324829;
srom_1(21058) <= 5773209;
srom_1(21059) <= 5233853;
srom_1(21060) <= 4709291;
srom_1(21061) <= 4201982;
srom_1(21062) <= 3714306;
srom_1(21063) <= 3248549;
srom_1(21064) <= 2806896;
srom_1(21065) <= 2391417;
srom_1(21066) <= 2004062;
srom_1(21067) <= 1646645;
srom_1(21068) <= 1320844;
srom_1(21069) <= 1028186;
srom_1(21070) <= 770044;
srom_1(21071) <= 547627;
srom_1(21072) <= 361980;
srom_1(21073) <= 213973;
srom_1(21074) <= 104299;
srom_1(21075) <= 33473;
srom_1(21076) <= 1827;
srom_1(21077) <= 9509;
srom_1(21078) <= 56484;
srom_1(21079) <= 142531;
srom_1(21080) <= 267247;
srom_1(21081) <= 430047;
srom_1(21082) <= 630167;
srom_1(21083) <= 866669;
srom_1(21084) <= 1138444;
srom_1(21085) <= 1444218;
srom_1(21086) <= 1782556;
srom_1(21087) <= 2151872;
srom_1(21088) <= 2550435;
srom_1(21089) <= 2976374;
srom_1(21090) <= 3427694;
srom_1(21091) <= 3902277;
srom_1(21092) <= 4397898;
srom_1(21093) <= 4912232;
srom_1(21094) <= 5442869;
srom_1(21095) <= 5987319;
srom_1(21096) <= 6543029;
srom_1(21097) <= 7107395;
srom_1(21098) <= 7677768;
srom_1(21099) <= 8251474;
srom_1(21100) <= 8825824;
srom_1(21101) <= 9398123;
srom_1(21102) <= 9965688;
srom_1(21103) <= 10525858;
srom_1(21104) <= 11076006;
srom_1(21105) <= 11613551;
srom_1(21106) <= 12135974;
srom_1(21107) <= 12640824;
srom_1(21108) <= 13125734;
srom_1(21109) <= 13588429;
srom_1(21110) <= 14026741;
srom_1(21111) <= 14438614;
srom_1(21112) <= 14822116;
srom_1(21113) <= 15175450;
srom_1(21114) <= 15496957;
srom_1(21115) <= 15785131;
srom_1(21116) <= 16038620;
srom_1(21117) <= 16256236;
srom_1(21118) <= 16436957;
srom_1(21119) <= 16579938;
srom_1(21120) <= 16684506;
srom_1(21121) <= 16750171;
srom_1(21122) <= 16776627;
srom_1(21123) <= 16763748;
srom_1(21124) <= 16711596;
srom_1(21125) <= 16620414;
srom_1(21126) <= 16490630;
srom_1(21127) <= 16322853;
srom_1(21128) <= 16117869;
srom_1(21129) <= 15876641;
srom_1(21130) <= 15600298;
srom_1(21131) <= 15290138;
srom_1(21132) <= 14947614;
srom_1(21133) <= 14574332;
srom_1(21134) <= 14172043;
srom_1(21135) <= 13742634;
srom_1(21136) <= 13288118;
srom_1(21137) <= 12810626;
srom_1(21138) <= 12312398;
srom_1(21139) <= 11795770;
srom_1(21140) <= 11263165;
srom_1(21141) <= 10717080;
srom_1(21142) <= 10160076;
srom_1(21143) <= 9594765;
srom_1(21144) <= 9023797;
srom_1(21145) <= 8449852;
srom_1(21146) <= 7875619;
srom_1(21147) <= 7303791;
srom_1(21148) <= 6737051;
srom_1(21149) <= 6178055;
srom_1(21150) <= 5629425;
srom_1(21151) <= 5093734;
srom_1(21152) <= 4573494;
srom_1(21153) <= 4071144;
srom_1(21154) <= 3589041;
srom_1(21155) <= 3129444;
srom_1(21156) <= 2694509;
srom_1(21157) <= 2286276;
srom_1(21158) <= 1906658;
srom_1(21159) <= 1557437;
srom_1(21160) <= 1240249;
srom_1(21161) <= 956583;
srom_1(21162) <= 707768;
srom_1(21163) <= 494971;
srom_1(21164) <= 319190;
srom_1(21165) <= 181249;
srom_1(21166) <= 81795;
srom_1(21167) <= 21295;
srom_1(21168) <= 32;
srom_1(21169) <= 18106;
srom_1(21170) <= 75432;
srom_1(21171) <= 171741;
srom_1(21172) <= 306582;
srom_1(21173) <= 479323;
srom_1(21174) <= 689152;
srom_1(21175) <= 935088;
srom_1(21176) <= 1215975;
srom_1(21177) <= 1530497;
srom_1(21178) <= 1877180;
srom_1(21179) <= 2254396;
srom_1(21180) <= 2660378;
srom_1(21181) <= 3093222;
srom_1(21182) <= 3550897;
srom_1(21183) <= 4031258;
srom_1(21184) <= 4532053;
srom_1(21185) <= 5050932;
srom_1(21186) <= 5585462;
srom_1(21187) <= 6133138;
srom_1(21188) <= 6691390;
srom_1(21189) <= 7257601;
srom_1(21190) <= 7829115;
srom_1(21191) <= 8403254;
srom_1(21192) <= 8977323;
srom_1(21193) <= 9548632;
srom_1(21194) <= 10114501;
srom_1(21195) <= 10672277;
srom_1(21196) <= 11219344;
srom_1(21197) <= 11753136;
srom_1(21198) <= 12271151;
srom_1(21199) <= 12770960;
srom_1(21200) <= 13250218;
srom_1(21201) <= 13706679;
srom_1(21202) <= 14138201;
srom_1(21203) <= 14542761;
srom_1(21204) <= 14918462;
srom_1(21205) <= 15263543;
srom_1(21206) <= 15576385;
srom_1(21207) <= 15855521;
srom_1(21208) <= 16099641;
srom_1(21209) <= 16307603;
srom_1(21210) <= 16478429;
srom_1(21211) <= 16611319;
srom_1(21212) <= 16705650;
srom_1(21213) <= 16760980;
srom_1(21214) <= 16777049;
srom_1(21215) <= 16753781;
srom_1(21216) <= 16691286;
srom_1(21217) <= 16589858;
srom_1(21218) <= 16449970;
srom_1(21219) <= 16272280;
srom_1(21220) <= 16057621;
srom_1(21221) <= 15807000;
srom_1(21222) <= 15521590;
srom_1(21223) <= 15202732;
srom_1(21224) <= 14851920;
srom_1(21225) <= 14470800;
srom_1(21226) <= 14061158;
srom_1(21227) <= 13624915;
srom_1(21228) <= 13164118;
srom_1(21229) <= 12680926;
srom_1(21230) <= 12177606;
srom_1(21231) <= 11656519;
srom_1(21232) <= 11120107;
srom_1(21233) <= 10570886;
srom_1(21234) <= 10011432;
srom_1(21235) <= 9444367;
srom_1(21236) <= 8872352;
srom_1(21237) <= 8298068;
srom_1(21238) <= 7724209;
srom_1(21239) <= 7153466;
srom_1(21240) <= 6588515;
srom_1(21241) <= 6032004;
srom_1(21242) <= 5486545;
srom_1(21243) <= 4954694;
srom_1(21244) <= 4438947;
srom_1(21245) <= 3941720;
srom_1(21246) <= 3465347;
srom_1(21247) <= 3012060;
srom_1(21248) <= 2583986;
srom_1(21249) <= 2183132;
srom_1(21250) <= 1811377;
srom_1(21251) <= 1470465;
srom_1(21252) <= 1161995;
srom_1(21253) <= 887413;
srom_1(21254) <= 648007;
srom_1(21255) <= 444898;
srom_1(21256) <= 279041;
srom_1(21257) <= 151212;
srom_1(21258) <= 62011;
srom_1(21259) <= 11857;
srom_1(21260) <= 983;
srom_1(21261) <= 29443;
srom_1(21262) <= 97101;
srom_1(21263) <= 203641;
srom_1(21264) <= 348563;
srom_1(21265) <= 531188;
srom_1(21266) <= 750659;
srom_1(21267) <= 1005946;
srom_1(21268) <= 1295854;
srom_1(21269) <= 1619022;
srom_1(21270) <= 1973935;
srom_1(21271) <= 2358928;
srom_1(21272) <= 2772197;
srom_1(21273) <= 3211803;
srom_1(21274) <= 3675684;
srom_1(21275) <= 4161667;
srom_1(21276) <= 4667471;
srom_1(21277) <= 5190724;
srom_1(21278) <= 5728974;
srom_1(21279) <= 6279695;
srom_1(21280) <= 6840306;
srom_1(21281) <= 7408177;
srom_1(21282) <= 7980646;
srom_1(21283) <= 8555028;
srom_1(21284) <= 9128630;
srom_1(21285) <= 9698761;
srom_1(21286) <= 10262749;
srom_1(21287) <= 10817948;
srom_1(21288) <= 11361755;
srom_1(21289) <= 11891620;
srom_1(21290) <= 12405058;
srom_1(21291) <= 12899661;
srom_1(21292) <= 13373111;
srom_1(21293) <= 13823187;
srom_1(21294) <= 14247778;
srom_1(21295) <= 14644893;
srom_1(21296) <= 15012671;
srom_1(21297) <= 15349386;
srom_1(21298) <= 15653459;
srom_1(21299) <= 15923465;
srom_1(21300) <= 16158138;
srom_1(21301) <= 16356377;
srom_1(21302) <= 16517252;
srom_1(21303) <= 16640008;
srom_1(21304) <= 16724072;
srom_1(21305) <= 16769047;
srom_1(21306) <= 16774724;
srom_1(21307) <= 16741075;
srom_1(21308) <= 16668259;
srom_1(21309) <= 16556616;
srom_1(21310) <= 16406671;
srom_1(21311) <= 16219127;
srom_1(21312) <= 15994862;
srom_1(21313) <= 15734929;
srom_1(21314) <= 15440547;
srom_1(21315) <= 15113096;
srom_1(21316) <= 14754111;
srom_1(21317) <= 14365276;
srom_1(21318) <= 13948415;
srom_1(21319) <= 13505482;
srom_1(21320) <= 13038554;
srom_1(21321) <= 12549821;
srom_1(21322) <= 12041574;
srom_1(21323) <= 11516197;
srom_1(21324) <= 10976154;
srom_1(21325) <= 10423977;
srom_1(21326) <= 9862256;
srom_1(21327) <= 9293624;
srom_1(21328) <= 8720748;
srom_1(21329) <= 8146315;
srom_1(21330) <= 7573018;
srom_1(21331) <= 7003545;
srom_1(21332) <= 6440568;
srom_1(21333) <= 5886725;
srom_1(21334) <= 5344615;
srom_1(21335) <= 4816779;
srom_1(21336) <= 4305692;
srom_1(21337) <= 3813752;
srom_1(21338) <= 3343265;
srom_1(21339) <= 2896437;
srom_1(21340) <= 2475364;
srom_1(21341) <= 2082020;
srom_1(21342) <= 1718249;
srom_1(21343) <= 1385759;
srom_1(21344) <= 1086107;
srom_1(21345) <= 820699;
srom_1(21346) <= 590779;
srom_1(21347) <= 397427;
srom_1(21348) <= 241547;
srom_1(21349) <= 123872;
srom_1(21350) <= 44953;
srom_1(21351) <= 5161;
srom_1(21352) <= 4681;
srom_1(21353) <= 43517;
srom_1(21354) <= 121485;
srom_1(21355) <= 238221;
srom_1(21356) <= 393176;
srom_1(21357) <= 585625;
srom_1(21358) <= 814665;
srom_1(21359) <= 1079222;
srom_1(21360) <= 1378055;
srom_1(21361) <= 1709763;
srom_1(21362) <= 2072790;
srom_1(21363) <= 2465434;
srom_1(21364) <= 2885854;
srom_1(21365) <= 3332078;
srom_1(21366) <= 3802015;
srom_1(21367) <= 4293459;
srom_1(21368) <= 4804107;
srom_1(21369) <= 5331563;
srom_1(21370) <= 5873356;
srom_1(21371) <= 6426943;
srom_1(21372) <= 6989729;
srom_1(21373) <= 7559075;
srom_1(21374) <= 8132310;
srom_1(21375) <= 8706748;
srom_1(21376) <= 9279694;
srom_1(21377) <= 9848461;
srom_1(21378) <= 10410383;
srom_1(21379) <= 10962823;
srom_1(21380) <= 11503192;
srom_1(21381) <= 12028956;
srom_1(21382) <= 12537649;
srom_1(21383) <= 13026886;
srom_1(21384) <= 13494372;
srom_1(21385) <= 13937916;
srom_1(21386) <= 14355437;
srom_1(21387) <= 14744977;
srom_1(21388) <= 15104710;
srom_1(21389) <= 15432950;
srom_1(21390) <= 15728155;
srom_1(21391) <= 15988943;
srom_1(21392) <= 16214091;
srom_1(21393) <= 16402542;
srom_1(21394) <= 16553413;
srom_1(21395) <= 16665996;
srom_1(21396) <= 16739764;
srom_1(21397) <= 16774371;
srom_1(21398) <= 16769654;
srom_1(21399) <= 16725635;
srom_1(21400) <= 16642521;
srom_1(21401) <= 16520701;
srom_1(21402) <= 16360747;
srom_1(21403) <= 16163410;
srom_1(21404) <= 15929613;
srom_1(21405) <= 15660454;
srom_1(21406) <= 15357195;
srom_1(21407) <= 15021258;
srom_1(21408) <= 14654218;
srom_1(21409) <= 14257796;
srom_1(21410) <= 13833852;
srom_1(21411) <= 13384373;
srom_1(21412) <= 12911468;
srom_1(21413) <= 12417353;
srom_1(21414) <= 11904346;
srom_1(21415) <= 11374852;
srom_1(21416) <= 10831355;
srom_1(21417) <= 10276403;
srom_1(21418) <= 9712598;
srom_1(21419) <= 9142585;
srom_1(21420) <= 8569036;
srom_1(21421) <= 7994641;
srom_1(21422) <= 7422093;
srom_1(21423) <= 6854078;
srom_1(21424) <= 6293259;
srom_1(21425) <= 5742265;
srom_1(21426) <= 5203681;
srom_1(21427) <= 4680033;
srom_1(21428) <= 4173775;
srom_1(21429) <= 3687282;
srom_1(21430) <= 3222835;
srom_1(21431) <= 2782612;
srom_1(21432) <= 2368677;
srom_1(21433) <= 1982972;
srom_1(21434) <= 1627305;
srom_1(21435) <= 1303345;
srom_1(21436) <= 1012609;
srom_1(21437) <= 756462;
srom_1(21438) <= 536105;
srom_1(21439) <= 352571;
srom_1(21440) <= 206721;
srom_1(21441) <= 99238;
srom_1(21442) <= 30627;
srom_1(21443) <= 1210;
srom_1(21444) <= 11124;
srom_1(21445) <= 60322;
srom_1(21446) <= 148575;
srom_1(21447) <= 275469;
srom_1(21448) <= 440407;
srom_1(21449) <= 642618;
srom_1(21450) <= 881152;
srom_1(21451) <= 1154891;
srom_1(21452) <= 1462551;
srom_1(21453) <= 1802690;
srom_1(21454) <= 2173713;
srom_1(21455) <= 2573879;
srom_1(21456) <= 3001313;
srom_1(21457) <= 3454010;
srom_1(21458) <= 3929846;
srom_1(21459) <= 4426592;
srom_1(21460) <= 4941916;
srom_1(21461) <= 5473403;
srom_1(21462) <= 6018561;
srom_1(21463) <= 6574833;
srom_1(21464) <= 7139610;
srom_1(21465) <= 7710244;
srom_1(21466) <= 8284059;
srom_1(21467) <= 8858364;
srom_1(21468) <= 9430466;
srom_1(21469) <= 9997683;
srom_1(21470) <= 10557355;
srom_1(21471) <= 11106856;
srom_1(21472) <= 11643610;
srom_1(21473) <= 12165101;
srom_1(21474) <= 12668882;
srom_1(21475) <= 13152592;
srom_1(21476) <= 13613962;
srom_1(21477) <= 14050828;
srom_1(21478) <= 14461142;
srom_1(21479) <= 14842980;
srom_1(21480) <= 15194551;
srom_1(21481) <= 15514207;
srom_1(21482) <= 15800448;
srom_1(21483) <= 16051933;
srom_1(21484) <= 16267482;
srom_1(21485) <= 16446084;
srom_1(21486) <= 16586901;
srom_1(21487) <= 16689275;
srom_1(21488) <= 16752723;
srom_1(21489) <= 16776949;
srom_1(21490) <= 16761839;
srom_1(21491) <= 16707465;
srom_1(21492) <= 16614080;
srom_1(21493) <= 16482124;
srom_1(21494) <= 16312214;
srom_1(21495) <= 16105147;
srom_1(21496) <= 15861895;
srom_1(21497) <= 15583598;
srom_1(21498) <= 15271562;
srom_1(21499) <= 14927249;
srom_1(21500) <= 14552273;
srom_1(21501) <= 14148395;
srom_1(21502) <= 13717507;
srom_1(21503) <= 13261629;
srom_1(21504) <= 12782901;
srom_1(21505) <= 12283566;
srom_1(21506) <= 11765966;
srom_1(21507) <= 11232529;
srom_1(21508) <= 10685755;
srom_1(21509) <= 10128210;
srom_1(21510) <= 9562507;
srom_1(21511) <= 8991299;
srom_1(21512) <= 8417264;
srom_1(21513) <= 7843096;
srom_1(21514) <= 7271485;
srom_1(21515) <= 6705113;
srom_1(21516) <= 6146636;
srom_1(21517) <= 5598672;
srom_1(21518) <= 5063790;
srom_1(21519) <= 4544501;
srom_1(21520) <= 4043237;
srom_1(21521) <= 3562350;
srom_1(21522) <= 3104096;
srom_1(21523) <= 2670622;
srom_1(21524) <= 2263961;
srom_1(21525) <= 1886022;
srom_1(21526) <= 1538575;
srom_1(21527) <= 1223250;
srom_1(21528) <= 941527;
srom_1(21529) <= 694725;
srom_1(21530) <= 484002;
srom_1(21531) <= 310347;
srom_1(21532) <= 174573;
srom_1(21533) <= 77318;
srom_1(21534) <= 19037;
srom_1(21535) <= 5;
srom_1(21536) <= 20309;
srom_1(21537) <= 79855;
srom_1(21538) <= 178364;
srom_1(21539) <= 315373;
srom_1(21540) <= 490240;
srom_1(21541) <= 702146;
srom_1(21542) <= 950096;
srom_1(21543) <= 1232928;
srom_1(21544) <= 1549315;
srom_1(21545) <= 1897774;
srom_1(21546) <= 2276671;
srom_1(21547) <= 2684228;
srom_1(21548) <= 3118536;
srom_1(21549) <= 3577557;
srom_1(21550) <= 4059138;
srom_1(21551) <= 4561022;
srom_1(21552) <= 5080854;
srom_1(21553) <= 5616198;
srom_1(21554) <= 6164542;
srom_1(21555) <= 6723316;
srom_1(21556) <= 7289899;
srom_1(21557) <= 7861635;
srom_1(21558) <= 8435841;
srom_1(21559) <= 9009826;
srom_1(21560) <= 9580898;
srom_1(21561) <= 10146379;
srom_1(21562) <= 10703617;
srom_1(21563) <= 11249999;
srom_1(21564) <= 11782963;
srom_1(21565) <= 12300009;
srom_1(21566) <= 12798714;
srom_1(21567) <= 13276738;
srom_1(21568) <= 13731841;
srom_1(21569) <= 14161887;
srom_1(21570) <= 14564860;
srom_1(21571) <= 14938870;
srom_1(21572) <= 15282164;
srom_1(21573) <= 15593132;
srom_1(21574) <= 15870315;
srom_1(21575) <= 16112414;
srom_1(21576) <= 16318293;
srom_1(21577) <= 16486988;
srom_1(21578) <= 16617706;
srom_1(21579) <= 16709835;
srom_1(21580) <= 16762943;
srom_1(21581) <= 16776781;
srom_1(21582) <= 16751284;
srom_1(21583) <= 16686571;
srom_1(21584) <= 16582947;
srom_1(21585) <= 16440896;
srom_1(21586) <= 16261086;
srom_1(21587) <= 16044358;
srom_1(21588) <= 15791730;
srom_1(21589) <= 15504387;
srom_1(21590) <= 15183675;
srom_1(21591) <= 14831098;
srom_1(21592) <= 14448311;
srom_1(21593) <= 14037108;
srom_1(21594) <= 13599416;
srom_1(21595) <= 13137290;
srom_1(21596) <= 12652895;
srom_1(21597) <= 12148504;
srom_1(21598) <= 11626481;
srom_1(21599) <= 11089275;
srom_1(21600) <= 10539404;
srom_1(21601) <= 9979447;
srom_1(21602) <= 9412031;
srom_1(21603) <= 8839815;
srom_1(21604) <= 8265483;
srom_1(21605) <= 7691729;
srom_1(21606) <= 7121243;
srom_1(21607) <= 6556699;
srom_1(21608) <= 6000747;
srom_1(21609) <= 5455991;
srom_1(21610) <= 4924988;
srom_1(21611) <= 4410227;
srom_1(21612) <= 3914122;
srom_1(21613) <= 3438999;
srom_1(21614) <= 2987087;
srom_1(21615) <= 2560504;
srom_1(21616) <= 2161251;
srom_1(21617) <= 1791200;
srom_1(21618) <= 1452087;
srom_1(21619) <= 1145502;
srom_1(21620) <= 872882;
srom_1(21621) <= 635506;
srom_1(21622) <= 434487;
srom_1(21623) <= 270767;
srom_1(21624) <= 145115;
srom_1(21625) <= 58119;
srom_1(21626) <= 10188;
srom_1(21627) <= 1546;
srom_1(21628) <= 32234;
srom_1(21629) <= 102108;
srom_1(21630) <= 210840;
srom_1(21631) <= 357920;
srom_1(21632) <= 542659;
srom_1(21633) <= 764191;
srom_1(21634) <= 1021475;
srom_1(21635) <= 1313307;
srom_1(21636) <= 1638318;
srom_1(21637) <= 1994983;
srom_1(21638) <= 2381629;
srom_1(21639) <= 2796445;
srom_1(21640) <= 3237484;
srom_1(21641) <= 3702678;
srom_1(21642) <= 4189847;
srom_1(21643) <= 4696705;
srom_1(21644) <= 5220875;
srom_1(21645) <= 5759900;
srom_1(21646) <= 6311252;
srom_1(21647) <= 6872345;
srom_1(21648) <= 7440549;
srom_1(21649) <= 8013198;
srom_1(21650) <= 8587608;
srom_1(21651) <= 9161085;
srom_1(21652) <= 9730939;
srom_1(21653) <= 10294498;
srom_1(21654) <= 10849121;
srom_1(21655) <= 11392205;
srom_1(21656) <= 11921204;
srom_1(21657) <= 12433637;
srom_1(21658) <= 12927102;
srom_1(21659) <= 13399284;
srom_1(21660) <= 13847970;
srom_1(21661) <= 14271055;
srom_1(21662) <= 14666555;
srom_1(21663) <= 15032615;
srom_1(21664) <= 15367520;
srom_1(21665) <= 15669698;
srom_1(21666) <= 15937732;
srom_1(21667) <= 16170366;
srom_1(21668) <= 16366509;
srom_1(21669) <= 16525240;
srom_1(21670) <= 16645816;
srom_1(21671) <= 16727671;
srom_1(21672) <= 16770422;
srom_1(21673) <= 16773867;
srom_1(21674) <= 16737991;
srom_1(21675) <= 16662961;
srom_1(21676) <= 16549131;
srom_1(21677) <= 16397032;
srom_1(21678) <= 16207380;
srom_1(21679) <= 15981063;
srom_1(21680) <= 15719142;
srom_1(21681) <= 15422846;
srom_1(21682) <= 15093563;
srom_1(21683) <= 14732839;
srom_1(21684) <= 14342365;
srom_1(21685) <= 13923971;
srom_1(21686) <= 13479620;
srom_1(21687) <= 13011396;
srom_1(21688) <= 12521493;
srom_1(21689) <= 12012211;
srom_1(21690) <= 11485936;
srom_1(21691) <= 10945136;
srom_1(21692) <= 10392348;
srom_1(21693) <= 9830164;
srom_1(21694) <= 9261220;
srom_1(21695) <= 8688184;
srom_1(21696) <= 8113743;
srom_1(21697) <= 7540591;
srom_1(21698) <= 6971415;
srom_1(21699) <= 6408886;
srom_1(21700) <= 5855639;
srom_1(21701) <= 5314271;
srom_1(21702) <= 4787320;
srom_1(21703) <= 4277256;
srom_1(21704) <= 3786472;
srom_1(21705) <= 3317268;
srom_1(21706) <= 2871846;
srom_1(21707) <= 2452294;
srom_1(21708) <= 2060579;
srom_1(21709) <= 1698539;
srom_1(21710) <= 1367871;
srom_1(21711) <= 1070125;
srom_1(21712) <= 806698;
srom_1(21713) <= 578825;
srom_1(21714) <= 387575;
srom_1(21715) <= 233845;
srom_1(21716) <= 118355;
srom_1(21717) <= 41647;
srom_1(21718) <= 4081;
srom_1(21719) <= 5833;
srom_1(21720) <= 46895;
srom_1(21721) <= 127073;
srom_1(21722) <= 245993;
srom_1(21723) <= 403097;
srom_1(21724) <= 597647;
srom_1(21725) <= 828731;
srom_1(21726) <= 1095267;
srom_1(21727) <= 1396003;
srom_1(21728) <= 1729531;
srom_1(21729) <= 2094285;
srom_1(21730) <= 2488555;
srom_1(21731) <= 2910492;
srom_1(21732) <= 3358119;
srom_1(21733) <= 3829334;
srom_1(21734) <= 4321930;
srom_1(21735) <= 4833596;
srom_1(21736) <= 5361933;
srom_1(21737) <= 5904463;
srom_1(21738) <= 6458642;
srom_1(21739) <= 7021871;
srom_1(21740) <= 7591509;
srom_1(21741) <= 8164885;
srom_1(21742) <= 8739310;
srom_1(21743) <= 9312091;
srom_1(21744) <= 9880541;
srom_1(21745) <= 10441994;
srom_1(21746) <= 10993819;
srom_1(21747) <= 11533427;
srom_1(21748) <= 12058288;
srom_1(21749) <= 12565941;
srom_1(21750) <= 13054004;
srom_1(21751) <= 13520190;
srom_1(21752) <= 13962312;
srom_1(21753) <= 14378297;
srom_1(21754) <= 14766195;
srom_1(21755) <= 15124185;
srom_1(21756) <= 15450591;
srom_1(21757) <= 15743880;
srom_1(21758) <= 16002678;
srom_1(21759) <= 16225770;
srom_1(21760) <= 16412112;
srom_1(21761) <= 16560829;
srom_1(21762) <= 16671223;
srom_1(21763) <= 16742777;
srom_1(21764) <= 16775156;
srom_1(21765) <= 16768207;
srom_1(21766) <= 16721964;
srom_1(21767) <= 16636642;
srom_1(21768) <= 16512643;
srom_1(21769) <= 16350547;
srom_1(21770) <= 16151115;
srom_1(21771) <= 15915282;
srom_1(21772) <= 15644153;
srom_1(21773) <= 15339001;
srom_1(21774) <= 15001256;
srom_1(21775) <= 14632503;
srom_1(21776) <= 14234469;
srom_1(21777) <= 13809022;
srom_1(21778) <= 13358157;
srom_1(21779) <= 12883988;
srom_1(21780) <= 12388739;
srom_1(21781) <= 11874731;
srom_1(21782) <= 11344376;
srom_1(21783) <= 10800161;
srom_1(21784) <= 10244637;
srom_1(21785) <= 9680409;
srom_1(21786) <= 9110123;
srom_1(21787) <= 8536454;
srom_1(21788) <= 7962092;
srom_1(21789) <= 7389730;
srom_1(21790) <= 6822052;
srom_1(21791) <= 6261720;
srom_1(21792) <= 5711361;
srom_1(21793) <= 5173558;
srom_1(21794) <= 4650830;
srom_1(21795) <= 4145631;
srom_1(21796) <= 3660328;
srom_1(21797) <= 3197198;
srom_1(21798) <= 2758412;
srom_1(21799) <= 2346028;
srom_1(21800) <= 1961979;
srom_1(21801) <= 1608068;
srom_1(21802) <= 1285952;
srom_1(21803) <= 997144;
srom_1(21804) <= 742996;
srom_1(21805) <= 524702;
srom_1(21806) <= 343283;
srom_1(21807) <= 199593;
srom_1(21808) <= 94303;
srom_1(21809) <= 27908;
srom_1(21810) <= 720;
srom_1(21811) <= 12865;
srom_1(21812) <= 64286;
srom_1(21813) <= 154744;
srom_1(21814) <= 283812;
srom_1(21815) <= 450887;
srom_1(21816) <= 655185;
srom_1(21817) <= 895747;
srom_1(21818) <= 1171446;
srom_1(21819) <= 1480989;
srom_1(21820) <= 1822924;
srom_1(21821) <= 2195647;
srom_1(21822) <= 2597412;
srom_1(21823) <= 3026333;
srom_1(21824) <= 3480400;
srom_1(21825) <= 3957483;
srom_1(21826) <= 4455345;
srom_1(21827) <= 4971652;
srom_1(21828) <= 5503982;
srom_1(21829) <= 6049839;
srom_1(21830) <= 6606663;
srom_1(21831) <= 7171844;
srom_1(21832) <= 7742730;
srom_1(21833) <= 8316645;
srom_1(21834) <= 8890897;
srom_1(21835) <= 9462794;
srom_1(21836) <= 10029654;
srom_1(21837) <= 10588818;
srom_1(21838) <= 11137665;
srom_1(21839) <= 11673620;
srom_1(21840) <= 12194171;
srom_1(21841) <= 12696876;
srom_1(21842) <= 13179379;
srom_1(21843) <= 13639416;
srom_1(21844) <= 14074829;
srom_1(21845) <= 14483579;
srom_1(21846) <= 14863747;
srom_1(21847) <= 15213550;
srom_1(21848) <= 15531349;
srom_1(21849) <= 15815654;
srom_1(21850) <= 16065130;
srom_1(21851) <= 16278609;
srom_1(21852) <= 16455089;
srom_1(21853) <= 16593742;
srom_1(21854) <= 16693918;
srom_1(21855) <= 16755148;
srom_1(21856) <= 16777145;
srom_1(21857) <= 16759804;
srom_1(21858) <= 16703208;
srom_1(21859) <= 16607623;
srom_1(21860) <= 16473495;
srom_1(21861) <= 16301455;
srom_1(21862) <= 16092308;
srom_1(21863) <= 15847036;
srom_1(21864) <= 15566790;
srom_1(21865) <= 15252882;
srom_1(21866) <= 14906785;
srom_1(21867) <= 14530122;
srom_1(21868) <= 14124660;
srom_1(21869) <= 13692299;
srom_1(21870) <= 13235067;
srom_1(21871) <= 12755109;
srom_1(21872) <= 12254674;
srom_1(21873) <= 11736111;
srom_1(21874) <= 11201849;
srom_1(21875) <= 10654396;
srom_1(21876) <= 10096317;
srom_1(21877) <= 9530231;
srom_1(21878) <= 8958790;
srom_1(21879) <= 8384677;
srom_1(21880) <= 7810581;
srom_1(21881) <= 7239196;
srom_1(21882) <= 6673201;
srom_1(21883) <= 6115250;
srom_1(21884) <= 5567960;
srom_1(21885) <= 5033897;
srom_1(21886) <= 4515565;
srom_1(21887) <= 4015395;
srom_1(21888) <= 3535733;
srom_1(21889) <= 3078827;
srom_1(21890) <= 2646821;
srom_1(21891) <= 2241740;
srom_1(21892) <= 1865483;
srom_1(21893) <= 1519816;
srom_1(21894) <= 1206359;
srom_1(21895) <= 926582;
srom_1(21896) <= 681797;
srom_1(21897) <= 473152;
srom_1(21898) <= 301626;
srom_1(21899) <= 168021;
srom_1(21900) <= 72966;
srom_1(21901) <= 16906;
srom_1(21902) <= 104;
srom_1(21903) <= 22638;
srom_1(21904) <= 84403;
srom_1(21905) <= 185110;
srom_1(21906) <= 324285;
srom_1(21907) <= 501277;
srom_1(21908) <= 715255;
srom_1(21909) <= 965216;
srom_1(21910) <= 1249988;
srom_1(21911) <= 1568236;
srom_1(21912) <= 1918466;
srom_1(21913) <= 2299037;
srom_1(21914) <= 2708165;
srom_1(21915) <= 3143929;
srom_1(21916) <= 3604288;
srom_1(21917) <= 4087083;
srom_1(21918) <= 4590048;
srom_1(21919) <= 5110826;
srom_1(21920) <= 5646975;
srom_1(21921) <= 6195981;
srom_1(21922) <= 6755268;
srom_1(21923) <= 7322215;
srom_1(21924) <= 7894162;
srom_1(21925) <= 8468428;
srom_1(21926) <= 9042320;
srom_1(21927) <= 9613146;
srom_1(21928) <= 10178230;
srom_1(21929) <= 10734921;
srom_1(21930) <= 11280610;
srom_1(21931) <= 11812738;
srom_1(21932) <= 12328808;
srom_1(21933) <= 12826402;
srom_1(21934) <= 13303185;
srom_1(21935) <= 13756922;
srom_1(21936) <= 14185485;
srom_1(21937) <= 14586865;
srom_1(21938) <= 14959179;
srom_1(21939) <= 15300681;
srom_1(21940) <= 15609770;
srom_1(21941) <= 15884996;
srom_1(21942) <= 16125070;
srom_1(21943) <= 16328864;
srom_1(21944) <= 16495424;
srom_1(21945) <= 16623968;
srom_1(21946) <= 16713894;
srom_1(21947) <= 16764780;
srom_1(21948) <= 16776387;
srom_1(21949) <= 16748661;
srom_1(21950) <= 16681731;
srom_1(21951) <= 16575912;
srom_1(21952) <= 16431700;
srom_1(21953) <= 16249772;
srom_1(21954) <= 16030979;
srom_1(21955) <= 15776349;
srom_1(21956) <= 15487076;
srom_1(21957) <= 15164515;
srom_1(21958) <= 14810179;
srom_1(21959) <= 14425731;
srom_1(21960) <= 14012972;
srom_1(21961) <= 13573839;
srom_1(21962) <= 13110390;
srom_1(21963) <= 12624800;
srom_1(21964) <= 12119344;
srom_1(21965) <= 11596394;
srom_1(21966) <= 11058401;
srom_1(21967) <= 10507889;
srom_1(21968) <= 9947439;
srom_1(21969) <= 9379679;
srom_1(21970) <= 8807271;
srom_1(21971) <= 8232900;
srom_1(21972) <= 7659259;
srom_1(21973) <= 7089039;
srom_1(21974) <= 6524912;
srom_1(21975) <= 5969525;
srom_1(21976) <= 5425482;
srom_1(21977) <= 4895334;
srom_1(21978) <= 4381567;
srom_1(21979) <= 3886591;
srom_1(21980) <= 3412726;
srom_1(21981) <= 2962194;
srom_1(21982) <= 2537109;
srom_1(21983) <= 2139464;
srom_1(21984) <= 1771123;
srom_1(21985) <= 1433814;
srom_1(21986) <= 1129118;
srom_1(21987) <= 858464;
srom_1(21988) <= 623122;
srom_1(21989) <= 424195;
srom_1(21990) <= 262615;
srom_1(21991) <= 139142;
srom_1(21992) <= 54352;
srom_1(21993) <= 8645;
srom_1(21994) <= 2235;
srom_1(21995) <= 35151;
srom_1(21996) <= 107239;
srom_1(21997) <= 218162;
srom_1(21998) <= 367398;
srom_1(21999) <= 554249;
srom_1(22000) <= 777838;
srom_1(22001) <= 1037116;
srom_1(22002) <= 1330868;
srom_1(22003) <= 1657716;
srom_1(22004) <= 2016127;
srom_1(22005) <= 2404421;
srom_1(22006) <= 2820777;
srom_1(22007) <= 3263243;
srom_1(22008) <= 3729743;
srom_1(22009) <= 4218090;
srom_1(22010) <= 4725995;
srom_1(22011) <= 5251074;
srom_1(22012) <= 5790866;
srom_1(22013) <= 6342840;
srom_1(22014) <= 6904408;
srom_1(22015) <= 7472935;
srom_1(22016) <= 8045756;
srom_1(22017) <= 8620185;
srom_1(22018) <= 9193528;
srom_1(22019) <= 9763097;
srom_1(22020) <= 10326220;
srom_1(22021) <= 10880256;
srom_1(22022) <= 11422609;
srom_1(22023) <= 11950734;
srom_1(22024) <= 12462155;
srom_1(22025) <= 12954474;
srom_1(22026) <= 13425382;
srom_1(22027) <= 13872671;
srom_1(22028) <= 14294243;
srom_1(22029) <= 14688122;
srom_1(22030) <= 15052459;
srom_1(22031) <= 15385548;
srom_1(22032) <= 15685826;
srom_1(22033) <= 15951885;
srom_1(22034) <= 16182477;
srom_1(22035) <= 16376520;
srom_1(22036) <= 16533106;
srom_1(22037) <= 16651499;
srom_1(22038) <= 16731145;
srom_1(22039) <= 16771669;
srom_1(22040) <= 16772883;
srom_1(22041) <= 16734780;
srom_1(22042) <= 16657539;
srom_1(22043) <= 16541522;
srom_1(22044) <= 16387273;
srom_1(22045) <= 16195515;
srom_1(22046) <= 15967149;
srom_1(22047) <= 15703244;
srom_1(22048) <= 15405038;
srom_1(22049) <= 15073929;
srom_1(22050) <= 14711471;
srom_1(22051) <= 14319363;
srom_1(22052) <= 13899443;
srom_1(22053) <= 13453682;
srom_1(22054) <= 12984168;
srom_1(22055) <= 12493104;
srom_1(22056) <= 11982793;
srom_1(22057) <= 11455627;
srom_1(22058) <= 10914079;
srom_1(22059) <= 10360689;
srom_1(22060) <= 9798050;
srom_1(22061) <= 9228802;
srom_1(22062) <= 8655614;
srom_1(22063) <= 8081175;
srom_1(22064) <= 7508176;
srom_1(22065) <= 6939307;
srom_1(22066) <= 6377233;
srom_1(22067) <= 5824592;
srom_1(22068) <= 5283974;
srom_1(22069) <= 4757915;
srom_1(22070) <= 4248881;
srom_1(22071) <= 3759261;
srom_1(22072) <= 3291348;
srom_1(22073) <= 2847339;
srom_1(22074) <= 2429314;
srom_1(22075) <= 2039234;
srom_1(22076) <= 1678929;
srom_1(22077) <= 1350088;
srom_1(22078) <= 1054253;
srom_1(22079) <= 792811;
srom_1(22080) <= 566989;
srom_1(22081) <= 377845;
srom_1(22082) <= 226266;
srom_1(22083) <= 112963;
srom_1(22084) <= 38467;
srom_1(22085) <= 3128;
srom_1(22086) <= 7111;
srom_1(22087) <= 50398;
srom_1(22088) <= 132786;
srom_1(22089) <= 253888;
srom_1(22090) <= 413137;
srom_1(22091) <= 609786;
srom_1(22092) <= 842912;
srom_1(22093) <= 1111422;
srom_1(22094) <= 1414057;
srom_1(22095) <= 1749399;
srom_1(22096) <= 2115874;
srom_1(22097) <= 2511764;
srom_1(22098) <= 2935213;
srom_1(22099) <= 3384234;
srom_1(22100) <= 3856723;
srom_1(22101) <= 4350463;
srom_1(22102) <= 4863140;
srom_1(22103) <= 5392349;
srom_1(22104) <= 5935608;
srom_1(22105) <= 6490370;
srom_1(22106) <= 7054033;
srom_1(22107) <= 7623955;
srom_1(22108) <= 8197463;
srom_1(22109) <= 8771867;
srom_1(22110) <= 9344473;
srom_1(22111) <= 9912598;
srom_1(22112) <= 10473575;
srom_1(22113) <= 11024776;
srom_1(22114) <= 11563615;
srom_1(22115) <= 12087565;
srom_1(22116) <= 12594169;
srom_1(22117) <= 13081052;
srom_1(22118) <= 13545930;
srom_1(22119) <= 13986624;
srom_1(22120) <= 14401067;
srom_1(22121) <= 14787316;
srom_1(22122) <= 15143559;
srom_1(22123) <= 15468125;
srom_1(22124) <= 15759493;
srom_1(22125) <= 16016297;
srom_1(22126) <= 16237332;
srom_1(22127) <= 16421561;
srom_1(22128) <= 16568121;
srom_1(22129) <= 16676324;
srom_1(22130) <= 16745664;
srom_1(22131) <= 16775814;
srom_1(22132) <= 16766634;
srom_1(22133) <= 16718167;
srom_1(22134) <= 16630639;
srom_1(22135) <= 16504462;
srom_1(22136) <= 16340226;
srom_1(22137) <= 16138703;
srom_1(22138) <= 15900837;
srom_1(22139) <= 15627743;
srom_1(22140) <= 15320703;
srom_1(22141) <= 14981155;
srom_1(22142) <= 14610693;
srom_1(22143) <= 14211053;
srom_1(22144) <= 13784110;
srom_1(22145) <= 13331866;
srom_1(22146) <= 12856441;
srom_1(22147) <= 12360064;
srom_1(22148) <= 11845065;
srom_1(22149) <= 11313856;
srom_1(22150) <= 10768930;
srom_1(22151) <= 10212842;
srom_1(22152) <= 9648200;
srom_1(22153) <= 9077651;
srom_1(22154) <= 8503870;
srom_1(22155) <= 7929550;
srom_1(22156) <= 7357381;
srom_1(22157) <= 6790049;
srom_1(22158) <= 6230213;
srom_1(22159) <= 5680498;
srom_1(22160) <= 5143483;
srom_1(22161) <= 4621685;
srom_1(22162) <= 4117551;
srom_1(22163) <= 3633446;
srom_1(22164) <= 3171639;
srom_1(22165) <= 2734297;
srom_1(22166) <= 2323469;
srom_1(22167) <= 1941084;
srom_1(22168) <= 1588932;
srom_1(22169) <= 1268667;
srom_1(22170) <= 981790;
srom_1(22171) <= 729645;
srom_1(22172) <= 513416;
srom_1(22173) <= 334117;
srom_1(22174) <= 192588;
srom_1(22175) <= 89493;
srom_1(22176) <= 25315;
srom_1(22177) <= 356;
srom_1(22178) <= 14732;
srom_1(22179) <= 68376;
srom_1(22180) <= 161036;
srom_1(22181) <= 292279;
srom_1(22182) <= 461487;
srom_1(22183) <= 667869;
srom_1(22184) <= 910456;
srom_1(22185) <= 1188111;
srom_1(22186) <= 1499531;
srom_1(22187) <= 1843256;
srom_1(22188) <= 2217675;
srom_1(22189) <= 2621031;
srom_1(22190) <= 3051434;
srom_1(22191) <= 3506864;
srom_1(22192) <= 3985187;
srom_1(22193) <= 4484159;
srom_1(22194) <= 5001440;
srom_1(22195) <= 5534604;
srom_1(22196) <= 6081152;
srom_1(22197) <= 6638521;
srom_1(22198) <= 7204096;
srom_1(22199) <= 7775226;
srom_1(22200) <= 8349232;
srom_1(22201) <= 8923423;
srom_1(22202) <= 9495105;
srom_1(22203) <= 10061599;
srom_1(22204) <= 10620248;
srom_1(22205) <= 11168432;
srom_1(22206) <= 11703581;
srom_1(22207) <= 12223184;
srom_1(22208) <= 12724805;
srom_1(22209) <= 13206093;
srom_1(22210) <= 13664790;
srom_1(22211) <= 14098745;
srom_1(22212) <= 14505923;
srom_1(22213) <= 14884415;
srom_1(22214) <= 15232446;
srom_1(22215) <= 15548384;
srom_1(22216) <= 15830747;
srom_1(22217) <= 16078212;
srom_1(22218) <= 16289617;
srom_1(22219) <= 16463972;
srom_1(22220) <= 16600458;
srom_1(22221) <= 16698436;
srom_1(22222) <= 16757447;
srom_1(22223) <= 16777213;
srom_1(22224) <= 16757643;
srom_1(22225) <= 16698827;
srom_1(22226) <= 16601041;
srom_1(22227) <= 16464745;
srom_1(22228) <= 16290576;
srom_1(22229) <= 16079353;
srom_1(22230) <= 15832065;
srom_1(22231) <= 15549872;
srom_1(22232) <= 15234098;
srom_1(22233) <= 14886223;
srom_1(22234) <= 14507878;
srom_1(22235) <= 14100838;
srom_1(22236) <= 13667011;
srom_1(22237) <= 13208432;
srom_1(22238) <= 12727251;
srom_1(22239) <= 12225725;
srom_1(22240) <= 11706205;
srom_1(22241) <= 11171128;
srom_1(22242) <= 10623002;
srom_1(22243) <= 10064399;
srom_1(22244) <= 9497937;
srom_1(22245) <= 8926274;
srom_1(22246) <= 8352089;
srom_1(22247) <= 7778075;
srom_1(22248) <= 7206924;
srom_1(22249) <= 6641315;
srom_1(22250) <= 6083899;
srom_1(22251) <= 5537291;
srom_1(22252) <= 5004054;
srom_1(22253) <= 4486688;
srom_1(22254) <= 3987619;
srom_1(22255) <= 3509188;
srom_1(22256) <= 3053638;
srom_1(22257) <= 2623106;
srom_1(22258) <= 2219611;
srom_1(22259) <= 1845043;
srom_1(22260) <= 1501161;
srom_1(22261) <= 1189577;
srom_1(22262) <= 911751;
srom_1(22263) <= 668987;
srom_1(22264) <= 462422;
srom_1(22265) <= 293027;
srom_1(22266) <= 161594;
srom_1(22267) <= 68740;
srom_1(22268) <= 14902;
srom_1(22269) <= 330;
srom_1(22270) <= 25094;
srom_1(22271) <= 89077;
srom_1(22272) <= 191980;
srom_1(22273) <= 333319;
srom_1(22274) <= 512433;
srom_1(22275) <= 728480;
srom_1(22276) <= 980449;
srom_1(22277) <= 1267157;
srom_1(22278) <= 1587259;
srom_1(22279) <= 1939256;
srom_1(22280) <= 2321496;
srom_1(22281) <= 2732187;
srom_1(22282) <= 3169402;
srom_1(22283) <= 3631092;
srom_1(22284) <= 4115092;
srom_1(22285) <= 4619132;
srom_1(22286) <= 5140848;
srom_1(22287) <= 5677794;
srom_1(22288) <= 6227452;
srom_1(22289) <= 6787244;
srom_1(22290) <= 7354546;
srom_1(22291) <= 7926697;
srom_1(22292) <= 8501014;
srom_1(22293) <= 9074803;
srom_1(22294) <= 9645375;
srom_1(22295) <= 10210054;
srom_1(22296) <= 10766191;
srom_1(22297) <= 11311178;
srom_1(22298) <= 11842461;
srom_1(22299) <= 12357548;
srom_1(22300) <= 12854022;
srom_1(22301) <= 13329557;
srom_1(22302) <= 13781922;
srom_1(22303) <= 14208996;
srom_1(22304) <= 14608776;
srom_1(22305) <= 14979388;
srom_1(22306) <= 15319093;
srom_1(22307) <= 15626299;
srom_1(22308) <= 15899565;
srom_1(22309) <= 16137609;
srom_1(22310) <= 16339316;
srom_1(22311) <= 16503739;
srom_1(22312) <= 16630107;
srom_1(22313) <= 16717828;
srom_1(22314) <= 16766490;
srom_1(22315) <= 16775866;
srom_1(22316) <= 16745911;
srom_1(22317) <= 16676766;
srom_1(22318) <= 16568754;
srom_1(22319) <= 16422383;
srom_1(22320) <= 16238339;
srom_1(22321) <= 16017485;
srom_1(22322) <= 15760857;
srom_1(22323) <= 15469657;
srom_1(22324) <= 15145252;
srom_1(22325) <= 14789163;
srom_1(22326) <= 14403059;
srom_1(22327) <= 13988752;
srom_1(22328) <= 13548183;
srom_1(22329) <= 13083420;
srom_1(22330) <= 12596641;
srom_1(22331) <= 12090129;
srom_1(22332) <= 11566259;
srom_1(22333) <= 11027488;
srom_1(22334) <= 10476343;
srom_1(22335) <= 9915407;
srom_1(22336) <= 9347312;
srom_1(22337) <= 8774721;
srom_1(22338) <= 8200319;
srom_1(22339) <= 7626800;
srom_1(22340) <= 7056854;
srom_1(22341) <= 6493153;
srom_1(22342) <= 5938340;
srom_1(22343) <= 5395017;
srom_1(22344) <= 4865733;
srom_1(22345) <= 4352968;
srom_1(22346) <= 3859128;
srom_1(22347) <= 3386528;
srom_1(22348) <= 2937384;
srom_1(22349) <= 2513803;
srom_1(22350) <= 2117772;
srom_1(22351) <= 1751146;
srom_1(22352) <= 1415645;
srom_1(22353) <= 1112843;
srom_1(22354) <= 844160;
srom_1(22355) <= 610855;
srom_1(22356) <= 414023;
srom_1(22357) <= 254587;
srom_1(22358) <= 133293;
srom_1(22359) <= 50712;
srom_1(22360) <= 7229;
srom_1(22361) <= 3050;
srom_1(22362) <= 38194;
srom_1(22363) <= 112496;
srom_1(22364) <= 225607;
srom_1(22365) <= 376997;
srom_1(22366) <= 565957;
srom_1(22367) <= 791599;
srom_1(22368) <= 1052867;
srom_1(22369) <= 1348534;
srom_1(22370) <= 1677215;
srom_1(22371) <= 2037368;
srom_1(22372) <= 2427303;
srom_1(22373) <= 2845194;
srom_1(22374) <= 3289079;
srom_1(22375) <= 3756878;
srom_1(22376) <= 4246397;
srom_1(22377) <= 4755340;
srom_1(22378) <= 5281320;
srom_1(22379) <= 5821872;
srom_1(22380) <= 6374460;
srom_1(22381) <= 6936493;
srom_1(22382) <= 7505335;
srom_1(22383) <= 8078319;
srom_1(22384) <= 8652759;
srom_1(22385) <= 9225960;
srom_1(22386) <= 9795234;
srom_1(22387) <= 10357912;
srom_1(22388) <= 10911355;
srom_1(22389) <= 11452968;
srom_1(22390) <= 11980211;
srom_1(22391) <= 12490612;
srom_1(22392) <= 12981777;
srom_1(22393) <= 13451404;
srom_1(22394) <= 13897289;
srom_1(22395) <= 14317342;
srom_1(22396) <= 14709593;
srom_1(22397) <= 15072203;
srom_1(22398) <= 15403471;
srom_1(22399) <= 15701844;
srom_1(22400) <= 15965923;
srom_1(22401) <= 16194469;
srom_1(22402) <= 16386411;
srom_1(22403) <= 16540849;
srom_1(22404) <= 16657057;
srom_1(22405) <= 16734492;
srom_1(22406) <= 16772791;
srom_1(22407) <= 16771773;
srom_1(22408) <= 16731443;
srom_1(22409) <= 16651991;
srom_1(22410) <= 16533790;
srom_1(22411) <= 16377392;
srom_1(22412) <= 16183533;
srom_1(22413) <= 15953120;
srom_1(22414) <= 15687235;
srom_1(22415) <= 15387124;
srom_1(22416) <= 15054194;
srom_1(22417) <= 14690008;
srom_1(22418) <= 14296272;
srom_1(22419) <= 13874833;
srom_1(22420) <= 13427667;
srom_1(22421) <= 12956871;
srom_1(22422) <= 12464653;
srom_1(22423) <= 11953321;
srom_1(22424) <= 11425273;
srom_1(22425) <= 10882984;
srom_1(22426) <= 10328999;
srom_1(22427) <= 9765915;
srom_1(22428) <= 9196372;
srom_1(22429) <= 8623041;
srom_1(22430) <= 8048611;
srom_1(22431) <= 7475775;
srom_1(22432) <= 6907220;
srom_1(22433) <= 6345611;
srom_1(22434) <= 5793583;
srom_1(22435) <= 5253724;
srom_1(22436) <= 4728565;
srom_1(22437) <= 4220570;
srom_1(22438) <= 3732119;
srom_1(22439) <= 3265505;
srom_1(22440) <= 2822915;
srom_1(22441) <= 2406424;
srom_1(22442) <= 2017985;
srom_1(22443) <= 1659421;
srom_1(22444) <= 1332412;
srom_1(22445) <= 1038492;
srom_1(22446) <= 779039;
srom_1(22447) <= 555271;
srom_1(22448) <= 368235;
srom_1(22449) <= 218809;
srom_1(22450) <= 107695;
srom_1(22451) <= 35413;
srom_1(22452) <= 2301;
srom_1(22453) <= 8516;
srom_1(22454) <= 54028;
srom_1(22455) <= 138624;
srom_1(22456) <= 261907;
srom_1(22457) <= 423298;
srom_1(22458) <= 622042;
srom_1(22459) <= 857206;
srom_1(22460) <= 1127687;
srom_1(22461) <= 1432217;
srom_1(22462) <= 1769368;
srom_1(22463) <= 2137558;
srom_1(22464) <= 2535063;
srom_1(22465) <= 2960016;
srom_1(22466) <= 3410426;
srom_1(22467) <= 3884180;
srom_1(22468) <= 4379057;
srom_1(22469) <= 4892737;
srom_1(22470) <= 5422809;
srom_1(22471) <= 5966790;
srom_1(22472) <= 6522127;
srom_1(22473) <= 7086216;
srom_1(22474) <= 7656413;
srom_1(22475) <= 8230043;
srom_1(22476) <= 8804417;
srom_1(22477) <= 9376842;
srom_1(22478) <= 9944631;
srom_1(22479) <= 10505125;
srom_1(22480) <= 11055693;
srom_1(22481) <= 11593754;
srom_1(22482) <= 12116785;
srom_1(22483) <= 12622334;
srom_1(22484) <= 13108029;
srom_1(22485) <= 13571593;
srom_1(22486) <= 14010852;
srom_1(22487) <= 14423747;
srom_1(22488) <= 14808341;
srom_1(22489) <= 15162830;
srom_1(22490) <= 15485553;
srom_1(22491) <= 15774996;
srom_1(22492) <= 16029801;
srom_1(22493) <= 16248774;
srom_1(22494) <= 16430888;
srom_1(22495) <= 16575290;
srom_1(22496) <= 16681301;
srom_1(22497) <= 16748425;
srom_1(22498) <= 16776346;
srom_1(22499) <= 16764935;
srom_1(22500) <= 16714244;
srom_1(22501) <= 16624512;
srom_1(22502) <= 16496158;
srom_1(22503) <= 16329785;
srom_1(22504) <= 16126174;
srom_1(22505) <= 15886278;
srom_1(22506) <= 15611223;
srom_1(22507) <= 15302299;
srom_1(22508) <= 14960954;
srom_1(22509) <= 14588790;
srom_1(22510) <= 14187550;
srom_1(22511) <= 13759117;
srom_1(22512) <= 13305500;
srom_1(22513) <= 12828826;
srom_1(22514) <= 12331330;
srom_1(22515) <= 11815346;
srom_1(22516) <= 11283292;
srom_1(22517) <= 10737664;
srom_1(22518) <= 10181021;
srom_1(22519) <= 9615972;
srom_1(22520) <= 9045168;
srom_1(22521) <= 8471285;
srom_1(22522) <= 7897014;
srom_1(22523) <= 7325049;
srom_1(22524) <= 6758071;
srom_1(22525) <= 6198739;
srom_1(22526) <= 5649676;
srom_1(22527) <= 5113457;
srom_1(22528) <= 4592596;
srom_1(22529) <= 4089536;
srom_1(22530) <= 3606636;
srom_1(22531) <= 3146160;
srom_1(22532) <= 2710267;
srom_1(22533) <= 2301003;
srom_1(22534) <= 1920285;
srom_1(22535) <= 1569899;
srom_1(22536) <= 1251489;
srom_1(22537) <= 966547;
srom_1(22538) <= 716410;
srom_1(22539) <= 502250;
srom_1(22540) <= 325072;
srom_1(22541) <= 185707;
srom_1(22542) <= 84808;
srom_1(22543) <= 22849;
srom_1(22544) <= 119;
srom_1(22545) <= 16726;
srom_1(22546) <= 72591;
srom_1(22547) <= 167453;
srom_1(22548) <= 300867;
srom_1(22549) <= 472207;
srom_1(22550) <= 680670;
srom_1(22551) <= 925278;
srom_1(22552) <= 1204884;
srom_1(22553) <= 1518177;
srom_1(22554) <= 1863687;
srom_1(22555) <= 2239796;
srom_1(22556) <= 2644738;
srom_1(22557) <= 3076615;
srom_1(22558) <= 3533402;
srom_1(22559) <= 4012957;
srom_1(22560) <= 4513031;
srom_1(22561) <= 5031278;
srom_1(22562) <= 5565269;
srom_1(22563) <= 6112500;
srom_1(22564) <= 6670405;
srom_1(22565) <= 7236366;
srom_1(22566) <= 7807731;
srom_1(22567) <= 8381819;
srom_1(22568) <= 8955940;
srom_1(22569) <= 9527400;
srom_1(22570) <= 10093520;
srom_1(22571) <= 10651645;
srom_1(22572) <= 11199158;
srom_1(22573) <= 11733491;
srom_1(22574) <= 12252139;
srom_1(22575) <= 12752669;
srom_1(22576) <= 13232735;
srom_1(22577) <= 13690085;
srom_1(22578) <= 14122574;
srom_1(22579) <= 14528176;
srom_1(22580) <= 14904986;
srom_1(22581) <= 15251239;
srom_1(22582) <= 15565311;
srom_1(22583) <= 15845728;
srom_1(22584) <= 16091177;
srom_1(22585) <= 16300506;
srom_1(22586) <= 16472733;
srom_1(22587) <= 16607051;
srom_1(22588) <= 16702829;
srom_1(22589) <= 16759620;
srom_1(22590) <= 16777156;
srom_1(22591) <= 16755355;
srom_1(22592) <= 16694319;
srom_1(22593) <= 16594336;
srom_1(22594) <= 16455872;
srom_1(22595) <= 16279579;
srom_1(22596) <= 16066282;
srom_1(22597) <= 15816982;
srom_1(22598) <= 15532847;
srom_1(22599) <= 15215211;
srom_1(22600) <= 14865563;
srom_1(22601) <= 14485541;
srom_1(22602) <= 14076930;
srom_1(22603) <= 13641643;
srom_1(22604) <= 13181724;
srom_1(22605) <= 12699328;
srom_1(22606) <= 12196717;
srom_1(22607) <= 11676249;
srom_1(22608) <= 11140364;
srom_1(22609) <= 10591575;
srom_1(22610) <= 10032455;
srom_1(22611) <= 9465627;
srom_1(22612) <= 8893749;
srom_1(22613) <= 8319502;
srom_1(22614) <= 7745578;
srom_1(22615) <= 7174670;
srom_1(22616) <= 6609455;
srom_1(22617) <= 6052583;
srom_1(22618) <= 5506665;
srom_1(22619) <= 4974262;
srom_1(22620) <= 4457869;
srom_1(22621) <= 3959909;
srom_1(22622) <= 3482717;
srom_1(22623) <= 3028531;
srom_1(22624) <= 2599479;
srom_1(22625) <= 2197575;
srom_1(22626) <= 1824702;
srom_1(22627) <= 1482610;
srom_1(22628) <= 1172903;
srom_1(22629) <= 897032;
srom_1(22630) <= 656292;
srom_1(22631) <= 451812;
srom_1(22632) <= 284550;
srom_1(22633) <= 155290;
srom_1(22634) <= 64640;
srom_1(22635) <= 13023;
srom_1(22636) <= 683;
srom_1(22637) <= 27676;
srom_1(22638) <= 93876;
srom_1(22639) <= 198974;
srom_1(22640) <= 342475;
srom_1(22641) <= 523707;
srom_1(22642) <= 741821;
srom_1(22643) <= 995793;
srom_1(22644) <= 1284433;
srom_1(22645) <= 1606386;
srom_1(22646) <= 1960143;
srom_1(22647) <= 2344046;
srom_1(22648) <= 2756294;
srom_1(22649) <= 3194954;
srom_1(22650) <= 3657968;
srom_1(22651) <= 4143166;
srom_1(22652) <= 4648273;
srom_1(22653) <= 5170919;
srom_1(22654) <= 5708654;
srom_1(22655) <= 6258956;
srom_1(22656) <= 6819245;
srom_1(22657) <= 7386893;
srom_1(22658) <= 7959239;
srom_1(22659) <= 8533598;
srom_1(22660) <= 9107277;
srom_1(22661) <= 9677586;
srom_1(22662) <= 10241850;
srom_1(22663) <= 10797424;
srom_1(22664) <= 11341702;
srom_1(22665) <= 11872133;
srom_1(22666) <= 12386227;
srom_1(22667) <= 12881576;
srom_1(22668) <= 13355855;
srom_1(22669) <= 13806841;
srom_1(22670) <= 14232420;
srom_1(22671) <= 14630594;
srom_1(22672) <= 14999498;
srom_1(22673) <= 15337401;
srom_1(22674) <= 15642719;
srom_1(22675) <= 15914020;
srom_1(22676) <= 16150031;
srom_1(22677) <= 16349647;
srom_1(22678) <= 16511930;
srom_1(22679) <= 16636121;
srom_1(22680) <= 16721636;
srom_1(22681) <= 16768074;
srom_1(22682) <= 16775219;
srom_1(22683) <= 16743035;
srom_1(22684) <= 16671675;
srom_1(22685) <= 16561473;
srom_1(22686) <= 16412945;
srom_1(22687) <= 16226789;
srom_1(22688) <= 16003876;
srom_1(22689) <= 15745253;
srom_1(22690) <= 15452132;
srom_1(22691) <= 15125888;
srom_1(22692) <= 14768050;
srom_1(22693) <= 14380297;
srom_1(22694) <= 13964447;
srom_1(22695) <= 13522450;
srom_1(22696) <= 13056378;
srom_1(22697) <= 12568418;
srom_1(22698) <= 12060857;
srom_1(22699) <= 11536076;
srom_1(22700) <= 10996535;
srom_1(22701) <= 10444764;
srom_1(22702) <= 9883352;
srom_1(22703) <= 9314930;
srom_1(22704) <= 8742165;
srom_1(22705) <= 8167741;
srom_1(22706) <= 7594353;
srom_1(22707) <= 7024690;
srom_1(22708) <= 6461422;
srom_1(22709) <= 5907192;
srom_1(22710) <= 5364598;
srom_1(22711) <= 4836184;
srom_1(22712) <= 4324430;
srom_1(22713) <= 3831733;
srom_1(22714) <= 3360405;
srom_1(22715) <= 2912656;
srom_1(22716) <= 2490586;
srom_1(22717) <= 2096174;
srom_1(22718) <= 1731269;
srom_1(22719) <= 1397582;
srom_1(22720) <= 1096679;
srom_1(22721) <= 829970;
srom_1(22722) <= 598706;
srom_1(22723) <= 403972;
srom_1(22724) <= 246680;
srom_1(22725) <= 127569;
srom_1(22726) <= 47197;
srom_1(22727) <= 5940;
srom_1(22728) <= 3993;
srom_1(22729) <= 41363;
srom_1(22730) <= 117877;
srom_1(22731) <= 233175;
srom_1(22732) <= 386717;
srom_1(22733) <= 577783;
srom_1(22734) <= 805476;
srom_1(22735) <= 1068729;
srom_1(22736) <= 1366307;
srom_1(22737) <= 1696816;
srom_1(22738) <= 2058704;
srom_1(22739) <= 2450276;
srom_1(22740) <= 2869694;
srom_1(22741) <= 3314993;
srom_1(22742) <= 3784083;
srom_1(22743) <= 4274766;
srom_1(22744) <= 4784740;
srom_1(22745) <= 5311613;
srom_1(22746) <= 5852916;
srom_1(22747) <= 6406109;
srom_1(22748) <= 6968599;
srom_1(22749) <= 7537748;
srom_1(22750) <= 8110887;
srom_1(22751) <= 8685328;
srom_1(22752) <= 9258378;
srom_1(22753) <= 9827349;
srom_1(22754) <= 10389574;
srom_1(22755) <= 10942415;
srom_1(22756) <= 11483280;
srom_1(22757) <= 12009634;
srom_1(22758) <= 12519007;
srom_1(22759) <= 13009011;
srom_1(22760) <= 13477349;
srom_1(22761) <= 13921824;
srom_1(22762) <= 14340352;
srom_1(22763) <= 14730969;
srom_1(22764) <= 15091846;
srom_1(22765) <= 15421288;
srom_1(22766) <= 15717752;
srom_1(22767) <= 15979847;
srom_1(22768) <= 16206345;
srom_1(22769) <= 16396182;
srom_1(22770) <= 16548468;
srom_1(22771) <= 16662491;
srom_1(22772) <= 16737714;
srom_1(22773) <= 16773786;
srom_1(22774) <= 16770536;
srom_1(22775) <= 16727981;
srom_1(22776) <= 16646319;
srom_1(22777) <= 16525935;
srom_1(22778) <= 16367391;
srom_1(22779) <= 16171432;
srom_1(22780) <= 15938977;
srom_1(22781) <= 15671116;
srom_1(22782) <= 15369105;
srom_1(22783) <= 15034359;
srom_1(22784) <= 14668449;
srom_1(22785) <= 14273091;
srom_1(22786) <= 13850139;
srom_1(22787) <= 13401576;
srom_1(22788) <= 12929505;
srom_1(22789) <= 12436140;
srom_1(22790) <= 11923795;
srom_1(22791) <= 11394872;
srom_1(22792) <= 10851852;
srom_1(22793) <= 10297281;
srom_1(22794) <= 9733759;
srom_1(22795) <= 9163930;
srom_1(22796) <= 8590464;
srom_1(22797) <= 8016053;
srom_1(22798) <= 7443388;
srom_1(22799) <= 6875155;
srom_1(22800) <= 6314020;
srom_1(22801) <= 5762613;
srom_1(22802) <= 5223521;
srom_1(22803) <= 4699270;
srom_1(22804) <= 4192321;
srom_1(22805) <= 3705048;
srom_1(22806) <= 3239739;
srom_1(22807) <= 2798575;
srom_1(22808) <= 2383624;
srom_1(22809) <= 1996833;
srom_1(22810) <= 1640014;
srom_1(22811) <= 1314843;
srom_1(22812) <= 1022842;
srom_1(22813) <= 765382;
srom_1(22814) <= 543670;
srom_1(22815) <= 358746;
srom_1(22816) <= 211477;
srom_1(22817) <= 102553;
srom_1(22818) <= 32485;
srom_1(22819) <= 1601;
srom_1(22820) <= 10048;
srom_1(22821) <= 57784;
srom_1(22822) <= 144586;
srom_1(22823) <= 270047;
srom_1(22824) <= 433579;
srom_1(22825) <= 634415;
srom_1(22826) <= 871613;
srom_1(22827) <= 1144061;
srom_1(22828) <= 1450481;
srom_1(22829) <= 1789436;
srom_1(22830) <= 2159337;
srom_1(22831) <= 2558449;
srom_1(22832) <= 2984901;
srom_1(22833) <= 3436693;
srom_1(22834) <= 3911705;
srom_1(22835) <= 4407712;
srom_1(22836) <= 4922386;
srom_1(22837) <= 5453315;
srom_1(22838) <= 5998008;
srom_1(22839) <= 6553911;
srom_1(22840) <= 7118419;
srom_1(22841) <= 7688882;
srom_1(22842) <= 8262627;
srom_1(22843) <= 8836962;
srom_1(22844) <= 9409195;
srom_1(22845) <= 9976642;
srom_1(22846) <= 10536642;
srom_1(22847) <= 11086569;
srom_1(22848) <= 11623845;
srom_1(22849) <= 12145950;
srom_1(22850) <= 12650435;
srom_1(22851) <= 13134934;
srom_1(22852) <= 13597177;
srom_1(22853) <= 14034995;
srom_1(22854) <= 14446335;
srom_1(22855) <= 14829268;
srom_1(22856) <= 15181999;
srom_1(22857) <= 15502873;
srom_1(22858) <= 15790386;
srom_1(22859) <= 16043190;
srom_1(22860) <= 16260098;
srom_1(22861) <= 16440095;
srom_1(22862) <= 16582335;
srom_1(22863) <= 16686152;
srom_1(22864) <= 16751059;
srom_1(22865) <= 16776752;
srom_1(22866) <= 16763109;
srom_1(22867) <= 16710196;
srom_1(22868) <= 16618260;
srom_1(22869) <= 16487732;
srom_1(22870) <= 16319225;
srom_1(22871) <= 16113528;
srom_1(22872) <= 15871607;
srom_1(22873) <= 15594595;
srom_1(22874) <= 15283792;
srom_1(22875) <= 14940654;
srom_1(22876) <= 14566793;
srom_1(22877) <= 14163959;
srom_1(22878) <= 13734043;
srom_1(22879) <= 13279060;
srom_1(22880) <= 12801144;
srom_1(22881) <= 12302537;
srom_1(22882) <= 11785575;
srom_1(22883) <= 11252684;
srom_1(22884) <= 10706363;
srom_1(22885) <= 10149172;
srom_1(22886) <= 9583726;
srom_1(22887) <= 9012675;
srom_1(22888) <= 8438698;
srom_1(22889) <= 7864486;
srom_1(22890) <= 7292732;
srom_1(22891) <= 6726117;
srom_1(22892) <= 6167297;
srom_1(22893) <= 5618895;
srom_1(22894) <= 5083480;
srom_1(22895) <= 4563564;
srom_1(22896) <= 4061585;
srom_1(22897) <= 3579897;
srom_1(22898) <= 3120759;
srom_1(22899) <= 2686323;
srom_1(22900) <= 2278628;
srom_1(22901) <= 1899584;
srom_1(22902) <= 1550970;
srom_1(22903) <= 1234419;
srom_1(22904) <= 951417;
srom_1(22905) <= 703291;
srom_1(22906) <= 491203;
srom_1(22907) <= 316149;
srom_1(22908) <= 178950;
srom_1(22909) <= 80249;
srom_1(22910) <= 20508;
srom_1(22911) <= 8;
srom_1(22912) <= 18846;
srom_1(22913) <= 76932;
srom_1(22914) <= 173994;
srom_1(22915) <= 309577;
srom_1(22916) <= 483046;
srom_1(22917) <= 693587;
srom_1(22918) <= 940212;
srom_1(22919) <= 1221765;
srom_1(22920) <= 1536926;
srom_1(22921) <= 1884217;
srom_1(22922) <= 2262010;
srom_1(22923) <= 2668532;
srom_1(22924) <= 3101877;
srom_1(22925) <= 3560014;
srom_1(22926) <= 4040793;
srom_1(22927) <= 4541961;
srom_1(22928) <= 5061168;
srom_1(22929) <= 5595977;
srom_1(22930) <= 6143883;
srom_1(22931) <= 6702314;
srom_1(22932) <= 7268654;
srom_1(22933) <= 7840245;
srom_1(22934) <= 8414407;
srom_1(22935) <= 8988449;
srom_1(22936) <= 9559677;
srom_1(22937) <= 10125415;
srom_1(22938) <= 10683007;
srom_1(22939) <= 11229841;
srom_1(22940) <= 11763351;
srom_1(22941) <= 12281035;
srom_1(22942) <= 12780467;
srom_1(22943) <= 13259303;
srom_1(22944) <= 13715300;
srom_1(22945) <= 14146317;
srom_1(22946) <= 14550335;
srom_1(22947) <= 14925458;
srom_1(22948) <= 15269928;
srom_1(22949) <= 15582129;
srom_1(22950) <= 15860597;
srom_1(22951) <= 16104026;
srom_1(22952) <= 16311275;
srom_1(22953) <= 16481372;
srom_1(22954) <= 16613519;
srom_1(22955) <= 16707097;
srom_1(22956) <= 16761666;
srom_1(22957) <= 16776971;
srom_1(22958) <= 16752941;
srom_1(22959) <= 16689687;
srom_1(22960) <= 16587506;
srom_1(22961) <= 16446878;
srom_1(22962) <= 16268462;
srom_1(22963) <= 16053095;
srom_1(22964) <= 15801786;
srom_1(22965) <= 15515714;
srom_1(22966) <= 15196221;
srom_1(22967) <= 14844805;
srom_1(22968) <= 14463113;
srom_1(22969) <= 14052936;
srom_1(22970) <= 13616197;
srom_1(22971) <= 13154943;
srom_1(22972) <= 12671339;
srom_1(22973) <= 12167652;
srom_1(22974) <= 11646243;
srom_1(22975) <= 11109559;
srom_1(22976) <= 10560114;
srom_1(22977) <= 10000487;
srom_1(22978) <= 9433301;
srom_1(22979) <= 8861217;
srom_1(22980) <= 8286916;
srom_1(22981) <= 7713091;
srom_1(22982) <= 7142435;
srom_1(22983) <= 6577622;
srom_1(22984) <= 6021302;
srom_1(22985) <= 5476083;
srom_1(22986) <= 4944521;
srom_1(22987) <= 4429110;
srom_1(22988) <= 3932267;
srom_1(22989) <= 3456320;
srom_1(22990) <= 3003503;
srom_1(22991) <= 2575939;
srom_1(22992) <= 2175632;
srom_1(22993) <= 1804460;
srom_1(22994) <= 1464163;
srom_1(22995) <= 1156338;
srom_1(22996) <= 882427;
srom_1(22997) <= 643715;
srom_1(22998) <= 441321;
srom_1(22999) <= 276195;
srom_1(23000) <= 149111;
srom_1(23001) <= 60665;
srom_1(23002) <= 11271;
srom_1(23003) <= 1162;
srom_1(23004) <= 30384;
srom_1(23005) <= 98801;
srom_1(23006) <= 206091;
srom_1(23007) <= 351752;
srom_1(23008) <= 535101;
srom_1(23009) <= 755277;
srom_1(23010) <= 1011249;
srom_1(23011) <= 1301816;
srom_1(23012) <= 1625615;
srom_1(23013) <= 1981128;
srom_1(23014) <= 2366688;
srom_1(23015) <= 2780487;
srom_1(23016) <= 3220584;
srom_1(23017) <= 3684916;
srom_1(23018) <= 4171305;
srom_1(23019) <= 4677470;
srom_1(23020) <= 5201038;
srom_1(23021) <= 5739554;
srom_1(23022) <= 6290492;
srom_1(23023) <= 6851269;
srom_1(23024) <= 7419255;
srom_1(23025) <= 7991787;
srom_1(23026) <= 8566179;
srom_1(23027) <= 9139739;
srom_1(23028) <= 9709777;
srom_1(23029) <= 10273619;
srom_1(23030) <= 10828621;
srom_1(23031) <= 11372182;
srom_1(23032) <= 11901751;
srom_1(23033) <= 12414846;
srom_1(23034) <= 12909061;
srom_1(23035) <= 13382078;
srom_1(23036) <= 13831679;
srom_1(23037) <= 14255755;
srom_1(23038) <= 14652318;
srom_1(23039) <= 15019508;
srom_1(23040) <= 15355604;
srom_1(23041) <= 15659029;
srom_1(23042) <= 15928361;
srom_1(23043) <= 16162336;
srom_1(23044) <= 16359858;
srom_1(23045) <= 16520000;
srom_1(23046) <= 16642010;
srom_1(23047) <= 16725318;
srom_1(23048) <= 16769532;
srom_1(23049) <= 16774445;
srom_1(23050) <= 16740034;
srom_1(23051) <= 16666460;
srom_1(23052) <= 16554068;
srom_1(23053) <= 16403386;
srom_1(23054) <= 16215120;
srom_1(23055) <= 15990152;
srom_1(23056) <= 15729538;
srom_1(23057) <= 15434500;
srom_1(23058) <= 15106422;
srom_1(23059) <= 14746841;
srom_1(23060) <= 14357445;
srom_1(23061) <= 13940058;
srom_1(23062) <= 13496639;
srom_1(23063) <= 13029266;
srom_1(23064) <= 12540132;
srom_1(23065) <= 12031530;
srom_1(23066) <= 11505845;
srom_1(23067) <= 10965542;
srom_1(23068) <= 10413155;
srom_1(23069) <= 9851274;
srom_1(23070) <= 9282535;
srom_1(23071) <= 8709603;
srom_1(23072) <= 8135166;
srom_1(23073) <= 7561918;
srom_1(23074) <= 6992546;
srom_1(23075) <= 6429721;
srom_1(23076) <= 5876081;
srom_1(23077) <= 5334224;
srom_1(23078) <= 4806690;
srom_1(23079) <= 4295953;
srom_1(23080) <= 3804407;
srom_1(23081) <= 3334358;
srom_1(23082) <= 2888011;
srom_1(23083) <= 2467458;
srom_1(23084) <= 2074671;
srom_1(23085) <= 1711492;
srom_1(23086) <= 1379624;
srom_1(23087) <= 1080624;
srom_1(23088) <= 815894;
srom_1(23089) <= 586675;
srom_1(23090) <= 394041;
srom_1(23091) <= 238897;
srom_1(23092) <= 121970;
srom_1(23093) <= 43808;
srom_1(23094) <= 4777;
srom_1(23095) <= 5061;
srom_1(23096) <= 44659;
srom_1(23097) <= 123384;
srom_1(23098) <= 240867;
srom_1(23099) <= 396558;
srom_1(23100) <= 589727;
srom_1(23101) <= 819467;
srom_1(23102) <= 1084701;
srom_1(23103) <= 1384186;
srom_1(23104) <= 1716517;
srom_1(23105) <= 2080136;
srom_1(23106) <= 2473337;
srom_1(23107) <= 2894278;
srom_1(23108) <= 3340983;
srom_1(23109) <= 3811358;
srom_1(23110) <= 4303197;
srom_1(23111) <= 4814194;
srom_1(23112) <= 5341953;
srom_1(23113) <= 5883998;
srom_1(23114) <= 6437789;
srom_1(23115) <= 7000728;
srom_1(23116) <= 7570174;
srom_1(23117) <= 8143459;
srom_1(23118) <= 8717894;
srom_1(23119) <= 9290784;
srom_1(23120) <= 9859443;
srom_1(23121) <= 10421206;
srom_1(23122) <= 10973436;
srom_1(23123) <= 11513546;
srom_1(23124) <= 12039002;
srom_1(23125) <= 12547340;
srom_1(23126) <= 13036176;
srom_1(23127) <= 13503218;
srom_1(23128) <= 13946275;
srom_1(23129) <= 14363271;
srom_1(23130) <= 14752250;
srom_1(23131) <= 15111387;
srom_1(23132) <= 15438999;
srom_1(23133) <= 15733550;
srom_1(23134) <= 15993657;
srom_1(23135) <= 16218102;
srom_1(23136) <= 16405831;
srom_1(23137) <= 16555965;
srom_1(23138) <= 16667799;
srom_1(23139) <= 16740810;
srom_1(23140) <= 16774654;
srom_1(23141) <= 16769173;
srom_1(23142) <= 16724392;
srom_1(23143) <= 16640523;
srom_1(23144) <= 16517957;
srom_1(23145) <= 16357270;
srom_1(23146) <= 16159215;
srom_1(23147) <= 15924721;
srom_1(23148) <= 15654887;
srom_1(23149) <= 15350980;
srom_1(23150) <= 15014423;
srom_1(23151) <= 14646796;
srom_1(23152) <= 14249822;
srom_1(23153) <= 13825363;
srom_1(23154) <= 13375409;
srom_1(23155) <= 12902070;
srom_1(23156) <= 12407566;
srom_1(23157) <= 11894216;
srom_1(23158) <= 11364426;
srom_1(23159) <= 10820682;
srom_1(23160) <= 10265533;
srom_1(23161) <= 9701583;
srom_1(23162) <= 9131476;
srom_1(23163) <= 8557885;
srom_1(23164) <= 7983500;
srom_1(23165) <= 7411015;
srom_1(23166) <= 6843114;
srom_1(23167) <= 6282460;
srom_1(23168) <= 5731683;
srom_1(23169) <= 5193366;
srom_1(23170) <= 4670031;
srom_1(23171) <= 4164135;
srom_1(23172) <= 3678048;
srom_1(23173) <= 3214051;
srom_1(23174) <= 2774319;
srom_1(23175) <= 2360915;
srom_1(23176) <= 1975776;
srom_1(23177) <= 1620709;
srom_1(23178) <= 1297380;
srom_1(23179) <= 1007303;
srom_1(23180) <= 751840;
srom_1(23181) <= 532189;
srom_1(23182) <= 349379;
srom_1(23183) <= 204267;
srom_1(23184) <= 97535;
srom_1(23185) <= 29682;
srom_1(23186) <= 1028;
srom_1(23187) <= 11705;
srom_1(23188) <= 61665;
srom_1(23189) <= 150673;
srom_1(23190) <= 278311;
srom_1(23191) <= 443981;
srom_1(23192) <= 646906;
srom_1(23193) <= 886135;
srom_1(23194) <= 1160545;
srom_1(23195) <= 1468850;
srom_1(23196) <= 1809604;
srom_1(23197) <= 2181210;
srom_1(23198) <= 2581924;
srom_1(23199) <= 3009867;
srom_1(23200) <= 3463034;
srom_1(23201) <= 3939298;
srom_1(23202) <= 4436426;
srom_1(23203) <= 4952088;
srom_1(23204) <= 5483865;
srom_1(23205) <= 6029262;
srom_1(23206) <= 6585724;
srom_1(23207) <= 7150640;
srom_1(23208) <= 7721361;
srom_1(23209) <= 8295212;
srom_1(23210) <= 8869500;
srom_1(23211) <= 9441533;
srom_1(23212) <= 10008628;
srom_1(23213) <= 10568127;
srom_1(23214) <= 11117405;
srom_1(23215) <= 11653887;
srom_1(23216) <= 12175057;
srom_1(23217) <= 12678471;
srom_1(23218) <= 13161768;
srom_1(23219) <= 13622683;
srom_1(23220) <= 14059053;
srom_1(23221) <= 14468832;
srom_1(23222) <= 14850099;
srom_1(23223) <= 15201066;
srom_1(23224) <= 15520086;
srom_1(23225) <= 15805665;
srom_1(23226) <= 16056463;
srom_1(23227) <= 16271304;
srom_1(23228) <= 16449180;
srom_1(23229) <= 16589257;
srom_1(23230) <= 16690878;
srom_1(23231) <= 16753567;
srom_1(23232) <= 16777030;
srom_1(23233) <= 16761157;
srom_1(23234) <= 16706022;
srom_1(23235) <= 16611884;
srom_1(23236) <= 16479184;
srom_1(23237) <= 16308545;
srom_1(23238) <= 16100766;
srom_1(23239) <= 15856822;
srom_1(23240) <= 15577857;
srom_1(23241) <= 15265180;
srom_1(23242) <= 14920256;
srom_1(23243) <= 14544702;
srom_1(23244) <= 14140281;
srom_1(23245) <= 13708888;
srom_1(23246) <= 13252546;
srom_1(23247) <= 12773396;
srom_1(23248) <= 12273684;
srom_1(23249) <= 11755753;
srom_1(23250) <= 11222033;
srom_1(23251) <= 10675026;
srom_1(23252) <= 10117297;
srom_1(23253) <= 9551462;
srom_1(23254) <= 8980173;
srom_1(23255) <= 8406111;
srom_1(23256) <= 7831966;
srom_1(23257) <= 7260432;
srom_1(23258) <= 6694188;
srom_1(23259) <= 6135890;
srom_1(23260) <= 5588155;
srom_1(23261) <= 5053553;
srom_1(23262) <= 4534590;
srom_1(23263) <= 4033700;
srom_1(23264) <= 3553232;
srom_1(23265) <= 3095438;
srom_1(23266) <= 2662466;
srom_1(23267) <= 2256345;
srom_1(23268) <= 1878981;
srom_1(23269) <= 1532143;
srom_1(23270) <= 1217457;
srom_1(23271) <= 936399;
srom_1(23272) <= 690287;
srom_1(23273) <= 480275;
srom_1(23274) <= 307348;
srom_1(23275) <= 172317;
srom_1(23276) <= 75815;
srom_1(23277) <= 18294;
srom_1(23278) <= 24;
srom_1(23279) <= 21092;
srom_1(23280) <= 81398;
srom_1(23281) <= 180659;
srom_1(23282) <= 318409;
srom_1(23283) <= 494004;
srom_1(23284) <= 706620;
srom_1(23285) <= 955258;
srom_1(23286) <= 1238755;
srom_1(23287) <= 1555779;
srom_1(23288) <= 1904845;
srom_1(23289) <= 2284316;
srom_1(23290) <= 2692411;
srom_1(23291) <= 3127218;
srom_1(23292) <= 3586698;
srom_1(23293) <= 4068695;
srom_1(23294) <= 4570950;
srom_1(23295) <= 5091107;
srom_1(23296) <= 5626727;
srom_1(23297) <= 6175299;
srom_1(23298) <= 6734250;
srom_1(23299) <= 7300958;
srom_1(23300) <= 7872767;
srom_1(23301) <= 8446995;
srom_1(23302) <= 9020949;
srom_1(23303) <= 9591937;
srom_1(23304) <= 10157283;
srom_1(23305) <= 10714335;
srom_1(23306) <= 11260481;
srom_1(23307) <= 11793159;
srom_1(23308) <= 12309873;
srom_1(23309) <= 12808198;
srom_1(23310) <= 13285799;
srom_1(23311) <= 13740434;
srom_1(23312) <= 14169973;
srom_1(23313) <= 14572402;
srom_1(23314) <= 14945832;
srom_1(23315) <= 15288513;
srom_1(23316) <= 15598839;
srom_1(23317) <= 15875353;
srom_1(23318) <= 16116759;
srom_1(23319) <= 16321925;
srom_1(23320) <= 16489889;
srom_1(23321) <= 16619863;
srom_1(23322) <= 16711239;
srom_1(23323) <= 16763586;
srom_1(23324) <= 16776660;
srom_1(23325) <= 16750400;
srom_1(23326) <= 16684929;
srom_1(23327) <= 16580553;
srom_1(23328) <= 16437762;
srom_1(23329) <= 16257227;
srom_1(23330) <= 16039792;
srom_1(23331) <= 15786478;
srom_1(23332) <= 15498474;
srom_1(23333) <= 15177128;
srom_1(23334) <= 14823949;
srom_1(23335) <= 14440593;
srom_1(23336) <= 14028856;
srom_1(23337) <= 13590671;
srom_1(23338) <= 13128091;
srom_1(23339) <= 12643286;
srom_1(23340) <= 12138530;
srom_1(23341) <= 11616189;
srom_1(23342) <= 11078712;
srom_1(23343) <= 10528621;
srom_1(23344) <= 9968495;
srom_1(23345) <= 9400959;
srom_1(23346) <= 8828677;
srom_1(23347) <= 8254331;
srom_1(23348) <= 7680615;
srom_1(23349) <= 7110218;
srom_1(23350) <= 6545817;
srom_1(23351) <= 5990057;
srom_1(23352) <= 5445544;
srom_1(23353) <= 4914833;
srom_1(23354) <= 4400411;
srom_1(23355) <= 3904691;
srom_1(23356) <= 3429998;
srom_1(23357) <= 2978558;
srom_1(23358) <= 2552487;
srom_1(23359) <= 2153783;
srom_1(23360) <= 1784317;
srom_1(23361) <= 1445821;
srom_1(23362) <= 1139882;
srom_1(23363) <= 867934;
srom_1(23364) <= 631254;
srom_1(23365) <= 430951;
srom_1(23366) <= 267963;
srom_1(23367) <= 143056;
srom_1(23368) <= 56816;
srom_1(23369) <= 9646;
srom_1(23370) <= 1767;
srom_1(23371) <= 33218;
srom_1(23372) <= 103850;
srom_1(23373) <= 213332;
srom_1(23374) <= 361150;
srom_1(23375) <= 546613;
srom_1(23376) <= 768848;
srom_1(23377) <= 1026816;
srom_1(23378) <= 1319306;
srom_1(23379) <= 1644946;
srom_1(23380) <= 2002209;
srom_1(23381) <= 2389420;
srom_1(23382) <= 2804764;
srom_1(23383) <= 3246292;
srom_1(23384) <= 3711934;
srom_1(23385) <= 4199507;
srom_1(23386) <= 4706723;
srom_1(23387) <= 5231206;
srom_1(23388) <= 5770494;
srom_1(23389) <= 6322060;
srom_1(23390) <= 6883317;
srom_1(23391) <= 7451632;
srom_1(23392) <= 8024341;
srom_1(23393) <= 8598759;
srom_1(23394) <= 9172190;
srom_1(23395) <= 9741948;
srom_1(23396) <= 10305359;
srom_1(23397) <= 10859782;
srom_1(23398) <= 11402616;
srom_1(23399) <= 11931317;
srom_1(23400) <= 12443405;
srom_1(23401) <= 12936478;
srom_1(23402) <= 13408225;
srom_1(23403) <= 13856434;
srom_1(23404) <= 14279001;
srom_1(23405) <= 14673947;
srom_1(23406) <= 15039419;
srom_1(23407) <= 15373702;
srom_1(23408) <= 15675230;
srom_1(23409) <= 15942589;
srom_1(23410) <= 16174524;
srom_1(23411) <= 16369949;
srom_1(23412) <= 16527946;
srom_1(23413) <= 16647775;
srom_1(23414) <= 16728874;
srom_1(23415) <= 16770863;
srom_1(23416) <= 16773544;
srom_1(23417) <= 16736906;
srom_1(23418) <= 16661119;
srom_1(23419) <= 16546540;
srom_1(23420) <= 16393706;
srom_1(23421) <= 16203332;
srom_1(23422) <= 15976313;
srom_1(23423) <= 15713713;
srom_1(23424) <= 15416762;
srom_1(23425) <= 15086855;
srom_1(23426) <= 14725536;
srom_1(23427) <= 14334502;
srom_1(23428) <= 13915585;
srom_1(23429) <= 13470751;
srom_1(23430) <= 13002084;
srom_1(23431) <= 12511784;
srom_1(23432) <= 12002148;
srom_1(23433) <= 11475567;
srom_1(23434) <= 10934511;
srom_1(23435) <= 10381516;
srom_1(23436) <= 9819175;
srom_1(23437) <= 9250126;
srom_1(23438) <= 8677037;
srom_1(23439) <= 8102595;
srom_1(23440) <= 7529495;
srom_1(23441) <= 6960423;
srom_1(23442) <= 6398049;
srom_1(23443) <= 5845009;
srom_1(23444) <= 5303896;
srom_1(23445) <= 4777249;
srom_1(23446) <= 4267537;
srom_1(23447) <= 3777150;
srom_1(23448) <= 3308388;
srom_1(23449) <= 2863449;
srom_1(23450) <= 2444419;
srom_1(23451) <= 2053263;
srom_1(23452) <= 1691816;
srom_1(23453) <= 1361772;
srom_1(23454) <= 1064680;
srom_1(23455) <= 801932;
srom_1(23456) <= 574761;
srom_1(23457) <= 384231;
srom_1(23458) <= 231237;
srom_1(23459) <= 116495;
srom_1(23460) <= 40545;
srom_1(23461) <= 3741;
srom_1(23462) <= 6256;
srom_1(23463) <= 48080;
srom_1(23464) <= 129015;
srom_1(23465) <= 248682;
srom_1(23466) <= 406520;
srom_1(23467) <= 601788;
srom_1(23468) <= 833572;
srom_1(23469) <= 1100784;
srom_1(23470) <= 1402171;
srom_1(23471) <= 1736320;
srom_1(23472) <= 2101663;
srom_1(23473) <= 2496489;
srom_1(23474) <= 2918944;
srom_1(23475) <= 3367049;
srom_1(23476) <= 3838701;
srom_1(23477) <= 4331689;
srom_1(23478) <= 4843702;
srom_1(23479) <= 5372338;
srom_1(23480) <= 5915119;
srom_1(23481) <= 6469498;
srom_1(23482) <= 7032877;
srom_1(23483) <= 7602613;
srom_1(23484) <= 8176035;
srom_1(23485) <= 8750454;
srom_1(23486) <= 9323176;
srom_1(23487) <= 9891515;
srom_1(23488) <= 10452807;
srom_1(23489) <= 11004419;
srom_1(23490) <= 11543765;
srom_1(23491) <= 12068315;
srom_1(23492) <= 12575609;
srom_1(23493) <= 13063270;
srom_1(23494) <= 13529009;
srom_1(23495) <= 13970643;
srom_1(23496) <= 14386101;
srom_1(23497) <= 14773435;
srom_1(23498) <= 15130828;
srom_1(23499) <= 15456604;
srom_1(23500) <= 15749236;
srom_1(23501) <= 16007352;
srom_1(23502) <= 16229741;
srom_1(23503) <= 16415360;
srom_1(23504) <= 16563338;
srom_1(23505) <= 16672983;
srom_1(23506) <= 16743779;
srom_1(23507) <= 16775396;
srom_1(23508) <= 16767683;
srom_1(23509) <= 16720678;
srom_1(23510) <= 16634601;
srom_1(23511) <= 16509856;
srom_1(23512) <= 16347028;
srom_1(23513) <= 16146880;
srom_1(23514) <= 15910350;
srom_1(23515) <= 15638549;
srom_1(23516) <= 15332750;
srom_1(23517) <= 14994388;
srom_1(23518) <= 14625049;
srom_1(23519) <= 14226465;
srom_1(23520) <= 13800505;
srom_1(23521) <= 13349167;
srom_1(23522) <= 12874567;
srom_1(23523) <= 12378931;
srom_1(23524) <= 11864583;
srom_1(23525) <= 11333935;
srom_1(23526) <= 10789476;
srom_1(23527) <= 10233758;
srom_1(23528) <= 9669387;
srom_1(23529) <= 9099010;
srom_1(23530) <= 8525302;
srom_1(23531) <= 7950953;
srom_1(23532) <= 7378656;
srom_1(23533) <= 6811096;
srom_1(23534) <= 6250932;
srom_1(23535) <= 5700793;
srom_1(23536) <= 5163259;
srom_1(23537) <= 4640848;
srom_1(23538) <= 4136013;
srom_1(23539) <= 3651119;
srom_1(23540) <= 3188441;
srom_1(23541) <= 2750148;
srom_1(23542) <= 2338296;
srom_1(23543) <= 1954816;
srom_1(23544) <= 1601507;
srom_1(23545) <= 1280024;
srom_1(23546) <= 991876;
srom_1(23547) <= 738414;
srom_1(23548) <= 520826;
srom_1(23549) <= 340132;
srom_1(23550) <= 197181;
srom_1(23551) <= 92643;
srom_1(23552) <= 27006;
srom_1(23553) <= 581;
srom_1(23554) <= 13489;
srom_1(23555) <= 65672;
srom_1(23556) <= 156883;
srom_1(23557) <= 286696;
srom_1(23558) <= 454502;
srom_1(23559) <= 659513;
srom_1(23560) <= 900769;
srom_1(23561) <= 1177138;
srom_1(23562) <= 1487323;
srom_1(23563) <= 1829872;
srom_1(23564) <= 2203176;
srom_1(23565) <= 2605486;
srom_1(23566) <= 3034915;
srom_1(23567) <= 3489450;
srom_1(23568) <= 3966958;
srom_1(23569) <= 4465201;
srom_1(23570) <= 4981842;
srom_1(23571) <= 5514458;
srom_1(23572) <= 6060553;
srom_1(23573) <= 6617564;
srom_1(23574) <= 7182880;
srom_1(23575) <= 7753851;
srom_1(23576) <= 8327798;
srom_1(23577) <= 8902030;
srom_1(23578) <= 9473855;
srom_1(23579) <= 10040590;
srom_1(23580) <= 10599579;
srom_1(23581) <= 11148200;
srom_1(23582) <= 11683880;
srom_1(23583) <= 12204108;
srom_1(23584) <= 12706443;
srom_1(23585) <= 13188530;
srom_1(23586) <= 13648109;
srom_1(23587) <= 14083025;
srom_1(23588) <= 14491237;
srom_1(23589) <= 14870832;
srom_1(23590) <= 15220029;
srom_1(23591) <= 15537192;
srom_1(23592) <= 15820832;
srom_1(23593) <= 16069621;
srom_1(23594) <= 16282390;
srom_1(23595) <= 16458143;
srom_1(23596) <= 16596054;
srom_1(23597) <= 16695479;
srom_1(23598) <= 16755949;
srom_1(23599) <= 16777182;
srom_1(23600) <= 16759079;
srom_1(23601) <= 16701723;
srom_1(23602) <= 16605384;
srom_1(23603) <= 16470514;
srom_1(23604) <= 16297745;
srom_1(23605) <= 16087887;
srom_1(23606) <= 15841925;
srom_1(23607) <= 15561012;
srom_1(23608) <= 15246464;
srom_1(23609) <= 14899758;
srom_1(23610) <= 14522519;
srom_1(23611) <= 14116516;
srom_1(23612) <= 13683653;
srom_1(23613) <= 13225959;
srom_1(23614) <= 12745581;
srom_1(23615) <= 12244772;
srom_1(23616) <= 11725881;
srom_1(23617) <= 11191339;
srom_1(23618) <= 10643655;
srom_1(23619) <= 10085396;
srom_1(23620) <= 9519180;
srom_1(23621) <= 8947662;
srom_1(23622) <= 8373523;
srom_1(23623) <= 7799454;
srom_1(23624) <= 7228149;
srom_1(23625) <= 6662285;
srom_1(23626) <= 6104516;
srom_1(23627) <= 5557458;
srom_1(23628) <= 5023677;
srom_1(23629) <= 4505674;
srom_1(23630) <= 4005881;
srom_1(23631) <= 3526639;
srom_1(23632) <= 3070197;
srom_1(23633) <= 2638694;
srom_1(23634) <= 2234155;
srom_1(23635) <= 1858476;
srom_1(23636) <= 1513420;
srom_1(23637) <= 1200603;
srom_1(23638) <= 921493;
srom_1(23639) <= 677400;
srom_1(23640) <= 469466;
srom_1(23641) <= 298669;
srom_1(23642) <= 165808;
srom_1(23643) <= 71506;
srom_1(23644) <= 16206;
srom_1(23645) <= 167;
srom_1(23646) <= 23465;
srom_1(23647) <= 85989;
srom_1(23648) <= 187447;
srom_1(23649) <= 327364;
srom_1(23650) <= 505082;
srom_1(23651) <= 719769;
srom_1(23652) <= 970417;
srom_1(23653) <= 1255852;
srom_1(23654) <= 1574735;
srom_1(23655) <= 1925571;
srom_1(23656) <= 2306714;
srom_1(23657) <= 2716377;
srom_1(23658) <= 3152639;
srom_1(23659) <= 3613454;
srom_1(23660) <= 4096662;
srom_1(23661) <= 4599996;
srom_1(23662) <= 5121096;
srom_1(23663) <= 5657519;
srom_1(23664) <= 6206749;
srom_1(23665) <= 6766210;
srom_1(23666) <= 7333279;
srom_1(23667) <= 7905297;
srom_1(23668) <= 8479581;
srom_1(23669) <= 9053439;
srom_1(23670) <= 9624179;
srom_1(23671) <= 10189125;
srom_1(23672) <= 10745628;
srom_1(23673) <= 11291078;
srom_1(23674) <= 11822917;
srom_1(23675) <= 12338652;
srom_1(23676) <= 12835863;
srom_1(23677) <= 13312220;
srom_1(23678) <= 13765488;
srom_1(23679) <= 14193542;
srom_1(23680) <= 14594375;
srom_1(23681) <= 14966107;
srom_1(23682) <= 15306995;
srom_1(23683) <= 15615440;
srom_1(23684) <= 15889995;
srom_1(23685) <= 16129375;
srom_1(23686) <= 16332455;
srom_1(23687) <= 16498284;
srom_1(23688) <= 16626083;
srom_1(23689) <= 16715255;
srom_1(23690) <= 16765380;
srom_1(23691) <= 16776223;
srom_1(23692) <= 16747734;
srom_1(23693) <= 16680046;
srom_1(23694) <= 16573476;
srom_1(23695) <= 16428525;
srom_1(23696) <= 16245872;
srom_1(23697) <= 16026374;
srom_1(23698) <= 15771059;
srom_1(23699) <= 15481126;
srom_1(23700) <= 15157933;
srom_1(23701) <= 14802997;
srom_1(23702) <= 14417981;
srom_1(23703) <= 14004692;
srom_1(23704) <= 13565067;
srom_1(23705) <= 13101167;
srom_1(23706) <= 12615169;
srom_1(23707) <= 12109351;
srom_1(23708) <= 11586085;
srom_1(23709) <= 11047825;
srom_1(23710) <= 10497095;
srom_1(23711) <= 9936478;
srom_1(23712) <= 9368602;
srom_1(23713) <= 8796131;
srom_1(23714) <= 8221748;
srom_1(23715) <= 7648148;
srom_1(23716) <= 7078021;
srom_1(23717) <= 6514039;
srom_1(23718) <= 5958847;
srom_1(23719) <= 5415050;
srom_1(23720) <= 4885197;
srom_1(23721) <= 4371772;
srom_1(23722) <= 3877183;
srom_1(23723) <= 3403751;
srom_1(23724) <= 2953694;
srom_1(23725) <= 2529123;
srom_1(23726) <= 2132029;
srom_1(23727) <= 1764274;
srom_1(23728) <= 1427584;
srom_1(23729) <= 1123535;
srom_1(23730) <= 853556;
srom_1(23731) <= 618910;
srom_1(23732) <= 420700;
srom_1(23733) <= 259854;
srom_1(23734) <= 137126;
srom_1(23735) <= 53092;
srom_1(23736) <= 8147;
srom_1(23737) <= 2500;
srom_1(23738) <= 36178;
srom_1(23739) <= 109024;
srom_1(23740) <= 220696;
srom_1(23741) <= 370670;
srom_1(23742) <= 558243;
srom_1(23743) <= 782535;
srom_1(23744) <= 1042494;
srom_1(23745) <= 1336902;
srom_1(23746) <= 1664378;
srom_1(23747) <= 2023386;
srom_1(23748) <= 2412243;
srom_1(23749) <= 2829125;
srom_1(23750) <= 3272077;
srom_1(23751) <= 3739023;
srom_1(23752) <= 4227772;
srom_1(23753) <= 4736032;
srom_1(23754) <= 5261421;
srom_1(23755) <= 5801474;
srom_1(23756) <= 6353659;
srom_1(23757) <= 6915387;
srom_1(23758) <= 7484023;
srom_1(23759) <= 8056901;
srom_1(23760) <= 8631334;
srom_1(23761) <= 9204630;
srom_1(23762) <= 9774098;
srom_1(23763) <= 10337070;
srom_1(23764) <= 10890905;
srom_1(23765) <= 11433005;
srom_1(23766) <= 11960829;
srom_1(23767) <= 12471902;
srom_1(23768) <= 12963827;
srom_1(23769) <= 13434297;
srom_1(23770) <= 13881106;
srom_1(23771) <= 14302159;
srom_1(23772) <= 14695481;
srom_1(23773) <= 15059228;
srom_1(23774) <= 15391695;
srom_1(23775) <= 15691321;
srom_1(23776) <= 15956703;
srom_1(23777) <= 16186595;
srom_1(23778) <= 16379919;
srom_1(23779) <= 16535770;
srom_1(23780) <= 16653415;
srom_1(23781) <= 16732305;
srom_1(23782) <= 16772067;
srom_1(23783) <= 16772517;
srom_1(23784) <= 16733652;
srom_1(23785) <= 16655654;
srom_1(23786) <= 16538889;
srom_1(23787) <= 16383905;
srom_1(23788) <= 16191427;
srom_1(23789) <= 15962360;
srom_1(23790) <= 15697777;
srom_1(23791) <= 15398918;
srom_1(23792) <= 15067186;
srom_1(23793) <= 14704136;
srom_1(23794) <= 14311470;
srom_1(23795) <= 13891029;
srom_1(23796) <= 13444786;
srom_1(23797) <= 12974833;
srom_1(23798) <= 12483373;
srom_1(23799) <= 11972712;
srom_1(23800) <= 11445243;
srom_1(23801) <= 10903441;
srom_1(23802) <= 10349846;
srom_1(23803) <= 9787054;
srom_1(23804) <= 9217704;
srom_1(23805) <= 8644466;
srom_1(23806) <= 8070029;
srom_1(23807) <= 7497085;
srom_1(23808) <= 6928322;
srom_1(23809) <= 6366407;
srom_1(23810) <= 5813974;
srom_1(23811) <= 5273615;
srom_1(23812) <= 4747863;
srom_1(23813) <= 4239184;
srom_1(23814) <= 3749963;
srom_1(23815) <= 3282494;
srom_1(23816) <= 2838970;
srom_1(23817) <= 2421469;
srom_1(23818) <= 2031951;
srom_1(23819) <= 1672241;
srom_1(23820) <= 1344026;
srom_1(23821) <= 1048846;
srom_1(23822) <= 788085;
srom_1(23823) <= 562965;
srom_1(23824) <= 374542;
srom_1(23825) <= 223700;
srom_1(23826) <= 111146;
srom_1(23827) <= 37407;
srom_1(23828) <= 2831;
srom_1(23829) <= 7578;
srom_1(23830) <= 51627;
srom_1(23831) <= 134770;
srom_1(23832) <= 256619;
srom_1(23833) <= 416601;
srom_1(23834) <= 613967;
srom_1(23835) <= 847791;
srom_1(23836) <= 1116976;
srom_1(23837) <= 1420261;
srom_1(23838) <= 1756222;
srom_1(23839) <= 2123285;
srom_1(23840) <= 2519729;
srom_1(23841) <= 2943693;
srom_1(23842) <= 3393190;
srom_1(23843) <= 3866113;
srom_1(23844) <= 4360243;
srom_1(23845) <= 4873264;
srom_1(23846) <= 5402769;
srom_1(23847) <= 5946276;
srom_1(23848) <= 6501236;
srom_1(23849) <= 7065046;
srom_1(23850) <= 7635063;
srom_1(23851) <= 8208614;
srom_1(23852) <= 8783008;
srom_1(23853) <= 9355553;
srom_1(23854) <= 9923564;
srom_1(23855) <= 10484377;
srom_1(23856) <= 11035362;
srom_1(23857) <= 11573936;
srom_1(23858) <= 12097572;
srom_1(23859) <= 12603816;
srom_1(23860) <= 13090293;
srom_1(23861) <= 13554723;
srom_1(23862) <= 13994926;
srom_1(23863) <= 14408840;
srom_1(23864) <= 14794523;
srom_1(23865) <= 15150166;
srom_1(23866) <= 15474102;
srom_1(23867) <= 15764812;
srom_1(23868) <= 16020932;
srom_1(23869) <= 16241261;
srom_1(23870) <= 16424767;
srom_1(23871) <= 16570588;
srom_1(23872) <= 16678042;
srom_1(23873) <= 16746623;
srom_1(23874) <= 16776011;
srom_1(23875) <= 16766067;
srom_1(23876) <= 16716838;
srom_1(23877) <= 16628556;
srom_1(23878) <= 16501633;
srom_1(23879) <= 16336666;
srom_1(23880) <= 16134428;
srom_1(23881) <= 15895867;
srom_1(23882) <= 15622101;
srom_1(23883) <= 15314416;
srom_1(23884) <= 14974252;
srom_1(23885) <= 14603207;
srom_1(23886) <= 14203019;
srom_1(23887) <= 13775565;
srom_1(23888) <= 13322850;
srom_1(23889) <= 12846997;
srom_1(23890) <= 12350236;
srom_1(23891) <= 11834899;
srom_1(23892) <= 11303400;
srom_1(23893) <= 10758233;
srom_1(23894) <= 10201954;
srom_1(23895) <= 9637172;
srom_1(23896) <= 9066534;
srom_1(23897) <= 8492718;
srom_1(23898) <= 7918413;
srom_1(23899) <= 7346313;
srom_1(23900) <= 6779101;
srom_1(23901) <= 6219437;
srom_1(23902) <= 5669944;
srom_1(23903) <= 5133200;
srom_1(23904) <= 4611722;
srom_1(23905) <= 4107955;
srom_1(23906) <= 3624262;
srom_1(23907) <= 3162910;
srom_1(23908) <= 2726063;
srom_1(23909) <= 2315770;
srom_1(23910) <= 1933954;
srom_1(23911) <= 1582406;
srom_1(23912) <= 1262776;
srom_1(23913) <= 976560;
srom_1(23914) <= 725102;
srom_1(23915) <= 509581;
srom_1(23916) <= 331008;
srom_1(23917) <= 190219;
srom_1(23918) <= 87875;
srom_1(23919) <= 24457;
srom_1(23920) <= 260;
srom_1(23921) <= 15400;
srom_1(23922) <= 69804;
srom_1(23923) <= 163219;
srom_1(23924) <= 295204;
srom_1(23925) <= 465143;
srom_1(23926) <= 672237;
srom_1(23927) <= 915516;
srom_1(23928) <= 1193839;
srom_1(23929) <= 1505901;
srom_1(23930) <= 1850238;
srom_1(23931) <= 2225236;
srom_1(23932) <= 2629136;
srom_1(23933) <= 3060044;
srom_1(23934) <= 3515939;
srom_1(23935) <= 3994684;
srom_1(23936) <= 4494034;
srom_1(23937) <= 5011647;
srom_1(23938) <= 5545095;
srom_1(23939) <= 6091878;
srom_1(23940) <= 6649430;
srom_1(23941) <= 7215139;
srom_1(23942) <= 7786350;
srom_1(23943) <= 8360385;
srom_1(23944) <= 8934553;
srom_1(23945) <= 9506161;
srom_1(23946) <= 10072528;
srom_1(23947) <= 10630998;
srom_1(23948) <= 11178953;
srom_1(23949) <= 11713823;
srom_1(23950) <= 12233101;
srom_1(23951) <= 12734350;
srom_1(23952) <= 13215220;
srom_1(23953) <= 13673457;
srom_1(23954) <= 14106911;
srom_1(23955) <= 14513550;
srom_1(23956) <= 14891467;
srom_1(23957) <= 15238890;
srom_1(23958) <= 15554190;
srom_1(23959) <= 15835887;
srom_1(23960) <= 16082662;
srom_1(23961) <= 16293357;
srom_1(23962) <= 16466984;
srom_1(23963) <= 16602728;
srom_1(23964) <= 16699954;
srom_1(23965) <= 16758205;
srom_1(23966) <= 16777208;
srom_1(23967) <= 16756874;
srom_1(23968) <= 16697298;
srom_1(23969) <= 16598760;
srom_1(23970) <= 16461722;
srom_1(23971) <= 16286826;
srom_1(23972) <= 16074892;
srom_1(23973) <= 15826915;
srom_1(23974) <= 15544057;
srom_1(23975) <= 15227645;
srom_1(23976) <= 14879162;
srom_1(23977) <= 14500243;
srom_1(23978) <= 14092664;
srom_1(23979) <= 13658337;
srom_1(23980) <= 13199299;
srom_1(23981) <= 12717701;
srom_1(23982) <= 12215803;
srom_1(23983) <= 11695958;
srom_1(23984) <= 11160603;
srom_1(23985) <= 10612250;
srom_1(23986) <= 10053469;
srom_1(23987) <= 9486881;
srom_1(23988) <= 8915142;
srom_1(23989) <= 8340935;
srom_1(23990) <= 7766951;
srom_1(23991) <= 7195883;
srom_1(23992) <= 6630407;
srom_1(23993) <= 6073177;
srom_1(23994) <= 5526804;
srom_1(23995) <= 4993851;
srom_1(23996) <= 4476817;
srom_1(23997) <= 3978127;
srom_1(23998) <= 3500120;
srom_1(23999) <= 3045036;
srom_1(24000) <= 2615010;
srom_1(24001) <= 2212058;
srom_1(24002) <= 1838070;
srom_1(24003) <= 1494800;
srom_1(24004) <= 1183858;
srom_1(24005) <= 906701;
srom_1(24006) <= 664629;
srom_1(24007) <= 458777;
srom_1(24008) <= 290112;
srom_1(24009) <= 159422;
srom_1(24010) <= 67323;
srom_1(24011) <= 14244;
srom_1(24012) <= 436;
srom_1(24013) <= 25963;
srom_1(24014) <= 90706;
srom_1(24015) <= 194360;
srom_1(24016) <= 336439;
srom_1(24017) <= 516278;
srom_1(24018) <= 733033;
srom_1(24019) <= 985688;
srom_1(24020) <= 1273058;
srom_1(24021) <= 1593794;
srom_1(24022) <= 1946394;
srom_1(24023) <= 2329204;
srom_1(24024) <= 2740428;
srom_1(24025) <= 3178139;
srom_1(24026) <= 3640283;
srom_1(24027) <= 4124694;
srom_1(24028) <= 4629100;
srom_1(24029) <= 5151135;
srom_1(24030) <= 5688352;
srom_1(24031) <= 6238231;
srom_1(24032) <= 6798195;
srom_1(24033) <= 7365616;
srom_1(24034) <= 7937834;
srom_1(24035) <= 8512166;
srom_1(24036) <= 9085919;
srom_1(24037) <= 9656402;
srom_1(24038) <= 10220940;
srom_1(24039) <= 10776885;
srom_1(24040) <= 11321631;
srom_1(24041) <= 11852623;
srom_1(24042) <= 12367370;
srom_1(24043) <= 12863461;
srom_1(24044) <= 13338567;
srom_1(24045) <= 13790460;
srom_1(24046) <= 14217023;
srom_1(24047) <= 14616255;
srom_1(24048) <= 14986282;
srom_1(24049) <= 15325371;
srom_1(24050) <= 15631931;
srom_1(24051) <= 15904525;
srom_1(24052) <= 16141874;
srom_1(24053) <= 16342865;
srom_1(24054) <= 16506556;
srom_1(24055) <= 16632179;
srom_1(24056) <= 16719145;
srom_1(24057) <= 16767047;
srom_1(24058) <= 16775659;
srom_1(24059) <= 16744941;
srom_1(24060) <= 16675037;
srom_1(24061) <= 16566276;
srom_1(24062) <= 16419167;
srom_1(24063) <= 16234399;
srom_1(24064) <= 16012840;
srom_1(24065) <= 15755529;
srom_1(24066) <= 15463671;
srom_1(24067) <= 15138636;
srom_1(24068) <= 14781948;
srom_1(24069) <= 14395279;
srom_1(24070) <= 13980443;
srom_1(24071) <= 13539384;
srom_1(24072) <= 13074172;
srom_1(24073) <= 12586988;
srom_1(24074) <= 12080116;
srom_1(24075) <= 11555934;
srom_1(24076) <= 11016898;
srom_1(24077) <= 10465538;
srom_1(24078) <= 9904438;
srom_1(24079) <= 9336230;
srom_1(24080) <= 8763578;
srom_1(24081) <= 8189168;
srom_1(24082) <= 7615693;
srom_1(24083) <= 7045843;
srom_1(24084) <= 6482289;
srom_1(24085) <= 5927675;
srom_1(24086) <= 5384601;
srom_1(24087) <= 4855613;
srom_1(24088) <= 4343193;
srom_1(24089) <= 3849744;
srom_1(24090) <= 3377578;
srom_1(24091) <= 2928911;
srom_1(24092) <= 2505847;
srom_1(24093) <= 2110369;
srom_1(24094) <= 1744331;
srom_1(24095) <= 1409451;
srom_1(24096) <= 1107299;
srom_1(24097) <= 839291;
srom_1(24098) <= 606684;
srom_1(24099) <= 410569;
srom_1(24100) <= 251867;
srom_1(24101) <= 131320;
srom_1(24102) <= 49494;
srom_1(24103) <= 6774;
srom_1(24104) <= 3359;
srom_1(24105) <= 39265;
srom_1(24106) <= 114324;
srom_1(24107) <= 228184;
srom_1(24108) <= 380311;
srom_1(24109) <= 569991;
srom_1(24110) <= 796336;
srom_1(24111) <= 1058283;
srom_1(24112) <= 1354605;
srom_1(24113) <= 1683912;
srom_1(24114) <= 2044660;
srom_1(24115) <= 2435156;
srom_1(24116) <= 2853570;
srom_1(24117) <= 3297940;
srom_1(24118) <= 3766182;
srom_1(24119) <= 4256100;
srom_1(24120) <= 4765396;
srom_1(24121) <= 5291683;
srom_1(24122) <= 5832493;
srom_1(24123) <= 6385289;
srom_1(24124) <= 6947479;
srom_1(24125) <= 7516428;
srom_1(24126) <= 8089466;
srom_1(24127) <= 8663907;
srom_1(24128) <= 9237057;
srom_1(24129) <= 9806228;
srom_1(24130) <= 10368752;
srom_1(24131) <= 10921990;
srom_1(24132) <= 11463348;
srom_1(24133) <= 11990288;
srom_1(24134) <= 12500338;
srom_1(24135) <= 12991107;
srom_1(24136) <= 13460293;
srom_1(24137) <= 13905696;
srom_1(24138) <= 14325228;
srom_1(24139) <= 14716920;
srom_1(24140) <= 15078938;
srom_1(24141) <= 15409581;
srom_1(24142) <= 15707302;
srom_1(24143) <= 15970702;
srom_1(24144) <= 16198547;
srom_1(24145) <= 16389769;
srom_1(24146) <= 16543470;
srom_1(24147) <= 16658931;
srom_1(24148) <= 16735609;
srom_1(24149) <= 16773145;
srom_1(24150) <= 16771364;
srom_1(24151) <= 16730272;
srom_1(24152) <= 16650064;
srom_1(24153) <= 16531115;
srom_1(24154) <= 16373983;
srom_1(24155) <= 16179404;
srom_1(24156) <= 15948292;
srom_1(24157) <= 15681730;
srom_1(24158) <= 15380968;
srom_1(24159) <= 15047417;
srom_1(24160) <= 14682640;
srom_1(24161) <= 14288348;
srom_1(24162) <= 13866390;
srom_1(24163) <= 13418745;
srom_1(24164) <= 12947512;
srom_1(24165) <= 12454901;
srom_1(24166) <= 11943221;
srom_1(24167) <= 11414873;
srom_1(24168) <= 10872333;
srom_1(24169) <= 10318146;
srom_1(24170) <= 9754911;
srom_1(24171) <= 9185269;
srom_1(24172) <= 8611892;
srom_1(24173) <= 8037467;
srom_1(24174) <= 7464688;
srom_1(24175) <= 6896243;
srom_1(24176) <= 6334795;
srom_1(24177) <= 5782979;
srom_1(24178) <= 5243381;
srom_1(24179) <= 4718532;
srom_1(24180) <= 4210894;
srom_1(24181) <= 3722846;
srom_1(24182) <= 3256678;
srom_1(24183) <= 2814574;
srom_1(24184) <= 2398610;
srom_1(24185) <= 2010735;
srom_1(24186) <= 1652767;
srom_1(24187) <= 1326387;
srom_1(24188) <= 1033123;
srom_1(24189) <= 774352;
srom_1(24190) <= 551287;
srom_1(24191) <= 364974;
srom_1(24192) <= 216286;
srom_1(24193) <= 105921;
srom_1(24194) <= 34396;
srom_1(24195) <= 2047;
srom_1(24196) <= 9026;
srom_1(24197) <= 55299;
srom_1(24198) <= 140651;
srom_1(24199) <= 264679;
srom_1(24200) <= 426804;
srom_1(24201) <= 626264;
srom_1(24202) <= 862124;
srom_1(24203) <= 1133279;
srom_1(24204) <= 1438456;
srom_1(24205) <= 1776225;
srom_1(24206) <= 2145002;
srom_1(24207) <= 2543057;
srom_1(24208) <= 2968524;
srom_1(24209) <= 3419408;
srom_1(24210) <= 3893594;
srom_1(24211) <= 4388858;
srom_1(24212) <= 4902879;
srom_1(24213) <= 5433245;
srom_1(24214) <= 5977470;
srom_1(24215) <= 6533002;
srom_1(24216) <= 7097236;
srom_1(24217) <= 7667525;
srom_1(24218) <= 8241195;
srom_1(24219) <= 8815557;
srom_1(24220) <= 9387917;
srom_1(24221) <= 9955590;
srom_1(24222) <= 10515916;
srom_1(24223) <= 11066265;
srom_1(24224) <= 11604059;
srom_1(24225) <= 12126773;
srom_1(24226) <= 12631959;
srom_1(24227) <= 13117246;
srom_1(24228) <= 13580358;
srom_1(24229) <= 14019125;
srom_1(24230) <= 14431488;
srom_1(24231) <= 14815514;
srom_1(24232) <= 15169402;
srom_1(24233) <= 15491493;
srom_1(24234) <= 15780276;
srom_1(24235) <= 16034397;
srom_1(24236) <= 16252663;
srom_1(24237) <= 16434053;
srom_1(24238) <= 16577715;
srom_1(24239) <= 16682975;
srom_1(24240) <= 16749340;
srom_1(24241) <= 16776499;
srom_1(24242) <= 16764324;
srom_1(24243) <= 16712873;
srom_1(24244) <= 16622386;
srom_1(24245) <= 16493288;
srom_1(24246) <= 16326184;
srom_1(24247) <= 16121859;
srom_1(24248) <= 15881269;
srom_1(24249) <= 15605544;
srom_1(24250) <= 15295976;
srom_1(24251) <= 14954018;
srom_1(24252) <= 14581271;
srom_1(24253) <= 14179485;
srom_1(24254) <= 13750544;
srom_1(24255) <= 13296459;
srom_1(24256) <= 12819359;
srom_1(24257) <= 12321482;
srom_1(24258) <= 11805162;
srom_1(24259) <= 11272821;
srom_1(24260) <= 10726955;
srom_1(24261) <= 10170123;
srom_1(24262) <= 9604937;
srom_1(24263) <= 9034048;
srom_1(24264) <= 8460132;
srom_1(24265) <= 7885880;
srom_1(24266) <= 7313986;
srom_1(24267) <= 6747131;
srom_1(24268) <= 6187974;
srom_1(24269) <= 5639136;
srom_1(24270) <= 5103191;
srom_1(24271) <= 4582653;
srom_1(24272) <= 4079962;
srom_1(24273) <= 3597476;
srom_1(24274) <= 3137457;
srom_1(24275) <= 2702062;
srom_1(24276) <= 2293334;
srom_1(24277) <= 1913189;
srom_1(24278) <= 1563409;
srom_1(24279) <= 1245635;
srom_1(24280) <= 961356;
srom_1(24281) <= 711907;
srom_1(24282) <= 498456;
srom_1(24283) <= 322005;
srom_1(24284) <= 183380;
srom_1(24285) <= 83233;
srom_1(24286) <= 22033;
srom_1(24287) <= 67;
srom_1(24288) <= 17437;
srom_1(24289) <= 74062;
srom_1(24290) <= 169678;
srom_1(24291) <= 303834;
srom_1(24292) <= 475903;
srom_1(24293) <= 685078;
srom_1(24294) <= 930376;
srom_1(24295) <= 1210649;
srom_1(24296) <= 1524582;
srom_1(24297) <= 1870703;
srom_1(24298) <= 2247388;
srom_1(24299) <= 2652872;
srom_1(24300) <= 3085253;
srom_1(24301) <= 3542502;
srom_1(24302) <= 4022477;
srom_1(24303) <= 4522926;
srom_1(24304) <= 5041503;
srom_1(24305) <= 5575775;
srom_1(24306) <= 6123238;
srom_1(24307) <= 6681323;
srom_1(24308) <= 7247415;
srom_1(24309) <= 7818858;
srom_1(24310) <= 8392973;
srom_1(24311) <= 8967068;
srom_1(24312) <= 9538449;
srom_1(24313) <= 10104439;
srom_1(24314) <= 10662383;
srom_1(24315) <= 11209664;
srom_1(24316) <= 11743716;
srom_1(24317) <= 12262036;
srom_1(24318) <= 12762191;
srom_1(24319) <= 13241837;
srom_1(24320) <= 13698724;
srom_1(24321) <= 14130711;
srom_1(24322) <= 14535770;
srom_1(24323) <= 14912004;
srom_1(24324) <= 15257647;
srom_1(24325) <= 15571079;
srom_1(24326) <= 15850830;
srom_1(24327) <= 16095588;
srom_1(24328) <= 16304205;
srom_1(24329) <= 16475703;
srom_1(24330) <= 16609278;
srom_1(24331) <= 16704304;
srom_1(24332) <= 16760334;
srom_1(24333) <= 16777107;
srom_1(24334) <= 16754543;
srom_1(24335) <= 16692748;
srom_1(24336) <= 16592012;
srom_1(24337) <= 16452808;
srom_1(24338) <= 16275787;
srom_1(24339) <= 16061781;
srom_1(24340) <= 15811793;
srom_1(24341) <= 15526995;
srom_1(24342) <= 15208723;
srom_1(24343) <= 14858469;
srom_1(24344) <= 14477875;
srom_1(24345) <= 14068727;
srom_1(24346) <= 13632943;
srom_1(24347) <= 13172566;
srom_1(24348) <= 12689755;
srom_1(24349) <= 12186775;
srom_1(24350) <= 11665985;
srom_1(24351) <= 11129825;
srom_1(24352) <= 10580811;
srom_1(24353) <= 10021517;
srom_1(24354) <= 9454565;
srom_1(24355) <= 8882615;
srom_1(24356) <= 8308348;
srom_1(24357) <= 7734458;
srom_1(24358) <= 7163635;
srom_1(24359) <= 6598557;
srom_1(24360) <= 6041872;
srom_1(24361) <= 5496193;
srom_1(24362) <= 4964077;
srom_1(24363) <= 4448019;
srom_1(24364) <= 3950441;
srom_1(24365) <= 3473674;
srom_1(24366) <= 3019955;
srom_1(24367) <= 2591412;
srom_1(24368) <= 2190054;
srom_1(24369) <= 1817763;
srom_1(24370) <= 1476285;
srom_1(24371) <= 1167221;
srom_1(24372) <= 892021;
srom_1(24373) <= 651974;
srom_1(24374) <= 448208;
srom_1(24375) <= 281677;
srom_1(24376) <= 153161;
srom_1(24377) <= 63265;
srom_1(24378) <= 12409;
srom_1(24379) <= 832;
srom_1(24380) <= 28588;
srom_1(24381) <= 95548;
srom_1(24382) <= 201396;
srom_1(24383) <= 345637;
srom_1(24384) <= 527594;
srom_1(24385) <= 746414;
srom_1(24386) <= 1001071;
srom_1(24387) <= 1290370;
srom_1(24388) <= 1612956;
srom_1(24389) <= 1967315;
srom_1(24390) <= 2351785;
srom_1(24391) <= 2764565;
srom_1(24392) <= 3203717;
srom_1(24393) <= 3667183;
srom_1(24394) <= 4152790;
srom_1(24395) <= 4658260;
srom_1(24396) <= 5181222;
srom_1(24397) <= 5719226;
srom_1(24398) <= 6269746;
srom_1(24399) <= 6830203;
srom_1(24400) <= 7397968;
srom_1(24401) <= 7970378;
srom_1(24402) <= 8544750;
srom_1(24403) <= 9118389;
srom_1(24404) <= 9688606;
srom_1(24405) <= 10252727;
srom_1(24406) <= 10808106;
srom_1(24407) <= 11352139;
srom_1(24408) <= 11882276;
srom_1(24409) <= 12396029;
srom_1(24410) <= 12890991;
srom_1(24411) <= 13364839;
srom_1(24412) <= 13815352;
srom_1(24413) <= 14240416;
srom_1(24414) <= 14638040;
srom_1(24415) <= 15006358;
srom_1(24416) <= 15343643;
srom_1(24417) <= 15648314;
srom_1(24418) <= 15918941;
srom_1(24419) <= 16154256;
srom_1(24420) <= 16353155;
srom_1(24421) <= 16514706;
srom_1(24422) <= 16638151;
srom_1(24423) <= 16722910;
srom_1(24424) <= 16768587;
srom_1(24425) <= 16774968;
srom_1(24426) <= 16742022;
srom_1(24427) <= 16669904;
srom_1(24428) <= 16558952;
srom_1(24429) <= 16409687;
srom_1(24430) <= 16222808;
srom_1(24431) <= 15999192;
srom_1(24432) <= 15739887;
srom_1(24433) <= 15446109;
srom_1(24434) <= 15119237;
srom_1(24435) <= 14760802;
srom_1(24436) <= 14372486;
srom_1(24437) <= 13956109;
srom_1(24438) <= 13513624;
srom_1(24439) <= 13047107;
srom_1(24440) <= 12558744;
srom_1(24441) <= 12050826;
srom_1(24442) <= 11525734;
srom_1(24443) <= 10985931;
srom_1(24444) <= 10433949;
srom_1(24445) <= 9872375;
srom_1(24446) <= 9303844;
srom_1(24447) <= 8731020;
srom_1(24448) <= 8156591;
srom_1(24449) <= 7583250;
srom_1(24450) <= 7013686;
srom_1(24451) <= 6450569;
srom_1(24452) <= 5896540;
srom_1(24453) <= 5354197;
srom_1(24454) <= 4826083;
srom_1(24455) <= 4314676;
srom_1(24456) <= 3822372;
srom_1(24457) <= 3351482;
srom_1(24458) <= 2904212;
srom_1(24459) <= 2482660;
srom_1(24460) <= 2088803;
srom_1(24461) <= 1724488;
srom_1(24462) <= 1391424;
srom_1(24463) <= 1091172;
srom_1(24464) <= 825139;
srom_1(24465) <= 594575;
srom_1(24466) <= 400559;
srom_1(24467) <= 244003;
srom_1(24468) <= 125639;
srom_1(24469) <= 46023;
srom_1(24470) <= 5528;
srom_1(24471) <= 4344;
srom_1(24472) <= 42477;
srom_1(24473) <= 119748;
srom_1(24474) <= 235794;
srom_1(24475) <= 390072;
srom_1(24476) <= 581857;
srom_1(24477) <= 810252;
srom_1(24478) <= 1074183;
srom_1(24479) <= 1372415;
srom_1(24480) <= 1703547;
srom_1(24481) <= 2066029;
srom_1(24482) <= 2458159;
srom_1(24483) <= 2878099;
srom_1(24484) <= 3323880;
srom_1(24485) <= 3793410;
srom_1(24486) <= 4284490;
srom_1(24487) <= 4794815;
srom_1(24488) <= 5321992;
srom_1(24489) <= 5863550;
srom_1(24490) <= 6416949;
srom_1(24491) <= 6979593;
srom_1(24492) <= 7548845;
srom_1(24493) <= 8122035;
srom_1(24494) <= 8696475;
srom_1(24495) <= 9269471;
srom_1(24496) <= 9838336;
srom_1(24497) <= 10400404;
srom_1(24498) <= 10953037;
srom_1(24499) <= 11493645;
srom_1(24500) <= 12019692;
srom_1(24501) <= 12528711;
srom_1(24502) <= 13018317;
srom_1(24503) <= 13486212;
srom_1(24504) <= 13930202;
srom_1(24505) <= 14348206;
srom_1(24506) <= 14738264;
srom_1(24507) <= 15098546;
srom_1(24508) <= 15427362;
srom_1(24509) <= 15723172;
srom_1(24510) <= 15984587;
srom_1(24511) <= 16210382;
srom_1(24512) <= 16399498;
srom_1(24513) <= 16551048;
srom_1(24514) <= 16664322;
srom_1(24515) <= 16738788;
srom_1(24516) <= 16774097;
srom_1(24517) <= 16770084;
srom_1(24518) <= 16726767;
srom_1(24519) <= 16644349;
srom_1(24520) <= 16523218;
srom_1(24521) <= 16363940;
srom_1(24522) <= 16167264;
srom_1(24523) <= 15934111;
srom_1(24524) <= 15665574;
srom_1(24525) <= 15362913;
srom_1(24526) <= 15027547;
srom_1(24527) <= 14661049;
srom_1(24528) <= 14265137;
srom_1(24529) <= 13841668;
srom_1(24530) <= 13392628;
srom_1(24531) <= 12920122;
srom_1(24532) <= 12426367;
srom_1(24533) <= 11913677;
srom_1(24534) <= 11384457;
srom_1(24535) <= 10841188;
srom_1(24536) <= 10286418;
srom_1(24537) <= 9722749;
srom_1(24538) <= 9152823;
srom_1(24539) <= 8579314;
srom_1(24540) <= 8004910;
srom_1(24541) <= 7432306;
srom_1(24542) <= 6864186;
srom_1(24543) <= 6303215;
srom_1(24544) <= 5752023;
srom_1(24545) <= 5213194;
srom_1(24546) <= 4689257;
srom_1(24547) <= 4182666;
srom_1(24548) <= 3695799;
srom_1(24549) <= 3230938;
srom_1(24550) <= 2790263;
srom_1(24551) <= 2375841;
srom_1(24552) <= 1989615;
srom_1(24553) <= 1633395;
srom_1(24554) <= 1308854;
srom_1(24555) <= 1017511;
srom_1(24556) <= 760734;
srom_1(24557) <= 539727;
srom_1(24558) <= 355526;
srom_1(24559) <= 208995;
srom_1(24560) <= 100821;
srom_1(24561) <= 31511;
srom_1(24562) <= 1391;
srom_1(24563) <= 10601;
srom_1(24564) <= 59098;
srom_1(24565) <= 146655;
srom_1(24566) <= 272862;
srom_1(24567) <= 437126;
srom_1(24568) <= 638677;
srom_1(24569) <= 876571;
srom_1(24570) <= 1149691;
srom_1(24571) <= 1456756;
srom_1(24572) <= 1796328;
srom_1(24573) <= 2166813;
srom_1(24574) <= 2566474;
srom_1(24575) <= 2993437;
srom_1(24576) <= 3445700;
srom_1(24577) <= 3921142;
srom_1(24578) <= 4417533;
srom_1(24579) <= 4932546;
srom_1(24580) <= 5463766;
srom_1(24581) <= 6008701;
srom_1(24582) <= 6564797;
srom_1(24583) <= 7129445;
srom_1(24584) <= 7699997;
srom_1(24585) <= 8273779;
srom_1(24586) <= 8848099;
srom_1(24587) <= 9420265;
srom_1(24588) <= 9987593;
srom_1(24589) <= 10547422;
srom_1(24590) <= 11097128;
srom_1(24591) <= 11634133;
srom_1(24592) <= 12155918;
srom_1(24593) <= 12660038;
srom_1(24594) <= 13144127;
srom_1(24595) <= 13605916;
srom_1(24596) <= 14043239;
srom_1(24597) <= 14454045;
srom_1(24598) <= 14836409;
srom_1(24599) <= 15188536;
srom_1(24600) <= 15508777;
srom_1(24601) <= 15795628;
srom_1(24602) <= 16047746;
srom_1(24603) <= 16263947;
srom_1(24604) <= 16443218;
srom_1(24605) <= 16584718;
srom_1(24606) <= 16687784;
srom_1(24607) <= 16751932;
srom_1(24608) <= 16776861;
srom_1(24609) <= 16762455;
srom_1(24610) <= 16708782;
srom_1(24611) <= 16616092;
srom_1(24612) <= 16484820;
srom_1(24613) <= 16315583;
srom_1(24614) <= 16109173;
srom_1(24615) <= 15866559;
srom_1(24616) <= 15588878;
srom_1(24617) <= 15277433;
srom_1(24618) <= 14933684;
srom_1(24619) <= 14559242;
srom_1(24620) <= 14155865;
srom_1(24621) <= 13725442;
srom_1(24622) <= 13269994;
srom_1(24623) <= 12791654;
srom_1(24624) <= 12292668;
srom_1(24625) <= 11775374;
srom_1(24626) <= 11242198;
srom_1(24627) <= 10695641;
srom_1(24628) <= 10138265;
srom_1(24629) <= 9572685;
srom_1(24630) <= 9001552;
srom_1(24631) <= 8427545;
srom_1(24632) <= 7853355;
srom_1(24633) <= 7281675;
srom_1(24634) <= 6715186;
srom_1(24635) <= 6156544;
srom_1(24636) <= 5608369;
srom_1(24637) <= 5073231;
srom_1(24638) <= 4553641;
srom_1(24639) <= 4052034;
srom_1(24640) <= 3570762;
srom_1(24641) <= 3112083;
srom_1(24642) <= 2678148;
srom_1(24643) <= 2270991;
srom_1(24644) <= 1892521;
srom_1(24645) <= 1544514;
srom_1(24646) <= 1228601;
srom_1(24647) <= 946264;
srom_1(24648) <= 698827;
srom_1(24649) <= 487449;
srom_1(24650) <= 313123;
srom_1(24651) <= 176666;
srom_1(24652) <= 78717;
srom_1(24653) <= 19736;
srom_1(24654) <= 0;
srom_1(24655) <= 19600;
srom_1(24656) <= 78446;
srom_1(24657) <= 176261;
srom_1(24658) <= 312586;
srom_1(24659) <= 486783;
srom_1(24660) <= 698034;
srom_1(24661) <= 945349;
srom_1(24662) <= 1227568;
srom_1(24663) <= 1543367;
srom_1(24664) <= 1891266;
srom_1(24665) <= 2269634;
srom_1(24666) <= 2676695;
srom_1(24667) <= 3110541;
srom_1(24668) <= 3569139;
srom_1(24669) <= 4050336;
srom_1(24670) <= 4551877;
srom_1(24671) <= 5071409;
srom_1(24672) <= 5606497;
srom_1(24673) <= 6154632;
srom_1(24674) <= 6713242;
srom_1(24675) <= 7279708;
srom_1(24676) <= 7851375;
srom_1(24677) <= 8425561;
srom_1(24678) <= 8999573;
srom_1(24679) <= 9570721;
srom_1(24680) <= 10136325;
srom_1(24681) <= 10693734;
srom_1(24682) <= 11240333;
srom_1(24683) <= 11773559;
srom_1(24684) <= 12290912;
srom_1(24685) <= 12789966;
srom_1(24686) <= 13268380;
srom_1(24687) <= 13723912;
srom_1(24688) <= 14154424;
srom_1(24689) <= 14557898;
srom_1(24690) <= 14932443;
srom_1(24691) <= 15276301;
srom_1(24692) <= 15587860;
srom_1(24693) <= 15865660;
srom_1(24694) <= 16108397;
srom_1(24695) <= 16314934;
srom_1(24696) <= 16484301;
srom_1(24697) <= 16615704;
srom_1(24698) <= 16708528;
srom_1(24699) <= 16762337;
srom_1(24700) <= 16776879;
srom_1(24701) <= 16752085;
srom_1(24702) <= 16688072;
srom_1(24703) <= 16585140;
srom_1(24704) <= 16443772;
srom_1(24705) <= 16264630;
srom_1(24706) <= 16048555;
srom_1(24707) <= 15796559;
srom_1(24708) <= 15509826;
srom_1(24709) <= 15189698;
srom_1(24710) <= 14837678;
srom_1(24711) <= 14455415;
srom_1(24712) <= 14044704;
srom_1(24713) <= 13607469;
srom_1(24714) <= 13145761;
srom_1(24715) <= 12661745;
srom_1(24716) <= 12157691;
srom_1(24717) <= 11635962;
srom_1(24718) <= 11099006;
srom_1(24719) <= 10549339;
srom_1(24720) <= 9989540;
srom_1(24721) <= 9422234;
srom_1(24722) <= 8850080;
srom_1(24723) <= 8275763;
srom_1(24724) <= 7701974;
srom_1(24725) <= 7131406;
srom_1(24726) <= 6566733;
srom_1(24727) <= 6010604;
srom_1(24728) <= 5465625;
srom_1(24729) <= 4934354;
srom_1(24730) <= 4419281;
srom_1(24731) <= 3922821;
srom_1(24732) <= 3447303;
srom_1(24733) <= 2994956;
srom_1(24734) <= 2567902;
srom_1(24735) <= 2168144;
srom_1(24736) <= 1797555;
srom_1(24737) <= 1457874;
srom_1(24738) <= 1150693;
srom_1(24739) <= 877454;
srom_1(24740) <= 639437;
srom_1(24741) <= 437758;
srom_1(24742) <= 273364;
srom_1(24743) <= 147025;
srom_1(24744) <= 59333;
srom_1(24745) <= 10701;
srom_1(24746) <= 1355;
srom_1(24747) <= 31340;
srom_1(24748) <= 100515;
srom_1(24749) <= 208555;
srom_1(24750) <= 354955;
srom_1(24751) <= 539028;
srom_1(24752) <= 759909;
srom_1(24753) <= 1016564;
srom_1(24754) <= 1307790;
srom_1(24755) <= 1632220;
srom_1(24756) <= 1988332;
srom_1(24757) <= 2374458;
srom_1(24758) <= 2788786;
srom_1(24759) <= 3229374;
srom_1(24760) <= 3694155;
srom_1(24761) <= 4180950;
srom_1(24762) <= 4687476;
srom_1(24763) <= 5211358;
srom_1(24764) <= 5750139;
srom_1(24765) <= 6301293;
srom_1(24766) <= 6862235;
srom_1(24767) <= 7430335;
srom_1(24768) <= 8002929;
srom_1(24769) <= 8577330;
srom_1(24770) <= 9150847;
srom_1(24771) <= 9720790;
srom_1(24772) <= 10284486;
srom_1(24773) <= 10839291;
srom_1(24774) <= 11382604;
srom_1(24775) <= 11911877;
srom_1(24776) <= 12424628;
srom_1(24777) <= 12918453;
srom_1(24778) <= 13391036;
srom_1(24779) <= 13840161;
srom_1(24780) <= 14263721;
srom_1(24781) <= 14659732;
srom_1(24782) <= 15026334;
srom_1(24783) <= 15361810;
srom_1(24784) <= 15664587;
srom_1(24785) <= 15933244;
srom_1(24786) <= 16166521;
srom_1(24787) <= 16363325;
srom_1(24788) <= 16522733;
srom_1(24789) <= 16643997;
srom_1(24790) <= 16726549;
srom_1(24791) <= 16770002;
srom_1(24792) <= 16774151;
srom_1(24793) <= 16738977;
srom_1(24794) <= 16664646;
srom_1(24795) <= 16551505;
srom_1(24796) <= 16400086;
srom_1(24797) <= 16211099;
srom_1(24798) <= 15985428;
srom_1(24799) <= 15724134;
srom_1(24800) <= 15428441;
srom_1(24801) <= 15099736;
srom_1(24802) <= 14739560;
srom_1(24803) <= 14349602;
srom_1(24804) <= 13931691;
srom_1(24805) <= 13487787;
srom_1(24806) <= 13019971;
srom_1(24807) <= 12530437;
srom_1(24808) <= 12021480;
srom_1(24809) <= 11495487;
srom_1(24810) <= 10954926;
srom_1(24811) <= 10402329;
srom_1(24812) <= 9840290;
srom_1(24813) <= 9271444;
srom_1(24814) <= 8698457;
srom_1(24815) <= 8124018;
srom_1(24816) <= 7550819;
srom_1(24817) <= 6981549;
srom_1(24818) <= 6418877;
srom_1(24819) <= 5865442;
srom_1(24820) <= 5323839;
srom_1(24821) <= 4796607;
srom_1(24822) <= 4286220;
srom_1(24823) <= 3795070;
srom_1(24824) <= 3325461;
srom_1(24825) <= 2879595;
srom_1(24826) <= 2459562;
srom_1(24827) <= 2067333;
srom_1(24828) <= 1704746;
srom_1(24829) <= 1373502;
srom_1(24830) <= 1075155;
srom_1(24831) <= 811102;
srom_1(24832) <= 582584;
srom_1(24833) <= 390670;
srom_1(24834) <= 236261;
srom_1(24835) <= 120082;
srom_1(24836) <= 42677;
srom_1(24837) <= 4408;
srom_1(24838) <= 5456;
srom_1(24839) <= 45815;
srom_1(24840) <= 125297;
srom_1(24841) <= 243528;
srom_1(24842) <= 399954;
srom_1(24843) <= 593842;
srom_1(24844) <= 824282;
srom_1(24845) <= 1090193;
srom_1(24846) <= 1390330;
srom_1(24847) <= 1723284;
srom_1(24848) <= 2087493;
srom_1(24849) <= 2481251;
srom_1(24850) <= 2902711;
srom_1(24851) <= 3349896;
srom_1(24852) <= 3820709;
srom_1(24853) <= 4312942;
srom_1(24854) <= 4824288;
srom_1(24855) <= 5352347;
srom_1(24856) <= 5894645;
srom_1(24857) <= 6448639;
srom_1(24858) <= 7011729;
srom_1(24859) <= 7581276;
srom_1(24860) <= 8154608;
srom_1(24861) <= 8729038;
srom_1(24862) <= 9301872;
srom_1(24863) <= 9870423;
srom_1(24864) <= 10432025;
srom_1(24865) <= 10984045;
srom_1(24866) <= 11523894;
srom_1(24867) <= 12049041;
srom_1(24868) <= 12557022;
srom_1(24869) <= 13045457;
srom_1(24870) <= 13512054;
srom_1(24871) <= 13954625;
srom_1(24872) <= 14371095;
srom_1(24873) <= 14759512;
srom_1(24874) <= 15118053;
srom_1(24875) <= 15445037;
srom_1(24876) <= 15738931;
srom_1(24877) <= 15998357;
srom_1(24878) <= 16222099;
srom_1(24879) <= 16409106;
srom_1(24880) <= 16558503;
srom_1(24881) <= 16669588;
srom_1(24882) <= 16741840;
srom_1(24883) <= 16774922;
srom_1(24884) <= 16768677;
srom_1(24885) <= 16723135;
srom_1(24886) <= 16638510;
srom_1(24887) <= 16515198;
srom_1(24888) <= 16353778;
srom_1(24889) <= 16155006;
srom_1(24890) <= 15919815;
srom_1(24891) <= 15649308;
srom_1(24892) <= 15344752;
srom_1(24893) <= 15007577;
srom_1(24894) <= 14639363;
srom_1(24895) <= 14241838;
srom_1(24896) <= 13816864;
srom_1(24897) <= 13366436;
srom_1(24898) <= 12892664;
srom_1(24899) <= 12397772;
srom_1(24900) <= 11884079;
srom_1(24901) <= 11353995;
srom_1(24902) <= 10810005;
srom_1(24903) <= 10254661;
srom_1(24904) <= 9690566;
srom_1(24905) <= 9120365;
srom_1(24906) <= 8546733;
srom_1(24907) <= 7972359;
srom_1(24908) <= 7399938;
srom_1(24909) <= 6832152;
srom_1(24910) <= 6271666;
srom_1(24911) <= 5721106;
srom_1(24912) <= 5183055;
srom_1(24913) <= 4660037;
srom_1(24914) <= 4154502;
srom_1(24915) <= 3668823;
srom_1(24916) <= 3205277;
srom_1(24917) <= 2766037;
srom_1(24918) <= 2353163;
srom_1(24919) <= 1968591;
srom_1(24920) <= 1614126;
srom_1(24921) <= 1291427;
srom_1(24922) <= 1002011;
srom_1(24923) <= 747232;
srom_1(24924) <= 528286;
srom_1(24925) <= 346200;
srom_1(24926) <= 201828;
srom_1(24927) <= 95846;
srom_1(24928) <= 28752;
srom_1(24929) <= 861;
srom_1(24930) <= 12302;
srom_1(24931) <= 63022;
srom_1(24932) <= 152784;
srom_1(24933) <= 281167;
srom_1(24934) <= 447568;
srom_1(24935) <= 651208;
srom_1(24936) <= 891131;
srom_1(24937) <= 1166212;
srom_1(24938) <= 1475161;
srom_1(24939) <= 1816530;
srom_1(24940) <= 2188718;
srom_1(24941) <= 2589979;
srom_1(24942) <= 3018431;
srom_1(24943) <= 3472067;
srom_1(24944) <= 3948757;
srom_1(24945) <= 4446268;
srom_1(24946) <= 4962266;
srom_1(24947) <= 5494331;
srom_1(24948) <= 6039968;
srom_1(24949) <= 6596619;
srom_1(24950) <= 7161673;
srom_1(24951) <= 7732480;
srom_1(24952) <= 8306365;
srom_1(24953) <= 8880635;
srom_1(24954) <= 9452597;
srom_1(24955) <= 10019571;
srom_1(24956) <= 10578896;
srom_1(24957) <= 11127950;
srom_1(24958) <= 11664158;
srom_1(24959) <= 12185007;
srom_1(24960) <= 12688052;
srom_1(24961) <= 13170936;
srom_1(24962) <= 13631394;
srom_1(24963) <= 14067267;
srom_1(24964) <= 14476511;
srom_1(24965) <= 14857206;
srom_1(24966) <= 15207568;
srom_1(24967) <= 15525953;
srom_1(24968) <= 15810869;
srom_1(24969) <= 16060980;
srom_1(24970) <= 16275112;
srom_1(24971) <= 16452261;
srom_1(24972) <= 16591597;
srom_1(24973) <= 16692467;
srom_1(24974) <= 16754397;
srom_1(24975) <= 16777097;
srom_1(24976) <= 16760460;
srom_1(24977) <= 16704565;
srom_1(24978) <= 16609673;
srom_1(24979) <= 16476230;
srom_1(24980) <= 16304862;
srom_1(24981) <= 16096371;
srom_1(24982) <= 15851736;
srom_1(24983) <= 15572104;
srom_1(24984) <= 15258786;
srom_1(24985) <= 14913251;
srom_1(24986) <= 14537120;
srom_1(24987) <= 14132157;
srom_1(24988) <= 13700260;
srom_1(24989) <= 13243455;
srom_1(24990) <= 12763883;
srom_1(24991) <= 12263795;
srom_1(24992) <= 11745535;
srom_1(24993) <= 11211532;
srom_1(24994) <= 10664292;
srom_1(24995) <= 10106381;
srom_1(24996) <= 9540414;
srom_1(24997) <= 8969047;
srom_1(24998) <= 8394957;
srom_1(24999) <= 7820837;
srom_1(25000) <= 7249380;
srom_1(25001) <= 6683266;
srom_1(25002) <= 6125148;
srom_1(25003) <= 5577644;
srom_1(25004) <= 5043322;
srom_1(25005) <= 4524687;
srom_1(25006) <= 4024171;
srom_1(25007) <= 3544122;
srom_1(25008) <= 3086790;
srom_1(25009) <= 2654320;
srom_1(25010) <= 2248740;
srom_1(25011) <= 1871952;
srom_1(25012) <= 1525723;
srom_1(25013) <= 1211676;
srom_1(25014) <= 931285;
srom_1(25015) <= 685863;
srom_1(25016) <= 476562;
srom_1(25017) <= 304364;
srom_1(25018) <= 170075;
srom_1(25019) <= 74326;
srom_1(25020) <= 17565;
srom_1(25021) <= 59;
srom_1(25022) <= 21890;
srom_1(25023) <= 82955;
srom_1(25024) <= 182968;
srom_1(25025) <= 321460;
srom_1(25026) <= 497782;
srom_1(25027) <= 711107;
srom_1(25028) <= 960434;
srom_1(25029) <= 1244595;
srom_1(25030) <= 1562256;
srom_1(25031) <= 1911928;
srom_1(25032) <= 2291971;
srom_1(25033) <= 2700604;
srom_1(25034) <= 3135910;
srom_1(25035) <= 3595848;
srom_1(25036) <= 4078260;
srom_1(25037) <= 4580885;
srom_1(25038) <= 5101366;
srom_1(25039) <= 5637262;
srom_1(25040) <= 6186059;
srom_1(25041) <= 6745186;
srom_1(25042) <= 7312019;
srom_1(25043) <= 7883900;
srom_1(25044) <= 8458148;
srom_1(25045) <= 9032070;
srom_1(25046) <= 9602975;
srom_1(25047) <= 10168185;
srom_1(25048) <= 10725049;
srom_1(25049) <= 11270958;
srom_1(25050) <= 11803350;
srom_1(25051) <= 12319730;
srom_1(25052) <= 12817674;
srom_1(25053) <= 13294850;
srom_1(25054) <= 13749018;
srom_1(25055) <= 14178050;
srom_1(25056) <= 14579933;
srom_1(25057) <= 14952783;
srom_1(25058) <= 15294851;
srom_1(25059) <= 15604533;
srom_1(25060) <= 15880377;
srom_1(25061) <= 16121090;
srom_1(25062) <= 16325542;
srom_1(25063) <= 16492776;
srom_1(25064) <= 16622006;
srom_1(25065) <= 16712627;
srom_1(25066) <= 16764214;
srom_1(25067) <= 16776525;
srom_1(25068) <= 16749502;
srom_1(25069) <= 16683272;
srom_1(25070) <= 16578145;
srom_1(25071) <= 16434615;
srom_1(25072) <= 16253354;
srom_1(25073) <= 16035212;
srom_1(25074) <= 15781214;
srom_1(25075) <= 15492548;
srom_1(25076) <= 15170570;
srom_1(25077) <= 14816789;
srom_1(25078) <= 14432864;
srom_1(25079) <= 14020595;
srom_1(25080) <= 13581916;
srom_1(25081) <= 13118884;
srom_1(25082) <= 12633670;
srom_1(25083) <= 12128549;
srom_1(25084) <= 11605891;
srom_1(25085) <= 11068145;
srom_1(25086) <= 10517834;
srom_1(25087) <= 9957539;
srom_1(25088) <= 9389886;
srom_1(25089) <= 8817538;
srom_1(25090) <= 8243179;
srom_1(25091) <= 7669501;
srom_1(25092) <= 7099196;
srom_1(25093) <= 6534937;
srom_1(25094) <= 5979371;
srom_1(25095) <= 5435102;
srom_1(25096) <= 4904683;
srom_1(25097) <= 4390602;
srom_1(25098) <= 3895269;
srom_1(25099) <= 3421006;
srom_1(25100) <= 2970038;
srom_1(25101) <= 2544480;
srom_1(25102) <= 2146327;
srom_1(25103) <= 1777446;
srom_1(25104) <= 1439567;
srom_1(25105) <= 1134275;
srom_1(25106) <= 863000;
srom_1(25107) <= 627016;
srom_1(25108) <= 427429;
srom_1(25109) <= 265174;
srom_1(25110) <= 141012;
srom_1(25111) <= 55527;
srom_1(25112) <= 9118;
srom_1(25113) <= 2004;
srom_1(25114) <= 34217;
srom_1(25115) <= 105607;
srom_1(25116) <= 215838;
srom_1(25117) <= 364395;
srom_1(25118) <= 550580;
srom_1(25119) <= 773520;
srom_1(25120) <= 1032170;
srom_1(25121) <= 1325316;
srom_1(25122) <= 1651585;
srom_1(25123) <= 2009446;
srom_1(25124) <= 2397221;
srom_1(25125) <= 2813092;
srom_1(25126) <= 3255108;
srom_1(25127) <= 3721198;
srom_1(25128) <= 4209174;
srom_1(25129) <= 4716749;
srom_1(25130) <= 5241542;
srom_1(25131) <= 5781093;
srom_1(25132) <= 6332872;
srom_1(25133) <= 6894291;
srom_1(25134) <= 7462717;
srom_1(25135) <= 8035485;
srom_1(25136) <= 8609909;
srom_1(25137) <= 9183295;
srom_1(25138) <= 9752954;
srom_1(25139) <= 10316216;
srom_1(25140) <= 10870438;
srom_1(25141) <= 11413022;
srom_1(25142) <= 11941424;
srom_1(25143) <= 12453165;
srom_1(25144) <= 12945847;
srom_1(25145) <= 13417157;
srom_1(25146) <= 13864888;
srom_1(25147) <= 14286937;
srom_1(25148) <= 14681328;
srom_1(25149) <= 15046210;
srom_1(25150) <= 15379872;
srom_1(25151) <= 15680750;
srom_1(25152) <= 15947432;
srom_1(25153) <= 16178669;
srom_1(25154) <= 16373375;
srom_1(25155) <= 16530638;
srom_1(25156) <= 16649720;
srom_1(25157) <= 16730063;
srom_1(25158) <= 16771289;
srom_1(25159) <= 16773207;
srom_1(25160) <= 16735806;
srom_1(25161) <= 16659263;
srom_1(25162) <= 16543935;
srom_1(25163) <= 16390365;
srom_1(25164) <= 16199271;
srom_1(25165) <= 15971550;
srom_1(25166) <= 15708271;
srom_1(25167) <= 15410667;
srom_1(25168) <= 15080134;
srom_1(25169) <= 14718222;
srom_1(25170) <= 14326629;
srom_1(25171) <= 13907190;
srom_1(25172) <= 13461873;
srom_1(25173) <= 12992765;
srom_1(25174) <= 12502067;
srom_1(25175) <= 11992079;
srom_1(25176) <= 11465194;
srom_1(25177) <= 10923881;
srom_1(25178) <= 10370679;
srom_1(25179) <= 9808183;
srom_1(25180) <= 9239030;
srom_1(25181) <= 8665889;
srom_1(25182) <= 8091448;
srom_1(25183) <= 7518401;
srom_1(25184) <= 6949434;
srom_1(25185) <= 6387215;
srom_1(25186) <= 5834382;
srom_1(25187) <= 5293527;
srom_1(25188) <= 4767185;
srom_1(25189) <= 4257826;
srom_1(25190) <= 3767837;
srom_1(25191) <= 3299517;
srom_1(25192) <= 2855061;
srom_1(25193) <= 2436554;
srom_1(25194) <= 2045958;
srom_1(25195) <= 1685105;
srom_1(25196) <= 1355687;
srom_1(25197) <= 1059248;
srom_1(25198) <= 797180;
srom_1(25199) <= 570710;
srom_1(25200) <= 380901;
srom_1(25201) <= 228643;
srom_1(25202) <= 114650;
srom_1(25203) <= 39457;
srom_1(25204) <= 3415;
srom_1(25205) <= 6694;
srom_1(25206) <= 49279;
srom_1(25207) <= 130971;
srom_1(25208) <= 251384;
srom_1(25209) <= 409957;
srom_1(25210) <= 605943;
srom_1(25211) <= 838426;
srom_1(25212) <= 1106314;
srom_1(25213) <= 1408351;
srom_1(25214) <= 1743120;
srom_1(25215) <= 2109053;
srom_1(25216) <= 2504433;
srom_1(25217) <= 2927405;
srom_1(25218) <= 3375988;
srom_1(25219) <= 3848076;
srom_1(25220) <= 4341456;
srom_1(25221) <= 4853814;
srom_1(25222) <= 5382749;
srom_1(25223) <= 5925779;
srom_1(25224) <= 6480357;
srom_1(25225) <= 7043885;
srom_1(25226) <= 7613718;
srom_1(25227) <= 8187185;
srom_1(25228) <= 8761597;
srom_1(25229) <= 9334259;
srom_1(25230) <= 9902487;
srom_1(25231) <= 10463616;
srom_1(25232) <= 11015014;
srom_1(25233) <= 11554097;
srom_1(25234) <= 12078335;
srom_1(25235) <= 12585271;
srom_1(25236) <= 13072527;
srom_1(25237) <= 13537818;
srom_1(25238) <= 13978964;
srom_1(25239) <= 14393894;
srom_1(25240) <= 14780663;
srom_1(25241) <= 15137458;
srom_1(25242) <= 15462605;
srom_1(25243) <= 15754580;
srom_1(25244) <= 16012013;
srom_1(25245) <= 16233697;
srom_1(25246) <= 16418593;
srom_1(25247) <= 16565834;
srom_1(25248) <= 16674729;
srom_1(25249) <= 16744767;
srom_1(25250) <= 16775620;
srom_1(25251) <= 16767144;
srom_1(25252) <= 16719378;
srom_1(25253) <= 16632546;
srom_1(25254) <= 16507056;
srom_1(25255) <= 16343495;
srom_1(25256) <= 16142631;
srom_1(25257) <= 15905406;
srom_1(25258) <= 15632932;
srom_1(25259) <= 15326487;
srom_1(25260) <= 14987507;
srom_1(25261) <= 14617583;
srom_1(25262) <= 14218450;
srom_1(25263) <= 13791978;
srom_1(25264) <= 13340168;
srom_1(25265) <= 12865138;
srom_1(25266) <= 12369117;
srom_1(25267) <= 11854429;
srom_1(25268) <= 11323489;
srom_1(25269) <= 10778786;
srom_1(25270) <= 10222875;
srom_1(25271) <= 9658363;
srom_1(25272) <= 9087896;
srom_1(25273) <= 8514150;
srom_1(25274) <= 7939815;
srom_1(25275) <= 7367585;
srom_1(25276) <= 6800142;
srom_1(25277) <= 6240149;
srom_1(25278) <= 5690230;
srom_1(25279) <= 5152965;
srom_1(25280) <= 4630873;
srom_1(25281) <= 4126402;
srom_1(25282) <= 3641919;
srom_1(25283) <= 3179694;
srom_1(25284) <= 2741895;
srom_1(25285) <= 2330576;
srom_1(25286) <= 1947665;
srom_1(25287) <= 1594958;
srom_1(25288) <= 1274108;
srom_1(25289) <= 986621;
srom_1(25290) <= 733845;
srom_1(25291) <= 516964;
srom_1(25292) <= 336996;
srom_1(25293) <= 194784;
srom_1(25294) <= 90997;
srom_1(25295) <= 26120;
srom_1(25296) <= 457;
srom_1(25297) <= 14129;
srom_1(25298) <= 67072;
srom_1(25299) <= 159038;
srom_1(25300) <= 289595;
srom_1(25301) <= 458130;
srom_1(25302) <= 663855;
srom_1(25303) <= 905804;
srom_1(25304) <= 1182842;
srom_1(25305) <= 1493670;
srom_1(25306) <= 1836831;
srom_1(25307) <= 2210716;
srom_1(25308) <= 2613571;
srom_1(25309) <= 3043507;
srom_1(25310) <= 3498508;
srom_1(25311) <= 3976440;
srom_1(25312) <= 4475063;
srom_1(25313) <= 4992037;
srom_1(25314) <= 5524939;
srom_1(25315) <= 6071270;
srom_1(25316) <= 6628468;
srom_1(25317) <= 7193919;
srom_1(25318) <= 7764973;
srom_1(25319) <= 8338952;
srom_1(25320) <= 8913163;
srom_1(25321) <= 9484914;
srom_1(25322) <= 10051524;
srom_1(25323) <= 10610337;
srom_1(25324) <= 11158731;
srom_1(25325) <= 11694134;
srom_1(25326) <= 12214037;
srom_1(25327) <= 12716002;
srom_1(25328) <= 13197673;
srom_1(25329) <= 13656794;
srom_1(25330) <= 14091210;
srom_1(25331) <= 14498884;
srom_1(25332) <= 14877906;
srom_1(25333) <= 15226496;
srom_1(25334) <= 15543022;
srom_1(25335) <= 15825998;
srom_1(25336) <= 16074097;
srom_1(25337) <= 16286157;
srom_1(25338) <= 16461182;
srom_1(25339) <= 16598353;
srom_1(25340) <= 16697025;
srom_1(25341) <= 16756735;
srom_1(25342) <= 16777205;
srom_1(25343) <= 16758338;
srom_1(25344) <= 16700222;
srom_1(25345) <= 16603131;
srom_1(25346) <= 16467518;
srom_1(25347) <= 16294021;
srom_1(25348) <= 16083453;
srom_1(25349) <= 15836800;
srom_1(25350) <= 15555221;
srom_1(25351) <= 15240035;
srom_1(25352) <= 14892720;
srom_1(25353) <= 14514905;
srom_1(25354) <= 14108362;
srom_1(25355) <= 13674997;
srom_1(25356) <= 13216842;
srom_1(25357) <= 12736046;
srom_1(25358) <= 12234864;
srom_1(25359) <= 11715645;
srom_1(25360) <= 11180824;
srom_1(25361) <= 10632910;
srom_1(25362) <= 10074471;
srom_1(25363) <= 9508127;
srom_1(25364) <= 8936533;
srom_1(25365) <= 8362369;
srom_1(25366) <= 7788329;
srom_1(25367) <= 7217103;
srom_1(25368) <= 6651371;
srom_1(25369) <= 6093786;
srom_1(25370) <= 5546961;
srom_1(25371) <= 5013463;
srom_1(25372) <= 4495791;
srom_1(25373) <= 3996374;
srom_1(25374) <= 3517554;
srom_1(25375) <= 3061576;
srom_1(25376) <= 2630578;
srom_1(25377) <= 2226582;
srom_1(25378) <= 1851481;
srom_1(25379) <= 1507035;
srom_1(25380) <= 1194859;
srom_1(25381) <= 916418;
srom_1(25382) <= 673016;
srom_1(25383) <= 465794;
srom_1(25384) <= 295726;
srom_1(25385) <= 163608;
srom_1(25386) <= 70060;
srom_1(25387) <= 15520;
srom_1(25388) <= 245;
srom_1(25389) <= 24306;
srom_1(25390) <= 87589;
srom_1(25391) <= 189799;
srom_1(25392) <= 330456;
srom_1(25393) <= 508901;
srom_1(25394) <= 724296;
srom_1(25395) <= 975631;
srom_1(25396) <= 1261729;
srom_1(25397) <= 1581247;
srom_1(25398) <= 1932687;
srom_1(25399) <= 2314401;
srom_1(25400) <= 2724599;
srom_1(25401) <= 3161358;
srom_1(25402) <= 3622629;
srom_1(25403) <= 4106249;
srom_1(25404) <= 4609951;
srom_1(25405) <= 5131372;
srom_1(25406) <= 5668067;
srom_1(25407) <= 6217520;
srom_1(25408) <= 6777154;
srom_1(25409) <= 7344345;
srom_1(25410) <= 7916432;
srom_1(25411) <= 8490734;
srom_1(25412) <= 9064557;
srom_1(25413) <= 9635210;
srom_1(25414) <= 10200017;
srom_1(25415) <= 10756330;
srom_1(25416) <= 11301540;
srom_1(25417) <= 11833090;
srom_1(25418) <= 12348488;
srom_1(25419) <= 12845316;
srom_1(25420) <= 13321246;
srom_1(25421) <= 13774044;
srom_1(25422) <= 14201589;
srom_1(25423) <= 14601874;
srom_1(25424) <= 14973023;
srom_1(25425) <= 15313296;
srom_1(25426) <= 15621096;
srom_1(25427) <= 15894981;
srom_1(25428) <= 16133666;
srom_1(25429) <= 16336032;
srom_1(25430) <= 16501129;
srom_1(25431) <= 16628184;
srom_1(25432) <= 16716601;
srom_1(25433) <= 16765964;
srom_1(25434) <= 16776044;
srom_1(25435) <= 16746792;
srom_1(25436) <= 16678346;
srom_1(25437) <= 16571026;
srom_1(25438) <= 16425336;
srom_1(25439) <= 16241959;
srom_1(25440) <= 16021755;
srom_1(25441) <= 15765756;
srom_1(25442) <= 15475164;
srom_1(25443) <= 15151340;
srom_1(25444) <= 14795803;
srom_1(25445) <= 14410221;
srom_1(25446) <= 13996402;
srom_1(25447) <= 13556285;
srom_1(25448) <= 13091936;
srom_1(25449) <= 12605531;
srom_1(25450) <= 12099351;
srom_1(25451) <= 11575771;
srom_1(25452) <= 11037244;
srom_1(25453) <= 10486298;
srom_1(25454) <= 9925514;
srom_1(25455) <= 9357524;
srom_1(25456) <= 8784990;
srom_1(25457) <= 8210597;
srom_1(25458) <= 7637039;
srom_1(25459) <= 7067005;
srom_1(25460) <= 6503169;
srom_1(25461) <= 5948174;
srom_1(25462) <= 5404623;
srom_1(25463) <= 4875065;
srom_1(25464) <= 4361984;
srom_1(25465) <= 3867784;
srom_1(25466) <= 3394784;
srom_1(25467) <= 2945202;
srom_1(25468) <= 2521146;
srom_1(25469) <= 2124605;
srom_1(25470) <= 1757437;
srom_1(25471) <= 1421366;
srom_1(25472) <= 1117966;
srom_1(25473) <= 848660;
srom_1(25474) <= 614712;
srom_1(25475) <= 417219;
srom_1(25476) <= 257106;
srom_1(25477) <= 135125;
srom_1(25478) <= 51847;
srom_1(25479) <= 7662;
srom_1(25480) <= 2779;
srom_1(25481) <= 37220;
srom_1(25482) <= 110824;
srom_1(25483) <= 223245;
srom_1(25484) <= 373956;
srom_1(25485) <= 562251;
srom_1(25486) <= 787246;
srom_1(25487) <= 1047886;
srom_1(25488) <= 1342950;
srom_1(25489) <= 1671053;
srom_1(25490) <= 2030657;
srom_1(25491) <= 2420075;
srom_1(25492) <= 2837482;
srom_1(25493) <= 3280920;
srom_1(25494) <= 3748310;
srom_1(25495) <= 4237460;
srom_1(25496) <= 4746076;
srom_1(25497) <= 5271773;
srom_1(25498) <= 5812086;
srom_1(25499) <= 6364482;
srom_1(25500) <= 6926369;
srom_1(25501) <= 7495112;
srom_1(25502) <= 8068046;
srom_1(25503) <= 8642483;
srom_1(25504) <= 9215730;
srom_1(25505) <= 9785098;
srom_1(25506) <= 10347917;
srom_1(25507) <= 10901548;
srom_1(25508) <= 11443396;
srom_1(25509) <= 11970918;
srom_1(25510) <= 12481642;
srom_1(25511) <= 12973172;
srom_1(25512) <= 13443203;
srom_1(25513) <= 13889532;
srom_1(25514) <= 14310065;
srom_1(25515) <= 14702830;
srom_1(25516) <= 15065986;
srom_1(25517) <= 15397829;
srom_1(25518) <= 15696803;
srom_1(25519) <= 15961507;
srom_1(25520) <= 16190699;
srom_1(25521) <= 16383304;
srom_1(25522) <= 16538419;
srom_1(25523) <= 16655317;
srom_1(25524) <= 16733450;
srom_1(25525) <= 16772451;
srom_1(25526) <= 16772137;
srom_1(25527) <= 16732509;
srom_1(25528) <= 16653755;
srom_1(25529) <= 16536242;
srom_1(25530) <= 16380522;
srom_1(25531) <= 16187326;
srom_1(25532) <= 15957558;
srom_1(25533) <= 15692297;
srom_1(25534) <= 15392787;
srom_1(25535) <= 15060431;
srom_1(25536) <= 14696789;
srom_1(25537) <= 14303566;
srom_1(25538) <= 13882605;
srom_1(25539) <= 13435882;
srom_1(25540) <= 12965490;
srom_1(25541) <= 12473635;
srom_1(25542) <= 11962624;
srom_1(25543) <= 11434853;
srom_1(25544) <= 10892798;
srom_1(25545) <= 10338999;
srom_1(25546) <= 9776055;
srom_1(25547) <= 9206604;
srom_1(25548) <= 8633317;
srom_1(25549) <= 8058883;
srom_1(25550) <= 7485995;
srom_1(25551) <= 6917340;
srom_1(25552) <= 6355584;
srom_1(25553) <= 5803361;
srom_1(25554) <= 5263262;
srom_1(25555) <= 4737818;
srom_1(25556) <= 4229494;
srom_1(25557) <= 3740674;
srom_1(25558) <= 3273649;
srom_1(25559) <= 2830611;
srom_1(25560) <= 2413635;
srom_1(25561) <= 2024678;
srom_1(25562) <= 1665564;
srom_1(25563) <= 1337977;
srom_1(25564) <= 1043452;
srom_1(25565) <= 783372;
srom_1(25566) <= 558955;
srom_1(25567) <= 371253;
srom_1(25568) <= 221148;
srom_1(25569) <= 109343;
srom_1(25570) <= 36363;
srom_1(25571) <= 2548;
srom_1(25572) <= 8059;
srom_1(25573) <= 52870;
srom_1(25574) <= 136769;
srom_1(25575) <= 259364;
srom_1(25576) <= 420080;
srom_1(25577) <= 618163;
srom_1(25578) <= 852684;
srom_1(25579) <= 1122544;
srom_1(25580) <= 1426477;
srom_1(25581) <= 1763057;
srom_1(25582) <= 2130708;
srom_1(25583) <= 2527703;
srom_1(25584) <= 2952183;
srom_1(25585) <= 3402155;
srom_1(25586) <= 3875511;
srom_1(25587) <= 4370030;
srom_1(25588) <= 4883394;
srom_1(25589) <= 5413195;
srom_1(25590) <= 5956949;
srom_1(25591) <= 6512105;
srom_1(25592) <= 7076061;
srom_1(25593) <= 7646172;
srom_1(25594) <= 8219765;
srom_1(25595) <= 8794149;
srom_1(25596) <= 9366632;
srom_1(25597) <= 9934528;
srom_1(25598) <= 10495175;
srom_1(25599) <= 11045944;
srom_1(25600) <= 11584251;
srom_1(25601) <= 12107573;
srom_1(25602) <= 12613455;
srom_1(25603) <= 13099526;
srom_1(25604) <= 13563506;
srom_1(25605) <= 14003218;
srom_1(25606) <= 14416602;
srom_1(25607) <= 14801718;
srom_1(25608) <= 15156762;
srom_1(25609) <= 15480066;
srom_1(25610) <= 15770117;
srom_1(25611) <= 16025553;
srom_1(25612) <= 16245177;
srom_1(25613) <= 16427959;
srom_1(25614) <= 16573042;
srom_1(25615) <= 16679744;
srom_1(25616) <= 16747567;
srom_1(25617) <= 16776192;
srom_1(25618) <= 16765485;
srom_1(25619) <= 16715495;
srom_1(25620) <= 16626458;
srom_1(25621) <= 16498791;
srom_1(25622) <= 16333092;
srom_1(25623) <= 16130139;
srom_1(25624) <= 15890883;
srom_1(25625) <= 15616447;
srom_1(25626) <= 15308116;
srom_1(25627) <= 14967338;
srom_1(25628) <= 14595710;
srom_1(25629) <= 14194974;
srom_1(25630) <= 13767010;
srom_1(25631) <= 13313826;
srom_1(25632) <= 12837545;
srom_1(25633) <= 12340401;
srom_1(25634) <= 11824727;
srom_1(25635) <= 11292939;
srom_1(25636) <= 10747532;
srom_1(25637) <= 10191062;
srom_1(25638) <= 9626141;
srom_1(25639) <= 9055416;
srom_1(25640) <= 8481565;
srom_1(25641) <= 7907277;
srom_1(25642) <= 7335247;
srom_1(25643) <= 6768156;
srom_1(25644) <= 6208664;
srom_1(25645) <= 5659395;
srom_1(25646) <= 5122924;
srom_1(25647) <= 4601766;
srom_1(25648) <= 4098367;
srom_1(25649) <= 3615086;
srom_1(25650) <= 3154189;
srom_1(25651) <= 2717839;
srom_1(25652) <= 2308080;
srom_1(25653) <= 1926836;
srom_1(25654) <= 1575893;
srom_1(25655) <= 1256897;
srom_1(25656) <= 971344;
srom_1(25657) <= 720573;
srom_1(25658) <= 505760;
srom_1(25659) <= 327913;
srom_1(25660) <= 187864;
srom_1(25661) <= 86273;
srom_1(25662) <= 23613;
srom_1(25663) <= 180;
srom_1(25664) <= 16083;
srom_1(25665) <= 71248;
srom_1(25666) <= 165415;
srom_1(25667) <= 298144;
srom_1(25668) <= 468812;
srom_1(25669) <= 676619;
srom_1(25670) <= 920590;
srom_1(25671) <= 1199581;
srom_1(25672) <= 1512283;
srom_1(25673) <= 1857231;
srom_1(25674) <= 2232807;
srom_1(25675) <= 2637250;
srom_1(25676) <= 3068663;
srom_1(25677) <= 3525023;
srom_1(25678) <= 4004189;
srom_1(25679) <= 4503916;
srom_1(25680) <= 5021860;
srom_1(25681) <= 5555591;
srom_1(25682) <= 6102607;
srom_1(25683) <= 6660343;
srom_1(25684) <= 7226184;
srom_1(25685) <= 7797475;
srom_1(25686) <= 8371539;
srom_1(25687) <= 8945683;
srom_1(25688) <= 9517214;
srom_1(25689) <= 10083453;
srom_1(25690) <= 10641744;
srom_1(25691) <= 11189469;
srom_1(25692) <= 11724061;
srom_1(25693) <= 12243011;
srom_1(25694) <= 12743886;
srom_1(25695) <= 13224338;
srom_1(25696) <= 13682114;
srom_1(25697) <= 14115066;
srom_1(25698) <= 14521166;
srom_1(25699) <= 14898507;
srom_1(25700) <= 15245322;
srom_1(25701) <= 15559983;
srom_1(25702) <= 15841014;
srom_1(25703) <= 16087099;
srom_1(25704) <= 16297084;
srom_1(25705) <= 16469982;
srom_1(25706) <= 16604984;
srom_1(25707) <= 16701457;
srom_1(25708) <= 16758948;
srom_1(25709) <= 16777188;
srom_1(25710) <= 16756090;
srom_1(25711) <= 16695755;
srom_1(25712) <= 16596464;
srom_1(25713) <= 16458684;
srom_1(25714) <= 16283061;
srom_1(25715) <= 16070418;
srom_1(25716) <= 15821752;
srom_1(25717) <= 15538230;
srom_1(25718) <= 15221180;
srom_1(25719) <= 14872091;
srom_1(25720) <= 14492598;
srom_1(25721) <= 14084481;
srom_1(25722) <= 13649655;
srom_1(25723) <= 13190157;
srom_1(25724) <= 12708144;
srom_1(25725) <= 12205874;
srom_1(25726) <= 11685704;
srom_1(25727) <= 11150073;
srom_1(25728) <= 10601493;
srom_1(25729) <= 10042535;
srom_1(25730) <= 9475822;
srom_1(25731) <= 8904010;
srom_1(25732) <= 8329782;
srom_1(25733) <= 7755829;
srom_1(25734) <= 7184844;
srom_1(25735) <= 6619503;
srom_1(25736) <= 6062458;
srom_1(25737) <= 5516322;
srom_1(25738) <= 4983654;
srom_1(25739) <= 4466954;
srom_1(25740) <= 3968644;
srom_1(25741) <= 3491060;
srom_1(25742) <= 3036443;
srom_1(25743) <= 2606923;
srom_1(25744) <= 2204516;
srom_1(25745) <= 1831109;
srom_1(25746) <= 1488451;
srom_1(25747) <= 1178151;
srom_1(25748) <= 901663;
srom_1(25749) <= 660284;
srom_1(25750) <= 455146;
srom_1(25751) <= 287211;
srom_1(25752) <= 157266;
srom_1(25753) <= 65920;
srom_1(25754) <= 13602;
srom_1(25755) <= 558;
srom_1(25756) <= 26848;
srom_1(25757) <= 92349;
srom_1(25758) <= 196754;
srom_1(25759) <= 339574;
srom_1(25760) <= 520138;
srom_1(25761) <= 737600;
srom_1(25762) <= 990940;
srom_1(25763) <= 1278971;
srom_1(25764) <= 1600341;
srom_1(25765) <= 1953544;
srom_1(25766) <= 2336923;
srom_1(25767) <= 2748680;
srom_1(25768) <= 3186885;
srom_1(25769) <= 3649482;
srom_1(25770) <= 4134303;
srom_1(25771) <= 4639074;
srom_1(25772) <= 5161427;
srom_1(25773) <= 5698914;
srom_1(25774) <= 6249014;
srom_1(25775) <= 6809147;
srom_1(25776) <= 7376687;
srom_1(25777) <= 7948972;
srom_1(25778) <= 8523319;
srom_1(25779) <= 9097034;
srom_1(25780) <= 9667426;
srom_1(25781) <= 10231822;
srom_1(25782) <= 10787575;
srom_1(25783) <= 11332078;
srom_1(25784) <= 11862778;
srom_1(25785) <= 12377186;
srom_1(25786) <= 12872891;
srom_1(25787) <= 13347567;
srom_1(25788) <= 13798989;
srom_1(25789) <= 14225040;
srom_1(25790) <= 14623722;
srom_1(25791) <= 14993165;
srom_1(25792) <= 15331637;
srom_1(25793) <= 15637551;
srom_1(25794) <= 15909472;
srom_1(25795) <= 16146125;
srom_1(25796) <= 16346401;
srom_1(25797) <= 16509359;
srom_1(25798) <= 16634237;
srom_1(25799) <= 16720448;
srom_1(25800) <= 16767588;
srom_1(25801) <= 16775437;
srom_1(25802) <= 16743956;
srom_1(25803) <= 16673295;
srom_1(25804) <= 16563783;
srom_1(25805) <= 16415936;
srom_1(25806) <= 16230445;
srom_1(25807) <= 16008182;
srom_1(25808) <= 15750188;
srom_1(25809) <= 15457672;
srom_1(25810) <= 15132008;
srom_1(25811) <= 14774721;
srom_1(25812) <= 14387488;
srom_1(25813) <= 13972124;
srom_1(25814) <= 13530576;
srom_1(25815) <= 13064917;
srom_1(25816) <= 12577328;
srom_1(25817) <= 12070097;
srom_1(25818) <= 11545603;
srom_1(25819) <= 11006304;
srom_1(25820) <= 10454730;
srom_1(25821) <= 9893467;
srom_1(25822) <= 9325147;
srom_1(25823) <= 8752436;
srom_1(25824) <= 8178018;
srom_1(25825) <= 7604588;
srom_1(25826) <= 7034834;
srom_1(25827) <= 6471429;
srom_1(25828) <= 5917014;
srom_1(25829) <= 5374189;
srom_1(25830) <= 4845500;
srom_1(25831) <= 4333426;
srom_1(25832) <= 3840368;
srom_1(25833) <= 3368638;
srom_1(25834) <= 2920448;
srom_1(25835) <= 2497901;
srom_1(25836) <= 2102977;
srom_1(25837) <= 1737528;
srom_1(25838) <= 1403269;
srom_1(25839) <= 1101766;
srom_1(25840) <= 834434;
srom_1(25841) <= 602526;
srom_1(25842) <= 407130;
srom_1(25843) <= 249161;
srom_1(25844) <= 129361;
srom_1(25845) <= 48292;
srom_1(25846) <= 6333;
srom_1(25847) <= 3682;
srom_1(25848) <= 40350;
srom_1(25849) <= 116166;
srom_1(25850) <= 230775;
srom_1(25851) <= 383638;
srom_1(25852) <= 574039;
srom_1(25853) <= 801086;
srom_1(25854) <= 1063713;
srom_1(25855) <= 1360689;
srom_1(25856) <= 1690621;
srom_1(25857) <= 2051963;
srom_1(25858) <= 2443019;
srom_1(25859) <= 2861956;
srom_1(25860) <= 3306810;
srom_1(25861) <= 3775493;
srom_1(25862) <= 4265810;
srom_1(25863) <= 4775459;
srom_1(25864) <= 5302052;
srom_1(25865) <= 5843118;
srom_1(25866) <= 6396122;
srom_1(25867) <= 6958468;
srom_1(25868) <= 7527522;
srom_1(25869) <= 8100613;
srom_1(25870) <= 8675054;
srom_1(25871) <= 9248153;
srom_1(25872) <= 9817220;
srom_1(25873) <= 10379589;
srom_1(25874) <= 10932621;
srom_1(25875) <= 11473723;
srom_1(25876) <= 12000358;
srom_1(25877) <= 12510056;
srom_1(25878) <= 13000427;
srom_1(25879) <= 13469172;
srom_1(25880) <= 13914093;
srom_1(25881) <= 14333103;
srom_1(25882) <= 14724236;
srom_1(25883) <= 15085660;
srom_1(25884) <= 15415679;
srom_1(25885) <= 15712746;
srom_1(25886) <= 15975467;
srom_1(25887) <= 16202611;
srom_1(25888) <= 16393112;
srom_1(25889) <= 16546078;
srom_1(25890) <= 16660790;
srom_1(25891) <= 16736711;
srom_1(25892) <= 16773485;
srom_1(25893) <= 16770940;
srom_1(25894) <= 16729087;
srom_1(25895) <= 16648122;
srom_1(25896) <= 16528426;
srom_1(25897) <= 16370559;
srom_1(25898) <= 16175262;
srom_1(25899) <= 15943451;
srom_1(25900) <= 15676213;
srom_1(25901) <= 15374800;
srom_1(25902) <= 15040627;
srom_1(25903) <= 14675261;
srom_1(25904) <= 14280414;
srom_1(25905) <= 13857938;
srom_1(25906) <= 13409815;
srom_1(25907) <= 12938145;
srom_1(25908) <= 12445141;
srom_1(25909) <= 11933115;
srom_1(25910) <= 11404467;
srom_1(25911) <= 10861677;
srom_1(25912) <= 10307290;
srom_1(25913) <= 9743905;
srom_1(25914) <= 9174165;
srom_1(25915) <= 8600742;
srom_1(25916) <= 8026323;
srom_1(25917) <= 7453603;
srom_1(25918) <= 6885268;
srom_1(25919) <= 6323983;
srom_1(25920) <= 5772379;
srom_1(25921) <= 5233044;
srom_1(25922) <= 4708506;
srom_1(25923) <= 4201225;
srom_1(25924) <= 3713581;
srom_1(25925) <= 3247859;
srom_1(25926) <= 2806244;
srom_1(25927) <= 2390807;
srom_1(25928) <= 2003495;
srom_1(25929) <= 1646126;
srom_1(25930) <= 1320374;
srom_1(25931) <= 1027767;
srom_1(25932) <= 769678;
srom_1(25933) <= 547317;
srom_1(25934) <= 361726;
srom_1(25935) <= 213777;
srom_1(25936) <= 104161;
srom_1(25937) <= 33395;
srom_1(25938) <= 1808;
srom_1(25939) <= 9551;
srom_1(25940) <= 56585;
srom_1(25941) <= 142692;
srom_1(25942) <= 267466;
srom_1(25943) <= 430323;
srom_1(25944) <= 630499;
srom_1(25945) <= 867056;
srom_1(25946) <= 1138884;
srom_1(25947) <= 1444708;
srom_1(25948) <= 1783094;
srom_1(25949) <= 2152456;
srom_1(25950) <= 2551062;
srom_1(25951) <= 2977042;
srom_1(25952) <= 3428398;
srom_1(25953) <= 3903015;
srom_1(25954) <= 4398666;
srom_1(25955) <= 4913027;
srom_1(25956) <= 5443686;
srom_1(25957) <= 5988156;
srom_1(25958) <= 6543881;
srom_1(25959) <= 7108258;
srom_1(25960) <= 7678638;
srom_1(25961) <= 8252347;
srom_1(25962) <= 8826696;
srom_1(25963) <= 9398990;
srom_1(25964) <= 9966546;
srom_1(25965) <= 10526703;
srom_1(25966) <= 11076833;
srom_1(25967) <= 11614358;
srom_1(25968) <= 12136755;
srom_1(25969) <= 12641577;
srom_1(25970) <= 13126454;
srom_1(25971) <= 13589115;
srom_1(25972) <= 14027388;
srom_1(25973) <= 14439219;
srom_1(25974) <= 14822677;
srom_1(25975) <= 15175963;
srom_1(25976) <= 15497421;
srom_1(25977) <= 15785543;
srom_1(25978) <= 16038979;
srom_1(25979) <= 16256539;
srom_1(25980) <= 16437204;
srom_1(25981) <= 16580126;
srom_1(25982) <= 16684635;
srom_1(25983) <= 16750242;
srom_1(25984) <= 16776637;
srom_1(25985) <= 16763699;
srom_1(25986) <= 16711487;
srom_1(25987) <= 16620246;
srom_1(25988) <= 16490403;
srom_1(25989) <= 16322569;
srom_1(25990) <= 16117530;
srom_1(25991) <= 15876247;
srom_1(25992) <= 15599852;
srom_1(25993) <= 15289641;
srom_1(25994) <= 14947069;
srom_1(25995) <= 14573742;
srom_1(25996) <= 14171411;
srom_1(25997) <= 13741962;
srom_1(25998) <= 13287409;
srom_1(25999) <= 12809884;
srom_1(26000) <= 12311626;
srom_1(26001) <= 11794972;
srom_1(26002) <= 11262345;
srom_1(26003) <= 10716241;
srom_1(26004) <= 10159222;
srom_1(26005) <= 9593900;
srom_1(26006) <= 9022927;
srom_1(26007) <= 8448978;
srom_1(26008) <= 7874747;
srom_1(26009) <= 7302925;
srom_1(26010) <= 6736194;
srom_1(26011) <= 6177212;
srom_1(26012) <= 5628601;
srom_1(26013) <= 5092931;
srom_1(26014) <= 4572716;
srom_1(26015) <= 4070396;
srom_1(26016) <= 3588325;
srom_1(26017) <= 3128764;
srom_1(26018) <= 2693868;
srom_1(26019) <= 2285676;
srom_1(26020) <= 1906104;
srom_1(26021) <= 1556930;
srom_1(26022) <= 1239793;
srom_1(26023) <= 956178;
srom_1(26024) <= 707417;
srom_1(26025) <= 494675;
srom_1(26026) <= 318951;
srom_1(26027) <= 181068;
srom_1(26028) <= 81673;
srom_1(26029) <= 21233;
srom_1(26030) <= 29;
srom_1(26031) <= 18163;
srom_1(26032) <= 75549;
srom_1(26033) <= 171917;
srom_1(26034) <= 306816;
srom_1(26035) <= 479614;
srom_1(26036) <= 689499;
srom_1(26037) <= 935488;
srom_1(26038) <= 1216428;
srom_1(26039) <= 1531000;
srom_1(26040) <= 1877730;
srom_1(26041) <= 2254992;
srom_1(26042) <= 2661016;
srom_1(26043) <= 3093899;
srom_1(26044) <= 3551611;
srom_1(26045) <= 4032005;
srom_1(26046) <= 4532828;
srom_1(26047) <= 5051733;
srom_1(26048) <= 5586285;
srom_1(26049) <= 6133979;
srom_1(26050) <= 6692245;
srom_1(26051) <= 7258466;
srom_1(26052) <= 7829987;
srom_1(26053) <= 8404127;
srom_1(26054) <= 8978194;
srom_1(26055) <= 9549497;
srom_1(26056) <= 10115356;
srom_1(26057) <= 10673117;
srom_1(26058) <= 11220166;
srom_1(26059) <= 11753936;
srom_1(26060) <= 12271926;
srom_1(26061) <= 12771705;
srom_1(26062) <= 13250930;
srom_1(26063) <= 13707354;
srom_1(26064) <= 14138837;
srom_1(26065) <= 14543355;
srom_1(26066) <= 14919011;
srom_1(26067) <= 15264043;
srom_1(26068) <= 15576835;
srom_1(26069) <= 15855919;
srom_1(26070) <= 16099985;
srom_1(26071) <= 16307891;
srom_1(26072) <= 16478660;
srom_1(26073) <= 16611492;
srom_1(26074) <= 16705764;
srom_1(26075) <= 16761034;
srom_1(26076) <= 16777043;
srom_1(26077) <= 16753716;
srom_1(26078) <= 16691162;
srom_1(26079) <= 16589674;
srom_1(26080) <= 16449729;
srom_1(26081) <= 16271982;
srom_1(26082) <= 16057267;
srom_1(26083) <= 15806592;
srom_1(26084) <= 15521131;
srom_1(26085) <= 15202223;
srom_1(26086) <= 14851364;
srom_1(26087) <= 14470198;
srom_1(26088) <= 14060514;
srom_1(26089) <= 13624233;
srom_1(26090) <= 13163400;
srom_1(26091) <= 12680176;
srom_1(26092) <= 12176827;
srom_1(26093) <= 11655714;
srom_1(26094) <= 11119281;
srom_1(26095) <= 10570043;
srom_1(26096) <= 10010575;
srom_1(26097) <= 9443501;
srom_1(26098) <= 8871480;
srom_1(26099) <= 8297195;
srom_1(26100) <= 7723339;
srom_1(26101) <= 7152602;
srom_1(26102) <= 6587662;
srom_1(26103) <= 6031166;
srom_1(26104) <= 5485726;
srom_1(26105) <= 4953898;
srom_1(26106) <= 4438176;
srom_1(26107) <= 3940980;
srom_1(26108) <= 3464640;
srom_1(26109) <= 3011390;
srom_1(26110) <= 2583356;
srom_1(26111) <= 2182544;
srom_1(26112) <= 1810835;
srom_1(26113) <= 1469972;
srom_1(26114) <= 1161552;
srom_1(26115) <= 887022;
srom_1(26116) <= 647670;
srom_1(26117) <= 444618;
srom_1(26118) <= 278818;
srom_1(26119) <= 151047;
srom_1(26120) <= 61905;
srom_1(26121) <= 11810;
srom_1(26122) <= 997;
srom_1(26123) <= 29516;
srom_1(26124) <= 97234;
srom_1(26125) <= 203832;
srom_1(26126) <= 348812;
srom_1(26127) <= 531494;
srom_1(26128) <= 751020;
srom_1(26129) <= 1006361;
srom_1(26130) <= 1296320;
srom_1(26131) <= 1619538;
srom_1(26132) <= 1974497;
srom_1(26133) <= 2359535;
srom_1(26134) <= 2772845;
srom_1(26135) <= 3212490;
srom_1(26136) <= 3676407;
srom_1(26137) <= 4162421;
srom_1(26138) <= 4668253;
srom_1(26139) <= 5191531;
srom_1(26140) <= 5729802;
srom_1(26141) <= 6280540;
srom_1(26142) <= 6841164;
srom_1(26143) <= 7409045;
srom_1(26144) <= 7981518;
srom_1(26145) <= 8555901;
srom_1(26146) <= 9129500;
srom_1(26147) <= 9699624;
srom_1(26148) <= 10263600;
srom_1(26149) <= 10818784;
srom_1(26150) <= 11362571;
srom_1(26151) <= 11892413;
srom_1(26152) <= 12405825;
srom_1(26153) <= 12900398;
srom_1(26154) <= 13373814;
srom_1(26155) <= 13823852;
srom_1(26156) <= 14248403;
srom_1(26157) <= 14645475;
srom_1(26158) <= 15013207;
srom_1(26159) <= 15349873;
srom_1(26160) <= 15653896;
srom_1(26161) <= 15923849;
srom_1(26162) <= 16158467;
srom_1(26163) <= 16356650;
srom_1(26164) <= 16517467;
srom_1(26165) <= 16640166;
srom_1(26166) <= 16724170;
srom_1(26167) <= 16769086;
srom_1(26168) <= 16774703;
srom_1(26169) <= 16740994;
srom_1(26170) <= 16668119;
srom_1(26171) <= 16556417;
srom_1(26172) <= 16406415;
srom_1(26173) <= 16218814;
srom_1(26174) <= 15994494;
srom_1(26175) <= 15734508;
srom_1(26176) <= 15440074;
srom_1(26177) <= 15112574;
srom_1(26178) <= 14753542;
srom_1(26179) <= 14364664;
srom_1(26180) <= 13947761;
srom_1(26181) <= 13504790;
srom_1(26182) <= 13037827;
srom_1(26183) <= 12549062;
srom_1(26184) <= 12040788;
srom_1(26185) <= 11515387;
srom_1(26186) <= 10975324;
srom_1(26187) <= 10423130;
srom_1(26188) <= 9861396;
srom_1(26189) <= 9292756;
srom_1(26190) <= 8719876;
srom_1(26191) <= 8145442;
srom_1(26192) <= 7572149;
srom_1(26193) <= 7002684;
srom_1(26194) <= 6439718;
srom_1(26195) <= 5885892;
srom_1(26196) <= 5343801;
srom_1(26197) <= 4815989;
srom_1(26198) <= 4304929;
srom_1(26199) <= 3813020;
srom_1(26200) <= 3342567;
srom_1(26201) <= 2895777;
srom_1(26202) <= 2474744;
srom_1(26203) <= 2081444;
srom_1(26204) <= 1717720;
srom_1(26205) <= 1385278;
srom_1(26206) <= 1085677;
srom_1(26207) <= 820322;
srom_1(26208) <= 590458;
srom_1(26209) <= 397161;
srom_1(26210) <= 241339;
srom_1(26211) <= 123723;
srom_1(26212) <= 44863;
srom_1(26213) <= 5130;
srom_1(26214) <= 4710;
srom_1(26215) <= 43605;
srom_1(26216) <= 121633;
srom_1(26217) <= 238427;
srom_1(26218) <= 393441;
srom_1(26219) <= 585946;
srom_1(26220) <= 815041;
srom_1(26221) <= 1079651;
srom_1(26222) <= 1378535;
srom_1(26223) <= 1710291;
srom_1(26224) <= 2073365;
srom_1(26225) <= 2466053;
srom_1(26226) <= 2886513;
srom_1(26227) <= 3332775;
srom_1(26228) <= 3802746;
srom_1(26229) <= 4294221;
srom_1(26230) <= 4804896;
srom_1(26231) <= 5332377;
srom_1(26232) <= 5874189;
srom_1(26233) <= 6427792;
srom_1(26234) <= 6990590;
srom_1(26235) <= 7559944;
srom_1(26236) <= 8133183;
srom_1(26237) <= 8707621;
srom_1(26238) <= 9280562;
srom_1(26239) <= 9849321;
srom_1(26240) <= 10411230;
srom_1(26241) <= 10963654;
srom_1(26242) <= 11504003;
srom_1(26243) <= 12029743;
srom_1(26244) <= 12538408;
srom_1(26245) <= 13027614;
srom_1(26246) <= 13495065;
srom_1(26247) <= 13938571;
srom_1(26248) <= 14356051;
srom_1(26249) <= 14745547;
srom_1(26250) <= 15105234;
srom_1(26251) <= 15433424;
srom_1(26252) <= 15728578;
srom_1(26253) <= 15989313;
srom_1(26254) <= 16214405;
srom_1(26255) <= 16402800;
srom_1(26256) <= 16553613;
srom_1(26257) <= 16666138;
srom_1(26258) <= 16739847;
srom_1(26259) <= 16774394;
srom_1(26260) <= 16769616;
srom_1(26261) <= 16725538;
srom_1(26262) <= 16642365;
srom_1(26263) <= 16520487;
srom_1(26264) <= 16360476;
srom_1(26265) <= 16163082;
srom_1(26266) <= 15929231;
srom_1(26267) <= 15660019;
srom_1(26268) <= 15356709;
srom_1(26269) <= 15020723;
srom_1(26270) <= 14653637;
srom_1(26271) <= 14257172;
srom_1(26272) <= 13833188;
srom_1(26273) <= 13383672;
srom_1(26274) <= 12910732;
srom_1(26275) <= 12416587;
srom_1(26276) <= 11903553;
srom_1(26277) <= 11374036;
srom_1(26278) <= 10830519;
srom_1(26279) <= 10275552;
srom_1(26280) <= 9711736;
srom_1(26281) <= 9141715;
srom_1(26282) <= 8568163;
srom_1(26283) <= 7993768;
srom_1(26284) <= 7421226;
srom_1(26285) <= 6853219;
srom_1(26286) <= 6292413;
srom_1(26287) <= 5741436;
srom_1(26288) <= 5202873;
srom_1(26289) <= 4679249;
srom_1(26290) <= 4173020;
srom_1(26291) <= 3686558;
srom_1(26292) <= 3222146;
srom_1(26293) <= 2781962;
srom_1(26294) <= 2368069;
srom_1(26295) <= 1982408;
srom_1(26296) <= 1626789;
srom_1(26297) <= 1302877;
srom_1(26298) <= 1012193;
srom_1(26299) <= 756100;
srom_1(26300) <= 535798;
srom_1(26301) <= 352321;
srom_1(26302) <= 206528;
srom_1(26303) <= 99104;
srom_1(26304) <= 30553;
srom_1(26305) <= 1195;
srom_1(26306) <= 11169;
srom_1(26307) <= 60427;
srom_1(26308) <= 148739;
srom_1(26309) <= 275691;
srom_1(26310) <= 440687;
srom_1(26311) <= 642953;
srom_1(26312) <= 881541;
srom_1(26313) <= 1155333;
srom_1(26314) <= 1463044;
srom_1(26315) <= 1803231;
srom_1(26316) <= 2174300;
srom_1(26317) <= 2574509;
srom_1(26318) <= 3001983;
srom_1(26319) <= 3454716;
srom_1(26320) <= 3930586;
srom_1(26321) <= 4427361;
srom_1(26322) <= 4942712;
srom_1(26323) <= 5474222;
srom_1(26324) <= 6019399;
srom_1(26325) <= 6575685;
srom_1(26326) <= 7140473;
srom_1(26327) <= 7711114;
srom_1(26328) <= 8284932;
srom_1(26329) <= 8859236;
srom_1(26330) <= 9431333;
srom_1(26331) <= 9998540;
srom_1(26332) <= 10558198;
srom_1(26333) <= 11107682;
srom_1(26334) <= 11644415;
srom_1(26335) <= 12165881;
srom_1(26336) <= 12669633;
srom_1(26337) <= 13153311;
srom_1(26338) <= 13614645;
srom_1(26339) <= 14051472;
srom_1(26340) <= 14461745;
srom_1(26341) <= 14843538;
srom_1(26342) <= 15195062;
srom_1(26343) <= 15514668;
srom_1(26344) <= 15800857;
srom_1(26345) <= 16052288;
srom_1(26346) <= 16267782;
srom_1(26347) <= 16446327;
srom_1(26348) <= 16587086;
srom_1(26349) <= 16689401;
srom_1(26350) <= 16752790;
srom_1(26351) <= 16776956;
srom_1(26352) <= 16761787;
srom_1(26353) <= 16707352;
srom_1(26354) <= 16613909;
srom_1(26355) <= 16481894;
srom_1(26356) <= 16311927;
srom_1(26357) <= 16104805;
srom_1(26358) <= 15861498;
srom_1(26359) <= 15583149;
srom_1(26360) <= 15271062;
srom_1(26361) <= 14926701;
srom_1(26362) <= 14551681;
srom_1(26363) <= 14147760;
srom_1(26364) <= 13716832;
srom_1(26365) <= 13260918;
srom_1(26366) <= 12782157;
srom_1(26367) <= 12282792;
srom_1(26368) <= 11765167;
srom_1(26369) <= 11231707;
srom_1(26370) <= 10684915;
srom_1(26371) <= 10127355;
srom_1(26372) <= 9561642;
srom_1(26373) <= 8990427;
srom_1(26374) <= 8416391;
srom_1(26375) <= 7842224;
srom_1(26376) <= 7270620;
srom_1(26377) <= 6704258;
srom_1(26378) <= 6145794;
srom_1(26379) <= 5597848;
srom_1(26380) <= 5062989;
srom_1(26381) <= 4543724;
srom_1(26382) <= 4042490;
srom_1(26383) <= 3561636;
srom_1(26384) <= 3103417;
srom_1(26385) <= 2669983;
srom_1(26386) <= 2263365;
srom_1(26387) <= 1885470;
srom_1(26388) <= 1538071;
srom_1(26389) <= 1222796;
srom_1(26390) <= 941125;
srom_1(26391) <= 694377;
srom_1(26392) <= 483710;
srom_1(26393) <= 310111;
srom_1(26394) <= 174396;
srom_1(26395) <= 77200;
srom_1(26396) <= 18979;
srom_1(26397) <= 6;
srom_1(26398) <= 20370;
srom_1(26399) <= 79975;
srom_1(26400) <= 178543;
srom_1(26401) <= 315610;
srom_1(26402) <= 490534;
srom_1(26403) <= 702496;
srom_1(26404) <= 950500;
srom_1(26405) <= 1233383;
srom_1(26406) <= 1549821;
srom_1(26407) <= 1898327;
srom_1(26408) <= 2277269;
srom_1(26409) <= 2684869;
srom_1(26410) <= 3119215;
srom_1(26411) <= 3578272;
srom_1(26412) <= 4059886;
srom_1(26413) <= 4561799;
srom_1(26414) <= 5081657;
srom_1(26415) <= 5617022;
srom_1(26416) <= 6165385;
srom_1(26417) <= 6724172;
srom_1(26418) <= 7290765;
srom_1(26419) <= 7862506;
srom_1(26420) <= 8436714;
srom_1(26421) <= 9010697;
srom_1(26422) <= 9581762;
srom_1(26423) <= 10147233;
srom_1(26424) <= 10704456;
srom_1(26425) <= 11250820;
srom_1(26426) <= 11783761;
srom_1(26427) <= 12300782;
srom_1(26428) <= 12799457;
srom_1(26429) <= 13277448;
srom_1(26430) <= 13732514;
srom_1(26431) <= 14162520;
srom_1(26432) <= 14565450;
srom_1(26433) <= 14939416;
srom_1(26434) <= 15282662;
srom_1(26435) <= 15593579;
srom_1(26436) <= 15870710;
srom_1(26437) <= 16112755;
srom_1(26438) <= 16318578;
srom_1(26439) <= 16487215;
srom_1(26440) <= 16617875;
srom_1(26441) <= 16709945;
srom_1(26442) <= 16762994;
srom_1(26443) <= 16776772;
srom_1(26444) <= 16751215;
srom_1(26445) <= 16686443;
srom_1(26446) <= 16582760;
srom_1(26447) <= 16440651;
srom_1(26448) <= 16260784;
srom_1(26449) <= 16044001;
srom_1(26450) <= 15791320;
srom_1(26451) <= 15503924;
srom_1(26452) <= 15183163;
srom_1(26453) <= 14830539;
srom_1(26454) <= 14447707;
srom_1(26455) <= 14036462;
srom_1(26456) <= 13598732;
srom_1(26457) <= 13136570;
srom_1(26458) <= 12652143;
srom_1(26459) <= 12147723;
srom_1(26460) <= 11625675;
srom_1(26461) <= 11088448;
srom_1(26462) <= 10538560;
srom_1(26463) <= 9978590;
srom_1(26464) <= 9411164;
srom_1(26465) <= 8838943;
srom_1(26466) <= 8264610;
srom_1(26467) <= 7690859;
srom_1(26468) <= 7120379;
srom_1(26469) <= 6555847;
srom_1(26470) <= 5999910;
srom_1(26471) <= 5455173;
srom_1(26472) <= 4924193;
srom_1(26473) <= 4409458;
srom_1(26474) <= 3913383;
srom_1(26475) <= 3438294;
srom_1(26476) <= 2986418;
srom_1(26477) <= 2559876;
srom_1(26478) <= 2160666;
srom_1(26479) <= 1790661;
srom_1(26480) <= 1451596;
srom_1(26481) <= 1145061;
srom_1(26482) <= 872494;
srom_1(26483) <= 635172;
srom_1(26484) <= 434209;
srom_1(26485) <= 270547;
srom_1(26486) <= 144953;
srom_1(26487) <= 58016;
srom_1(26488) <= 10145;
srom_1(26489) <= 1563;
srom_1(26490) <= 32310;
srom_1(26491) <= 102243;
srom_1(26492) <= 211034;
srom_1(26493) <= 358172;
srom_1(26494) <= 542968;
srom_1(26495) <= 764555;
srom_1(26496) <= 1021893;
srom_1(26497) <= 1313777;
srom_1(26498) <= 1638836;
srom_1(26499) <= 1995548;
srom_1(26500) <= 2382239;
srom_1(26501) <= 2797096;
srom_1(26502) <= 3238173;
srom_1(26503) <= 3703403;
srom_1(26504) <= 4190603;
srom_1(26505) <= 4697489;
srom_1(26506) <= 5221684;
srom_1(26507) <= 5760729;
srom_1(26508) <= 6312098;
srom_1(26509) <= 6873204;
srom_1(26510) <= 7441417;
srom_1(26511) <= 8014071;
srom_1(26512) <= 8588481;
srom_1(26513) <= 9161954;
srom_1(26514) <= 9731801;
srom_1(26515) <= 10295349;
srom_1(26516) <= 10849956;
srom_1(26517) <= 11393020;
srom_1(26518) <= 11921996;
srom_1(26519) <= 12434402;
srom_1(26520) <= 12927837;
srom_1(26521) <= 13399985;
srom_1(26522) <= 13848633;
srom_1(26523) <= 14271677;
srom_1(26524) <= 14667134;
srom_1(26525) <= 15033148;
srom_1(26526) <= 15368004;
srom_1(26527) <= 15670131;
srom_1(26528) <= 15938113;
srom_1(26529) <= 16170692;
srom_1(26530) <= 16366778;
srom_1(26531) <= 16525452;
srom_1(26532) <= 16645970;
srom_1(26533) <= 16727766;
srom_1(26534) <= 16770457;
srom_1(26535) <= 16773842;
srom_1(26536) <= 16737906;
srom_1(26537) <= 16662818;
srom_1(26538) <= 16548928;
srom_1(26539) <= 16396772;
srom_1(26540) <= 16207064;
srom_1(26541) <= 15980691;
srom_1(26542) <= 15718717;
srom_1(26543) <= 15422370;
srom_1(26544) <= 15093038;
srom_1(26545) <= 14732268;
srom_1(26546) <= 14341749;
srom_1(26547) <= 13923315;
srom_1(26548) <= 13478926;
srom_1(26549) <= 13010667;
srom_1(26550) <= 12520733;
srom_1(26551) <= 12011423;
srom_1(26552) <= 11485124;
srom_1(26553) <= 10944304;
srom_1(26554) <= 10391500;
srom_1(26555) <= 9829304;
srom_1(26556) <= 9260351;
srom_1(26557) <= 8687311;
srom_1(26558) <= 8112870;
srom_1(26559) <= 7539722;
srom_1(26560) <= 6970554;
srom_1(26561) <= 6408037;
srom_1(26562) <= 5854807;
srom_1(26563) <= 5313459;
srom_1(26564) <= 4786531;
srom_1(26565) <= 4276495;
srom_1(26566) <= 3785741;
srom_1(26567) <= 3316573;
srom_1(26568) <= 2871188;
srom_1(26569) <= 2451677;
srom_1(26570) <= 2060006;
srom_1(26571) <= 1698012;
srom_1(26572) <= 1367393;
srom_1(26573) <= 1069698;
srom_1(26574) <= 806324;
srom_1(26575) <= 578506;
srom_1(26576) <= 387313;
srom_1(26577) <= 233640;
srom_1(26578) <= 118209;
srom_1(26579) <= 41560;
srom_1(26580) <= 4054;
srom_1(26581) <= 5866;
srom_1(26582) <= 46987;
srom_1(26583) <= 127225;
srom_1(26584) <= 246203;
srom_1(26585) <= 403364;
srom_1(26586) <= 597970;
srom_1(26587) <= 829110;
srom_1(26588) <= 1095698;
srom_1(26589) <= 1396486;
srom_1(26590) <= 1730062;
srom_1(26591) <= 2094862;
srom_1(26592) <= 2489176;
srom_1(26593) <= 2911154;
srom_1(26594) <= 3358817;
srom_1(26595) <= 3830068;
srom_1(26596) <= 4322694;
srom_1(26597) <= 4834387;
srom_1(26598) <= 5362748;
srom_1(26599) <= 5905297;
srom_1(26600) <= 6459492;
srom_1(26601) <= 7022732;
srom_1(26602) <= 7592378;
srom_1(26603) <= 8165758;
srom_1(26604) <= 8740183;
srom_1(26605) <= 9312959;
srom_1(26606) <= 9881400;
srom_1(26607) <= 10442841;
srom_1(26608) <= 10994649;
srom_1(26609) <= 11534237;
srom_1(26610) <= 12059073;
srom_1(26611) <= 12566698;
srom_1(26612) <= 13054730;
srom_1(26613) <= 13520881;
srom_1(26614) <= 13962965;
srom_1(26615) <= 14378909;
srom_1(26616) <= 14766762;
srom_1(26617) <= 15124706;
srom_1(26618) <= 15451062;
srom_1(26619) <= 15744300;
srom_1(26620) <= 16003044;
srom_1(26621) <= 16226082;
srom_1(26622) <= 16412367;
srom_1(26623) <= 16561026;
srom_1(26624) <= 16671361;
srom_1(26625) <= 16742856;
srom_1(26626) <= 16775175;
srom_1(26627) <= 16768167;
srom_1(26628) <= 16721864;
srom_1(26629) <= 16636483;
srom_1(26630) <= 16512425;
srom_1(26631) <= 16350272;
srom_1(26632) <= 16150784;
srom_1(26633) <= 15914896;
srom_1(26634) <= 15643715;
srom_1(26635) <= 15338512;
srom_1(26636) <= 15000719;
srom_1(26637) <= 14631919;
srom_1(26638) <= 14233843;
srom_1(26639) <= 13808356;
srom_1(26640) <= 13357454;
srom_1(26641) <= 12883251;
srom_1(26642) <= 12387971;
srom_1(26643) <= 11873937;
srom_1(26644) <= 11343559;
srom_1(26645) <= 10799324;
srom_1(26646) <= 10243785;
srom_1(26647) <= 9679546;
srom_1(26648) <= 9109253;
srom_1(26649) <= 8535581;
srom_1(26650) <= 7961220;
srom_1(26651) <= 7388863;
srom_1(26652) <= 6821194;
srom_1(26653) <= 6260875;
srom_1(26654) <= 5710534;
srom_1(26655) <= 5172751;
srom_1(26656) <= 4650049;
srom_1(26657) <= 4144877;
srom_1(26658) <= 3659607;
srom_1(26659) <= 3196512;
srom_1(26660) <= 2757764;
srom_1(26661) <= 2345422;
srom_1(26662) <= 1961418;
srom_1(26663) <= 1607554;
srom_1(26664) <= 1285488;
srom_1(26665) <= 996731;
srom_1(26666) <= 742637;
srom_1(26667) <= 524398;
srom_1(26668) <= 343036;
srom_1(26669) <= 199403;
srom_1(26670) <= 94172;
srom_1(26671) <= 27837;
srom_1(26672) <= 708;
srom_1(26673) <= 12913;
srom_1(26674) <= 64394;
srom_1(26675) <= 154911;
srom_1(26676) <= 284038;
srom_1(26677) <= 451170;
srom_1(26678) <= 655523;
srom_1(26679) <= 896140;
srom_1(26680) <= 1171891;
srom_1(26681) <= 1481484;
srom_1(26682) <= 1823467;
srom_1(26683) <= 2196236;
srom_1(26684) <= 2598044;
srom_1(26685) <= 3027005;
srom_1(26686) <= 3481108;
srom_1(26687) <= 3958225;
srom_1(26688) <= 4456117;
srom_1(26689) <= 4972450;
srom_1(26690) <= 5504802;
srom_1(26691) <= 6050678;
srom_1(26692) <= 6607517;
srom_1(26693) <= 7172708;
srom_1(26694) <= 7743600;
srom_1(26695) <= 8317518;
srom_1(26696) <= 8891769;
srom_1(26697) <= 9463660;
srom_1(26698) <= 10030510;
srom_1(26699) <= 10589661;
srom_1(26700) <= 11138490;
srom_1(26701) <= 11674424;
srom_1(26702) <= 12194949;
srom_1(26703) <= 12697626;
srom_1(26704) <= 13180096;
srom_1(26705) <= 13640097;
srom_1(26706) <= 14075472;
srom_1(26707) <= 14484179;
srom_1(26708) <= 14864302;
srom_1(26709) <= 15214058;
srom_1(26710) <= 15531807;
srom_1(26711) <= 15816060;
srom_1(26712) <= 16065482;
srom_1(26713) <= 16278905;
srom_1(26714) <= 16455328;
srom_1(26715) <= 16593923;
srom_1(26716) <= 16694041;
srom_1(26717) <= 16755211;
srom_1(26718) <= 16777148;
srom_1(26719) <= 16759748;
srom_1(26720) <= 16703093;
srom_1(26721) <= 16607448;
srom_1(26722) <= 16473262;
srom_1(26723) <= 16301165;
srom_1(26724) <= 16091963;
srom_1(26725) <= 15846637;
srom_1(26726) <= 15566338;
srom_1(26727) <= 15252380;
srom_1(26728) <= 14906235;
srom_1(26729) <= 14529527;
srom_1(26730) <= 14124022;
srom_1(26731) <= 13691622;
srom_1(26732) <= 13234354;
srom_1(26733) <= 12754363;
srom_1(26734) <= 12253899;
srom_1(26735) <= 11735310;
srom_1(26736) <= 11201027;
srom_1(26737) <= 10653555;
srom_1(26738) <= 10095462;
srom_1(26739) <= 9529365;
srom_1(26740) <= 8957919;
srom_1(26741) <= 8383803;
srom_1(26742) <= 7809710;
srom_1(26743) <= 7238331;
srom_1(26744) <= 6672346;
srom_1(26745) <= 6114410;
srom_1(26746) <= 5567138;
srom_1(26747) <= 5033096;
srom_1(26748) <= 4514790;
srom_1(26749) <= 4014650;
srom_1(26750) <= 3535020;
srom_1(26751) <= 3078151;
srom_1(26752) <= 2646184;
srom_1(26753) <= 2241145;
srom_1(26754) <= 1864934;
srom_1(26755) <= 1519315;
srom_1(26756) <= 1205908;
srom_1(26757) <= 926184;
srom_1(26758) <= 681453;
srom_1(26759) <= 472863;
srom_1(26760) <= 301394;
srom_1(26761) <= 167848;
srom_1(26762) <= 72852;
srom_1(26763) <= 16851;
srom_1(26764) <= 108;
srom_1(26765) <= 22702;
srom_1(26766) <= 84527;
srom_1(26767) <= 185292;
srom_1(26768) <= 324526;
srom_1(26769) <= 501574;
srom_1(26770) <= 715608;
srom_1(26771) <= 965623;
srom_1(26772) <= 1250447;
srom_1(26773) <= 1568744;
srom_1(26774) <= 1919022;
srom_1(26775) <= 2299638;
srom_1(26776) <= 2708807;
srom_1(26777) <= 3144611;
srom_1(26778) <= 3605006;
srom_1(26779) <= 4087832;
srom_1(26780) <= 4590827;
srom_1(26781) <= 5111630;
srom_1(26782) <= 5647801;
srom_1(26783) <= 6196824;
srom_1(26784) <= 6756125;
srom_1(26785) <= 7323081;
srom_1(26786) <= 7895034;
srom_1(26787) <= 8469301;
srom_1(26788) <= 9043190;
srom_1(26789) <= 9614010;
srom_1(26790) <= 10179083;
srom_1(26791) <= 10735760;
srom_1(26792) <= 11281430;
srom_1(26793) <= 11813535;
srom_1(26794) <= 12329579;
srom_1(26795) <= 12827143;
srom_1(26796) <= 13303893;
srom_1(26797) <= 13757593;
srom_1(26798) <= 14186116;
srom_1(26799) <= 14587453;
srom_1(26800) <= 14959722;
srom_1(26801) <= 15301176;
srom_1(26802) <= 15610214;
srom_1(26803) <= 15885388;
srom_1(26804) <= 16125407;
srom_1(26805) <= 16329146;
srom_1(26806) <= 16495649;
srom_1(26807) <= 16624135;
srom_1(26808) <= 16714001;
srom_1(26809) <= 16764827;
srom_1(26810) <= 16776375;
srom_1(26811) <= 16748589;
srom_1(26812) <= 16681600;
srom_1(26813) <= 16575722;
srom_1(26814) <= 16431452;
srom_1(26815) <= 16249467;
srom_1(26816) <= 16030619;
srom_1(26817) <= 15775936;
srom_1(26818) <= 15486610;
srom_1(26819) <= 15164000;
srom_1(26820) <= 14809617;
srom_1(26821) <= 14425124;
srom_1(26822) <= 14012324;
srom_1(26823) <= 13573152;
srom_1(26824) <= 13109669;
srom_1(26825) <= 12624046;
srom_1(26826) <= 12118562;
srom_1(26827) <= 11595587;
srom_1(26828) <= 11057573;
srom_1(26829) <= 10507044;
srom_1(26830) <= 9946581;
srom_1(26831) <= 9378811;
srom_1(26832) <= 8806399;
srom_1(26833) <= 8232027;
srom_1(26834) <= 7658389;
srom_1(26835) <= 7088176;
srom_1(26836) <= 6524061;
srom_1(26837) <= 5968689;
srom_1(26838) <= 5424665;
srom_1(26839) <= 4894540;
srom_1(26840) <= 4380800;
srom_1(26841) <= 3885854;
srom_1(26842) <= 3412023;
srom_1(26843) <= 2961529;
srom_1(26844) <= 2536484;
srom_1(26845) <= 2138882;
srom_1(26846) <= 1770586;
srom_1(26847) <= 1433326;
srom_1(26848) <= 1128680;
srom_1(26849) <= 858079;
srom_1(26850) <= 622792;
srom_1(26851) <= 423921;
srom_1(26852) <= 262399;
srom_1(26853) <= 138983;
srom_1(26854) <= 54253;
srom_1(26855) <= 8606;
srom_1(26856) <= 2255;
srom_1(26857) <= 35231;
srom_1(26858) <= 107378;
srom_1(26859) <= 218360;
srom_1(26860) <= 367654;
srom_1(26861) <= 554561;
srom_1(26862) <= 778205;
srom_1(26863) <= 1037536;
srom_1(26864) <= 1331340;
srom_1(26865) <= 1658237;
srom_1(26866) <= 2016695;
srom_1(26867) <= 2405033;
srom_1(26868) <= 2821431;
srom_1(26869) <= 3263934;
srom_1(26870) <= 3730469;
srom_1(26871) <= 4218848;
srom_1(26872) <= 4726780;
srom_1(26873) <= 5251884;
srom_1(26874) <= 5791697;
srom_1(26875) <= 6343687;
srom_1(26876) <= 6905267;
srom_1(26877) <= 7473803;
srom_1(26878) <= 8046629;
srom_1(26879) <= 8621058;
srom_1(26880) <= 9194397;
srom_1(26881) <= 9763958;
srom_1(26882) <= 10327069;
srom_1(26883) <= 10881090;
srom_1(26884) <= 11423423;
srom_1(26885) <= 11951525;
srom_1(26886) <= 12462919;
srom_1(26887) <= 12955207;
srom_1(26888) <= 13426081;
srom_1(26889) <= 13873332;
srom_1(26890) <= 14294863;
srom_1(26891) <= 14688698;
srom_1(26892) <= 15052990;
srom_1(26893) <= 15386030;
srom_1(26894) <= 15686257;
srom_1(26895) <= 15952262;
srom_1(26896) <= 16182799;
srom_1(26897) <= 16376787;
srom_1(26898) <= 16533315;
srom_1(26899) <= 16651650;
srom_1(26900) <= 16731236;
srom_1(26901) <= 16771701;
srom_1(26902) <= 16772855;
srom_1(26903) <= 16734692;
srom_1(26904) <= 16657392;
srom_1(26905) <= 16541316;
srom_1(26906) <= 16387009;
srom_1(26907) <= 16195196;
srom_1(26908) <= 15966774;
srom_1(26909) <= 15702816;
srom_1(26910) <= 15404559;
srom_1(26911) <= 15073402;
srom_1(26912) <= 14710897;
srom_1(26913) <= 14318745;
srom_1(26914) <= 13898785;
srom_1(26915) <= 13452985;
srom_1(26916) <= 12983437;
srom_1(26917) <= 12492342;
srom_1(26918) <= 11982004;
srom_1(26919) <= 11454814;
srom_1(26920) <= 10913247;
srom_1(26921) <= 10359840;
srom_1(26922) <= 9797189;
srom_1(26923) <= 9227933;
srom_1(26924) <= 8654742;
srom_1(26925) <= 8080302;
srom_1(26926) <= 7507308;
srom_1(26927) <= 6938446;
srom_1(26928) <= 6376385;
srom_1(26929) <= 5823760;
srom_1(26930) <= 5283163;
srom_1(26931) <= 4757128;
srom_1(26932) <= 4248122;
srom_1(26933) <= 3758532;
srom_1(26934) <= 3290655;
srom_1(26935) <= 2846683;
srom_1(26936) <= 2428699;
srom_1(26937) <= 2038664;
srom_1(26938) <= 1678405;
srom_1(26939) <= 1349613;
srom_1(26940) <= 1053829;
srom_1(26941) <= 792441;
srom_1(26942) <= 566673;
srom_1(26943) <= 377586;
srom_1(26944) <= 226064;
srom_1(26945) <= 112820;
srom_1(26946) <= 38383;
srom_1(26947) <= 3104;
srom_1(26948) <= 7147;
srom_1(26949) <= 50494;
srom_1(26950) <= 132941;
srom_1(26951) <= 254102;
srom_1(26952) <= 413408;
srom_1(26953) <= 610113;
srom_1(26954) <= 843293;
srom_1(26955) <= 1111856;
srom_1(26956) <= 1414543;
srom_1(26957) <= 1749933;
srom_1(26958) <= 2116454;
srom_1(26959) <= 2512388;
srom_1(26960) <= 2935877;
srom_1(26961) <= 3384935;
srom_1(26962) <= 3857458;
srom_1(26963) <= 4351229;
srom_1(26964) <= 4863932;
srom_1(26965) <= 5393164;
srom_1(26966) <= 5936443;
srom_1(26967) <= 6491220;
srom_1(26968) <= 7054896;
srom_1(26969) <= 7624825;
srom_1(26970) <= 8198336;
srom_1(26971) <= 8772739;
srom_1(26972) <= 9345341;
srom_1(26973) <= 9913456;
srom_1(26974) <= 10474421;
srom_1(26975) <= 11025605;
srom_1(26976) <= 11564423;
srom_1(26977) <= 12088348;
srom_1(26978) <= 12594924;
srom_1(26979) <= 13081776;
srom_1(26980) <= 13546619;
srom_1(26981) <= 13987275;
srom_1(26982) <= 14401676;
srom_1(26983) <= 14787881;
srom_1(26984) <= 15144076;
srom_1(26985) <= 15468594;
srom_1(26986) <= 15759910;
srom_1(26987) <= 16016660;
srom_1(26988) <= 16237640;
srom_1(26989) <= 16421812;
srom_1(26990) <= 16568315;
srom_1(26991) <= 16676459;
srom_1(26992) <= 16745740;
srom_1(26993) <= 16775830;
srom_1(26994) <= 16766590;
srom_1(26995) <= 16718063;
srom_1(26996) <= 16630476;
srom_1(26997) <= 16504241;
srom_1(26998) <= 16339948;
srom_1(26999) <= 16138369;
srom_1(27000) <= 15900448;
srom_1(27001) <= 15627302;
srom_1(27002) <= 15320211;
srom_1(27003) <= 14980615;
srom_1(27004) <= 14610107;
srom_1(27005) <= 14210425;
srom_1(27006) <= 13783442;
srom_1(27007) <= 13331160;
srom_1(27008) <= 12855702;
srom_1(27009) <= 12359295;
srom_1(27010) <= 11844269;
srom_1(27011) <= 11313038;
srom_1(27012) <= 10768093;
srom_1(27013) <= 10211990;
srom_1(27014) <= 9647337;
srom_1(27015) <= 9076780;
srom_1(27016) <= 8502997;
srom_1(27017) <= 7928678;
srom_1(27018) <= 7356515;
srom_1(27019) <= 6789192;
srom_1(27020) <= 6229369;
srom_1(27021) <= 5679672;
srom_1(27022) <= 5142677;
srom_1(27023) <= 4620904;
srom_1(27024) <= 4116799;
srom_1(27025) <= 3632726;
srom_1(27026) <= 3170955;
srom_1(27027) <= 2733652;
srom_1(27028) <= 2322866;
srom_1(27029) <= 1940525;
srom_1(27030) <= 1588421;
srom_1(27031) <= 1268205;
srom_1(27032) <= 981380;
srom_1(27033) <= 729289;
srom_1(27034) <= 513116;
srom_1(27035) <= 333873;
srom_1(27036) <= 192402;
srom_1(27037) <= 89366;
srom_1(27038) <= 25247;
srom_1(27039) <= 348;
srom_1(27040) <= 14784;
srom_1(27041) <= 68487;
srom_1(27042) <= 161207;
srom_1(27043) <= 292507;
srom_1(27044) <= 461773;
srom_1(27045) <= 668211;
srom_1(27046) <= 910852;
srom_1(27047) <= 1188559;
srom_1(27048) <= 1500029;
srom_1(27049) <= 1843802;
srom_1(27050) <= 2218267;
srom_1(27051) <= 2621666;
srom_1(27052) <= 3052108;
srom_1(27053) <= 3507575;
srom_1(27054) <= 3985930;
srom_1(27055) <= 4484932;
srom_1(27056) <= 5002239;
srom_1(27057) <= 5535425;
srom_1(27058) <= 6081992;
srom_1(27059) <= 6639375;
srom_1(27060) <= 7204960;
srom_1(27061) <= 7776097;
srom_1(27062) <= 8350105;
srom_1(27063) <= 8924294;
srom_1(27064) <= 9495971;
srom_1(27065) <= 10062455;
srom_1(27066) <= 10621090;
srom_1(27067) <= 11169256;
srom_1(27068) <= 11704383;
srom_1(27069) <= 12223961;
srom_1(27070) <= 12725553;
srom_1(27071) <= 13206808;
srom_1(27072) <= 13665469;
srom_1(27073) <= 14099385;
srom_1(27074) <= 14506521;
srom_1(27075) <= 14884968;
srom_1(27076) <= 15232951;
srom_1(27077) <= 15548839;
srom_1(27078) <= 15831150;
srom_1(27079) <= 16078561;
srom_1(27080) <= 16289910;
srom_1(27081) <= 16464208;
srom_1(27082) <= 16600636;
srom_1(27083) <= 16698556;
srom_1(27084) <= 16757507;
srom_1(27085) <= 16777213;
srom_1(27086) <= 16757583;
srom_1(27087) <= 16698707;
srom_1(27088) <= 16600863;
srom_1(27089) <= 16464508;
srom_1(27090) <= 16290283;
srom_1(27091) <= 16079004;
srom_1(27092) <= 15831662;
srom_1(27093) <= 15549418;
srom_1(27094) <= 15233593;
srom_1(27095) <= 14885670;
srom_1(27096) <= 14507281;
srom_1(27097) <= 14100198;
srom_1(27098) <= 13666332;
srom_1(27099) <= 13207717;
srom_1(27100) <= 12726503;
srom_1(27101) <= 12224948;
srom_1(27102) <= 11705403;
srom_1(27103) <= 11170304;
srom_1(27104) <= 10622160;
srom_1(27105) <= 10063543;
srom_1(27106) <= 9497072;
srom_1(27107) <= 8925402;
srom_1(27108) <= 8351215;
srom_1(27109) <= 7777204;
srom_1(27110) <= 7206060;
srom_1(27111) <= 6640461;
srom_1(27112) <= 6083059;
srom_1(27113) <= 5536470;
srom_1(27114) <= 5003255;
srom_1(27115) <= 4485914;
srom_1(27116) <= 3986875;
srom_1(27117) <= 3508478;
srom_1(27118) <= 3052965;
srom_1(27119) <= 2622472;
srom_1(27120) <= 2219019;
srom_1(27121) <= 1844497;
srom_1(27122) <= 1500663;
srom_1(27123) <= 1189129;
srom_1(27124) <= 911355;
srom_1(27125) <= 668645;
srom_1(27126) <= 462136;
srom_1(27127) <= 292798;
srom_1(27128) <= 161423;
srom_1(27129) <= 68629;
srom_1(27130) <= 14850;
srom_1(27131) <= 338;
srom_1(27132) <= 25161;
srom_1(27133) <= 89204;
srom_1(27134) <= 192166;
srom_1(27135) <= 333563;
srom_1(27136) <= 512733;
srom_1(27137) <= 728836;
srom_1(27138) <= 980859;
srom_1(27139) <= 1267618;
srom_1(27140) <= 1587771;
srom_1(27141) <= 1939815;
srom_1(27142) <= 2322099;
srom_1(27143) <= 2732832;
srom_1(27144) <= 3170086;
srom_1(27145) <= 3631812;
srom_1(27146) <= 4115844;
srom_1(27147) <= 4619912;
srom_1(27148) <= 5141653;
srom_1(27149) <= 5678621;
srom_1(27150) <= 6228296;
srom_1(27151) <= 6788102;
srom_1(27152) <= 7355413;
srom_1(27153) <= 7927569;
srom_1(27154) <= 8501887;
srom_1(27155) <= 9075674;
srom_1(27156) <= 9646239;
srom_1(27157) <= 10210906;
srom_1(27158) <= 10767028;
srom_1(27159) <= 11311997;
srom_1(27160) <= 11843257;
srom_1(27161) <= 12358317;
srom_1(27162) <= 12854762;
srom_1(27163) <= 13330263;
srom_1(27164) <= 13782591;
srom_1(27165) <= 14209625;
srom_1(27166) <= 14609362;
srom_1(27167) <= 14979928;
srom_1(27168) <= 15319585;
srom_1(27169) <= 15626741;
srom_1(27170) <= 15899954;
srom_1(27171) <= 16137943;
srom_1(27172) <= 16339594;
srom_1(27173) <= 16503960;
srom_1(27174) <= 16630270;
srom_1(27175) <= 16717932;
srom_1(27176) <= 16766534;
srom_1(27177) <= 16775850;
srom_1(27178) <= 16745836;
srom_1(27179) <= 16676631;
srom_1(27180) <= 16568561;
srom_1(27181) <= 16422132;
srom_1(27182) <= 16238031;
srom_1(27183) <= 16017122;
srom_1(27184) <= 15760440;
srom_1(27185) <= 15469189;
srom_1(27186) <= 15144735;
srom_1(27187) <= 14788598;
srom_1(27188) <= 14402451;
srom_1(27189) <= 13988102;
srom_1(27190) <= 13547495;
srom_1(27191) <= 13082696;
srom_1(27192) <= 12595885;
srom_1(27193) <= 12089345;
srom_1(27194) <= 11565451;
srom_1(27195) <= 11026659;
srom_1(27196) <= 10475497;
srom_1(27197) <= 9914548;
srom_1(27198) <= 9346444;
srom_1(27199) <= 8773848;
srom_1(27200) <= 8199446;
srom_1(27201) <= 7625931;
srom_1(27202) <= 7055992;
srom_1(27203) <= 6492302;
srom_1(27204) <= 5937505;
srom_1(27205) <= 5394202;
srom_1(27206) <= 4864940;
srom_1(27207) <= 4352202;
srom_1(27208) <= 3858393;
srom_1(27209) <= 3385827;
srom_1(27210) <= 2936720;
srom_1(27211) <= 2513180;
srom_1(27212) <= 2117191;
srom_1(27213) <= 1750612;
srom_1(27214) <= 1415160;
srom_1(27215) <= 1112409;
srom_1(27216) <= 843778;
srom_1(27217) <= 610528;
srom_1(27218) <= 413752;
srom_1(27219) <= 254373;
srom_1(27220) <= 133138;
srom_1(27221) <= 50616;
srom_1(27222) <= 7193;
srom_1(27223) <= 3074;
srom_1(27224) <= 38277;
srom_1(27225) <= 112638;
srom_1(27226) <= 225808;
srom_1(27227) <= 377256;
srom_1(27228) <= 566272;
srom_1(27229) <= 791970;
srom_1(27230) <= 1053291;
srom_1(27231) <= 1349009;
srom_1(27232) <= 1677739;
srom_1(27233) <= 2037938;
srom_1(27234) <= 2427918;
srom_1(27235) <= 2845849;
srom_1(27236) <= 3289773;
srom_1(27237) <= 3757606;
srom_1(27238) <= 4247156;
srom_1(27239) <= 4756127;
srom_1(27240) <= 5282131;
srom_1(27241) <= 5822703;
srom_1(27242) <= 6375307;
srom_1(27243) <= 6937353;
srom_1(27244) <= 7506203;
srom_1(27245) <= 8079192;
srom_1(27246) <= 8653632;
srom_1(27247) <= 9226828;
srom_1(27248) <= 9796095;
srom_1(27249) <= 10358760;
srom_1(27250) <= 10912188;
srom_1(27251) <= 11453781;
srom_1(27252) <= 11981000;
srom_1(27253) <= 12491374;
srom_1(27254) <= 12982508;
srom_1(27255) <= 13452100;
srom_1(27256) <= 13897948;
srom_1(27257) <= 14317960;
srom_1(27258) <= 14710167;
srom_1(27259) <= 15072731;
srom_1(27260) <= 15403950;
srom_1(27261) <= 15702272;
srom_1(27262) <= 15966298;
srom_1(27263) <= 16194789;
srom_1(27264) <= 16386675;
srom_1(27265) <= 16541054;
srom_1(27266) <= 16657205;
srom_1(27267) <= 16734580;
srom_1(27268) <= 16772819;
srom_1(27269) <= 16771741;
srom_1(27270) <= 16731352;
srom_1(27271) <= 16651841;
srom_1(27272) <= 16533581;
srom_1(27273) <= 16377126;
srom_1(27274) <= 16183210;
srom_1(27275) <= 15952743;
srom_1(27276) <= 15686804;
srom_1(27277) <= 15386642;
srom_1(27278) <= 15053664;
srom_1(27279) <= 14689431;
srom_1(27280) <= 14295652;
srom_1(27281) <= 13874172;
srom_1(27282) <= 13426968;
srom_1(27283) <= 12956138;
srom_1(27284) <= 12463889;
srom_1(27285) <= 11952530;
srom_1(27286) <= 11424458;
srom_1(27287) <= 10882151;
srom_1(27288) <= 10328150;
srom_1(27289) <= 9765054;
srom_1(27290) <= 9195503;
srom_1(27291) <= 8622168;
srom_1(27292) <= 8047738;
srom_1(27293) <= 7474907;
srom_1(27294) <= 6906360;
srom_1(27295) <= 6344764;
srom_1(27296) <= 5792753;
srom_1(27297) <= 5252914;
srom_1(27298) <= 4727779;
srom_1(27299) <= 4219812;
srom_1(27300) <= 3731393;
srom_1(27301) <= 3264814;
srom_1(27302) <= 2822261;
srom_1(27303) <= 2405812;
srom_1(27304) <= 2017417;
srom_1(27305) <= 1658900;
srom_1(27306) <= 1331940;
srom_1(27307) <= 1038071;
srom_1(27308) <= 778672;
srom_1(27309) <= 554958;
srom_1(27310) <= 367979;
srom_1(27311) <= 218611;
srom_1(27312) <= 107556;
srom_1(27313) <= 35333;
srom_1(27314) <= 2281;
srom_1(27315) <= 8556;
srom_1(27316) <= 54127;
srom_1(27317) <= 138782;
srom_1(27318) <= 262123;
srom_1(27319) <= 423572;
srom_1(27320) <= 622372;
srom_1(27321) <= 857590;
srom_1(27322) <= 1128124;
srom_1(27323) <= 1432705;
srom_1(27324) <= 1769904;
srom_1(27325) <= 2138141;
srom_1(27326) <= 2535688;
srom_1(27327) <= 2960682;
srom_1(27328) <= 3411129;
srom_1(27329) <= 3884917;
srom_1(27330) <= 4379825;
srom_1(27331) <= 4893531;
srom_1(27332) <= 5423626;
srom_1(27333) <= 5967626;
srom_1(27334) <= 6522978;
srom_1(27335) <= 7087079;
srom_1(27336) <= 7657283;
srom_1(27337) <= 8230917;
srom_1(27338) <= 8805290;
srom_1(27339) <= 9377709;
srom_1(27340) <= 9945490;
srom_1(27341) <= 10505970;
srom_1(27342) <= 11056521;
srom_1(27343) <= 11594561;
srom_1(27344) <= 12117567;
srom_1(27345) <= 12623088;
srom_1(27346) <= 13108751;
srom_1(27347) <= 13572279;
srom_1(27348) <= 14011500;
srom_1(27349) <= 14424353;
srom_1(27350) <= 14808903;
srom_1(27351) <= 15163345;
srom_1(27352) <= 15486018;
srom_1(27353) <= 15775409;
srom_1(27354) <= 16030161;
srom_1(27355) <= 16249079;
srom_1(27356) <= 16431137;
srom_1(27357) <= 16575480;
srom_1(27358) <= 16681432;
srom_1(27359) <= 16748497;
srom_1(27360) <= 16776359;
srom_1(27361) <= 16764888;
srom_1(27362) <= 16714137;
srom_1(27363) <= 16624346;
srom_1(27364) <= 16495934;
srom_1(27365) <= 16329504;
srom_1(27366) <= 16125837;
srom_1(27367) <= 15885887;
srom_1(27368) <= 15610779;
srom_1(27369) <= 15301805;
srom_1(27370) <= 14960412;
srom_1(27371) <= 14588201;
srom_1(27372) <= 14186919;
srom_1(27373) <= 13758446;
srom_1(27374) <= 13304792;
srom_1(27375) <= 12828085;
srom_1(27376) <= 12330559;
srom_1(27377) <= 11814549;
srom_1(27378) <= 11282472;
srom_1(27379) <= 10736826;
srom_1(27380) <= 10180168;
srom_1(27381) <= 9615108;
srom_1(27382) <= 9044297;
srom_1(27383) <= 8470412;
srom_1(27384) <= 7896142;
srom_1(27385) <= 7324182;
srom_1(27386) <= 6757214;
srom_1(27387) <= 6197896;
srom_1(27388) <= 5648850;
srom_1(27389) <= 5112653;
srom_1(27390) <= 4591817;
srom_1(27391) <= 4088786;
srom_1(27392) <= 3605918;
srom_1(27393) <= 3145478;
srom_1(27394) <= 2709625;
srom_1(27395) <= 2300402;
srom_1(27396) <= 1919729;
srom_1(27397) <= 1569391;
srom_1(27398) <= 1251030;
srom_1(27399) <= 966140;
srom_1(27400) <= 716057;
srom_1(27401) <= 501953;
srom_1(27402) <= 324832;
srom_1(27403) <= 185524;
srom_1(27404) <= 84684;
srom_1(27405) <= 22784;
srom_1(27406) <= 114;
srom_1(27407) <= 16781;
srom_1(27408) <= 72706;
srom_1(27409) <= 167627;
srom_1(27410) <= 301099;
srom_1(27411) <= 472496;
srom_1(27412) <= 681014;
srom_1(27413) <= 925676;
srom_1(27414) <= 1205335;
srom_1(27415) <= 1518678;
srom_1(27416) <= 1864236;
srom_1(27417) <= 2240390;
srom_1(27418) <= 2645375;
srom_1(27419) <= 3077291;
srom_1(27420) <= 3534115;
srom_1(27421) <= 4013702;
srom_1(27422) <= 4513805;
srom_1(27423) <= 5032079;
srom_1(27424) <= 5566092;
srom_1(27425) <= 6113341;
srom_1(27426) <= 6671259;
srom_1(27427) <= 7237231;
srom_1(27428) <= 7808602;
srom_1(27429) <= 8382693;
srom_1(27430) <= 8956811;
srom_1(27431) <= 9528265;
srom_1(27432) <= 10094375;
srom_1(27433) <= 10652486;
srom_1(27434) <= 11199980;
srom_1(27435) <= 11734292;
srom_1(27436) <= 12252914;
srom_1(27437) <= 12753415;
srom_1(27438) <= 13233448;
srom_1(27439) <= 13690762;
srom_1(27440) <= 14123212;
srom_1(27441) <= 14528771;
srom_1(27442) <= 14905536;
srom_1(27443) <= 15251741;
srom_1(27444) <= 15565763;
srom_1(27445) <= 15846128;
srom_1(27446) <= 16091523;
srom_1(27447) <= 16300796;
srom_1(27448) <= 16472966;
srom_1(27449) <= 16607226;
srom_1(27450) <= 16702945;
srom_1(27451) <= 16759676;
srom_1(27452) <= 16777152;
srom_1(27453) <= 16755292;
srom_1(27454) <= 16694197;
srom_1(27455) <= 16594154;
srom_1(27456) <= 16455633;
srom_1(27457) <= 16279282;
srom_1(27458) <= 16065930;
srom_1(27459) <= 15816576;
srom_1(27460) <= 15532390;
srom_1(27461) <= 15214704;
srom_1(27462) <= 14865008;
srom_1(27463) <= 14484942;
srom_1(27464) <= 14076288;
srom_1(27465) <= 13640962;
srom_1(27466) <= 13181007;
srom_1(27467) <= 12698578;
srom_1(27468) <= 12195939;
srom_1(27469) <= 11675445;
srom_1(27470) <= 11139539;
srom_1(27471) <= 10590732;
srom_1(27472) <= 10031599;
srom_1(27473) <= 9464761;
srom_1(27474) <= 8892877;
srom_1(27475) <= 8318628;
srom_1(27476) <= 7744708;
srom_1(27477) <= 7173806;
srom_1(27478) <= 6608602;
srom_1(27479) <= 6051744;
srom_1(27480) <= 5505845;
srom_1(27481) <= 4973464;
srom_1(27482) <= 4457098;
srom_1(27483) <= 3959168;
srom_1(27484) <= 3482009;
srom_1(27485) <= 3027859;
srom_1(27486) <= 2598847;
srom_1(27487) <= 2196985;
srom_1(27488) <= 1824159;
srom_1(27489) <= 1482115;
srom_1(27490) <= 1172457;
srom_1(27491) <= 896639;
srom_1(27492) <= 655954;
srom_1(27493) <= 451529;
srom_1(27494) <= 284324;
srom_1(27495) <= 155123;
srom_1(27496) <= 64532;
srom_1(27497) <= 12975;
srom_1(27498) <= 694;
srom_1(27499) <= 27747;
srom_1(27500) <= 94007;
srom_1(27501) <= 199163;
srom_1(27502) <= 342722;
srom_1(27503) <= 524011;
srom_1(27504) <= 742180;
srom_1(27505) <= 996206;
srom_1(27506) <= 1284897;
srom_1(27507) <= 1606900;
srom_1(27508) <= 1960705;
srom_1(27509) <= 2344652;
srom_1(27510) <= 2756941;
srom_1(27511) <= 3195640;
srom_1(27512) <= 3658690;
srom_1(27513) <= 4143920;
srom_1(27514) <= 4649055;
srom_1(27515) <= 5171726;
srom_1(27516) <= 5709482;
srom_1(27517) <= 6259801;
srom_1(27518) <= 6820103;
srom_1(27519) <= 7387760;
srom_1(27520) <= 7960111;
srom_1(27521) <= 8534471;
srom_1(27522) <= 9108147;
srom_1(27523) <= 9678449;
srom_1(27524) <= 10242702;
srom_1(27525) <= 10798261;
srom_1(27526) <= 11342520;
srom_1(27527) <= 11872927;
srom_1(27528) <= 12386995;
srom_1(27529) <= 12882313;
srom_1(27530) <= 13356559;
srom_1(27531) <= 13807508;
srom_1(27532) <= 14233046;
srom_1(27533) <= 14631178;
srom_1(27534) <= 15000036;
srom_1(27535) <= 15337890;
srom_1(27536) <= 15643158;
srom_1(27537) <= 15914406;
srom_1(27538) <= 16150363;
srom_1(27539) <= 16349922;
srom_1(27540) <= 16512148;
srom_1(27541) <= 16636280;
srom_1(27542) <= 16721736;
srom_1(27543) <= 16768115;
srom_1(27544) <= 16775200;
srom_1(27545) <= 16742957;
srom_1(27546) <= 16671537;
srom_1(27547) <= 16561276;
srom_1(27548) <= 16412691;
srom_1(27549) <= 16226478;
srom_1(27550) <= 16003510;
srom_1(27551) <= 15744833;
srom_1(27552) <= 15451661;
srom_1(27553) <= 15125368;
srom_1(27554) <= 14767483;
srom_1(27555) <= 14379686;
srom_1(27556) <= 13963795;
srom_1(27557) <= 13521759;
srom_1(27558) <= 13055653;
srom_1(27559) <= 12567661;
srom_1(27560) <= 12060072;
srom_1(27561) <= 11535266;
srom_1(27562) <= 10995705;
srom_1(27563) <= 10443918;
srom_1(27564) <= 9882493;
srom_1(27565) <= 9314062;
srom_1(27566) <= 8741292;
srom_1(27567) <= 8166868;
srom_1(27568) <= 7593484;
srom_1(27569) <= 7023828;
srom_1(27570) <= 6460572;
srom_1(27571) <= 5906358;
srom_1(27572) <= 5363783;
srom_1(27573) <= 4835393;
srom_1(27574) <= 4323666;
srom_1(27575) <= 3831000;
srom_1(27576) <= 3359706;
srom_1(27577) <= 2911995;
srom_1(27578) <= 2489965;
srom_1(27579) <= 2095596;
srom_1(27580) <= 1730737;
srom_1(27581) <= 1397099;
srom_1(27582) <= 1096247;
srom_1(27583) <= 829591;
srom_1(27584) <= 598382;
srom_1(27585) <= 403704;
srom_1(27586) <= 246470;
srom_1(27587) <= 127417;
srom_1(27588) <= 47104;
srom_1(27589) <= 5907;
srom_1(27590) <= 4019;
srom_1(27591) <= 41450;
srom_1(27592) <= 118023;
srom_1(27593) <= 233380;
srom_1(27594) <= 386979;
srom_1(27595) <= 578101;
srom_1(27596) <= 805849;
srom_1(27597) <= 1069155;
srom_1(27598) <= 1366785;
srom_1(27599) <= 1697342;
srom_1(27600) <= 2059277;
srom_1(27601) <= 2450893;
srom_1(27602) <= 2870352;
srom_1(27603) <= 3315688;
srom_1(27604) <= 3784813;
srom_1(27605) <= 4275527;
srom_1(27606) <= 4785528;
srom_1(27607) <= 5312426;
srom_1(27608) <= 5853748;
srom_1(27609) <= 6406958;
srom_1(27610) <= 6969460;
srom_1(27611) <= 7538617;
srom_1(27612) <= 8111760;
srom_1(27613) <= 8686201;
srom_1(27614) <= 9259247;
srom_1(27615) <= 9828210;
srom_1(27616) <= 10390422;
srom_1(27617) <= 10943247;
srom_1(27618) <= 11484092;
srom_1(27619) <= 12010422;
srom_1(27620) <= 12519767;
srom_1(27621) <= 13009740;
srom_1(27622) <= 13478043;
srom_1(27623) <= 13922480;
srom_1(27624) <= 14340967;
srom_1(27625) <= 14731541;
srom_1(27626) <= 15092371;
srom_1(27627) <= 15421765;
srom_1(27628) <= 15718177;
srom_1(27629) <= 15980219;
srom_1(27630) <= 16206661;
srom_1(27631) <= 16396442;
srom_1(27632) <= 16548671;
srom_1(27633) <= 16662635;
srom_1(27634) <= 16737799;
srom_1(27635) <= 16773810;
srom_1(27636) <= 16770501;
srom_1(27637) <= 16727886;
srom_1(27638) <= 16646166;
srom_1(27639) <= 16525722;
srom_1(27640) <= 16367121;
srom_1(27641) <= 16171107;
srom_1(27642) <= 15938597;
srom_1(27643) <= 15670683;
srom_1(27644) <= 15368620;
srom_1(27645) <= 15033826;
srom_1(27646) <= 14667870;
srom_1(27647) <= 14272469;
srom_1(27648) <= 13849476;
srom_1(27649) <= 13400875;
srom_1(27650) <= 12928770;
srom_1(27651) <= 12435375;
srom_1(27652) <= 11923003;
srom_1(27653) <= 11394057;
srom_1(27654) <= 10851017;
srom_1(27655) <= 10296430;
srom_1(27656) <= 9732897;
srom_1(27657) <= 9163060;
srom_1(27658) <= 8589591;
srom_1(27659) <= 8015180;
srom_1(27660) <= 7442520;
srom_1(27661) <= 6874296;
srom_1(27662) <= 6313174;
srom_1(27663) <= 5761784;
srom_1(27664) <= 5222712;
srom_1(27665) <= 4698486;
srom_1(27666) <= 4191564;
srom_1(27667) <= 3704324;
srom_1(27668) <= 3239050;
srom_1(27669) <= 2797924;
srom_1(27670) <= 2383014;
srom_1(27671) <= 1996267;
srom_1(27672) <= 1639496;
srom_1(27673) <= 1314373;
srom_1(27674) <= 1022424;
srom_1(27675) <= 765018;
srom_1(27676) <= 543361;
srom_1(27677) <= 358494;
srom_1(27678) <= 211282;
srom_1(27679) <= 102416;
srom_1(27680) <= 32408;
srom_1(27681) <= 1584;
srom_1(27682) <= 10090;
srom_1(27683) <= 57886;
srom_1(27684) <= 144748;
srom_1(27685) <= 270267;
srom_1(27686) <= 433857;
srom_1(27687) <= 634749;
srom_1(27688) <= 872001;
srom_1(27689) <= 1144501;
srom_1(27690) <= 1450972;
srom_1(27691) <= 1789975;
srom_1(27692) <= 2159922;
srom_1(27693) <= 2559077;
srom_1(27694) <= 2985569;
srom_1(27695) <= 3437397;
srom_1(27696) <= 3912444;
srom_1(27697) <= 4408481;
srom_1(27698) <= 4923181;
srom_1(27699) <= 5454133;
srom_1(27700) <= 5998845;
srom_1(27701) <= 6554764;
srom_1(27702) <= 7119282;
srom_1(27703) <= 7689752;
srom_1(27704) <= 8263500;
srom_1(27705) <= 8837834;
srom_1(27706) <= 9410062;
srom_1(27707) <= 9977499;
srom_1(27708) <= 10537486;
srom_1(27709) <= 11087396;
srom_1(27710) <= 11624651;
srom_1(27711) <= 12146730;
srom_1(27712) <= 12651187;
srom_1(27713) <= 13135654;
srom_1(27714) <= 13597862;
srom_1(27715) <= 14035641;
srom_1(27716) <= 14446939;
srom_1(27717) <= 14829828;
srom_1(27718) <= 15182511;
srom_1(27719) <= 15503336;
srom_1(27720) <= 15790797;
srom_1(27721) <= 16043547;
srom_1(27722) <= 16260400;
srom_1(27723) <= 16440340;
srom_1(27724) <= 16582522;
srom_1(27725) <= 16686280;
srom_1(27726) <= 16751128;
srom_1(27727) <= 16776761;
srom_1(27728) <= 16763059;
srom_1(27729) <= 16710086;
srom_1(27730) <= 16618091;
srom_1(27731) <= 16487505;
srom_1(27732) <= 16318940;
srom_1(27733) <= 16113188;
srom_1(27734) <= 15871212;
srom_1(27735) <= 15594148;
srom_1(27736) <= 15283294;
srom_1(27737) <= 14940109;
srom_1(27738) <= 14566202;
srom_1(27739) <= 14163326;
srom_1(27740) <= 13733370;
srom_1(27741) <= 13278350;
srom_1(27742) <= 12800402;
srom_1(27743) <= 12301764;
srom_1(27744) <= 11784777;
srom_1(27745) <= 11251863;
srom_1(27746) <= 10705523;
srom_1(27747) <= 10148318;
srom_1(27748) <= 9582861;
srom_1(27749) <= 9011804;
srom_1(27750) <= 8437825;
srom_1(27751) <= 7863615;
srom_1(27752) <= 7291866;
srom_1(27753) <= 6725261;
srom_1(27754) <= 6166455;
srom_1(27755) <= 5618070;
srom_1(27756) <= 5082677;
srom_1(27757) <= 4562787;
srom_1(27758) <= 4060837;
srom_1(27759) <= 3579182;
srom_1(27760) <= 3120079;
srom_1(27761) <= 2685683;
srom_1(27762) <= 2278030;
srom_1(27763) <= 1899031;
srom_1(27764) <= 1550464;
srom_1(27765) <= 1233963;
srom_1(27766) <= 951013;
srom_1(27767) <= 702941;
srom_1(27768) <= 490909;
srom_1(27769) <= 315912;
srom_1(27770) <= 178771;
srom_1(27771) <= 80128;
srom_1(27772) <= 20447;
srom_1(27773) <= 7;
srom_1(27774) <= 18904;
srom_1(27775) <= 77050;
srom_1(27776) <= 174171;
srom_1(27777) <= 309812;
srom_1(27778) <= 483338;
srom_1(27779) <= 693934;
srom_1(27780) <= 940614;
srom_1(27781) <= 1222219;
srom_1(27782) <= 1537430;
srom_1(27783) <= 1884769;
srom_1(27784) <= 2262606;
srom_1(27785) <= 2669170;
srom_1(27786) <= 3102555;
srom_1(27787) <= 3560728;
srom_1(27788) <= 4041540;
srom_1(27789) <= 4542737;
srom_1(27790) <= 5061969;
srom_1(27791) <= 5596801;
srom_1(27792) <= 6144724;
srom_1(27793) <= 6703170;
srom_1(27794) <= 7269519;
srom_1(27795) <= 7841116;
srom_1(27796) <= 8415281;
srom_1(27797) <= 8989320;
srom_1(27798) <= 9560542;
srom_1(27799) <= 10126269;
srom_1(27800) <= 10683847;
srom_1(27801) <= 11230662;
srom_1(27802) <= 11764150;
srom_1(27803) <= 12281809;
srom_1(27804) <= 12781211;
srom_1(27805) <= 13260014;
srom_1(27806) <= 13715974;
srom_1(27807) <= 14146952;
srom_1(27808) <= 14550928;
srom_1(27809) <= 14926006;
srom_1(27810) <= 15270428;
srom_1(27811) <= 15582578;
srom_1(27812) <= 15860994;
srom_1(27813) <= 16104369;
srom_1(27814) <= 16311562;
srom_1(27815) <= 16481602;
srom_1(27816) <= 16613691;
srom_1(27817) <= 16707209;
srom_1(27818) <= 16761719;
srom_1(27819) <= 16776965;
srom_1(27820) <= 16752874;
srom_1(27821) <= 16689561;
srom_1(27822) <= 16587321;
srom_1(27823) <= 16446635;
srom_1(27824) <= 16268163;
srom_1(27825) <= 16052740;
srom_1(27826) <= 15801377;
srom_1(27827) <= 15515254;
srom_1(27828) <= 15195711;
srom_1(27829) <= 14844247;
srom_1(27830) <= 14462511;
srom_1(27831) <= 14052292;
srom_1(27832) <= 13615514;
srom_1(27833) <= 13154225;
srom_1(27834) <= 12670588;
srom_1(27835) <= 12166872;
srom_1(27836) <= 11645439;
srom_1(27837) <= 11108732;
srom_1(27838) <= 10559271;
srom_1(27839) <= 9999630;
srom_1(27840) <= 9432435;
srom_1(27841) <= 8860345;
srom_1(27842) <= 8286042;
srom_1(27843) <= 7712221;
srom_1(27844) <= 7141571;
srom_1(27845) <= 6576769;
srom_1(27846) <= 6020464;
srom_1(27847) <= 5475264;
srom_1(27848) <= 4943725;
srom_1(27849) <= 4428340;
srom_1(27850) <= 3931527;
srom_1(27851) <= 3455614;
srom_1(27852) <= 3002834;
srom_1(27853) <= 2575309;
srom_1(27854) <= 2175045;
srom_1(27855) <= 1803919;
srom_1(27856) <= 1463671;
srom_1(27857) <= 1155895;
srom_1(27858) <= 882037;
srom_1(27859) <= 643379;
srom_1(27860) <= 441042;
srom_1(27861) <= 275973;
srom_1(27862) <= 148947;
srom_1(27863) <= 60560;
srom_1(27864) <= 11226;
srom_1(27865) <= 1176;
srom_1(27866) <= 30458;
srom_1(27867) <= 98934;
srom_1(27868) <= 206283;
srom_1(27869) <= 352002;
srom_1(27870) <= 535408;
srom_1(27871) <= 755639;
srom_1(27872) <= 1011665;
srom_1(27873) <= 1302283;
srom_1(27874) <= 1626131;
srom_1(27875) <= 1981691;
srom_1(27876) <= 2367296;
srom_1(27877) <= 2781136;
srom_1(27878) <= 3221272;
srom_1(27879) <= 3685639;
srom_1(27880) <= 4172060;
srom_1(27881) <= 4678253;
srom_1(27882) <= 5201846;
srom_1(27883) <= 5740383;
srom_1(27884) <= 6291338;
srom_1(27885) <= 6852128;
srom_1(27886) <= 7420123;
srom_1(27887) <= 7992659;
srom_1(27888) <= 8567053;
srom_1(27889) <= 9140609;
srom_1(27890) <= 9710639;
srom_1(27891) <= 10274470;
srom_1(27892) <= 10829457;
srom_1(27893) <= 11372998;
srom_1(27894) <= 11902544;
srom_1(27895) <= 12415613;
srom_1(27896) <= 12909797;
srom_1(27897) <= 13382780;
srom_1(27898) <= 13832343;
srom_1(27899) <= 14256379;
srom_1(27900) <= 14652899;
srom_1(27901) <= 15020043;
srom_1(27902) <= 15356091;
srom_1(27903) <= 15659465;
srom_1(27904) <= 15928744;
srom_1(27905) <= 16162665;
srom_1(27906) <= 16360130;
srom_1(27907) <= 16520214;
srom_1(27908) <= 16642166;
srom_1(27909) <= 16725415;
srom_1(27910) <= 16769569;
srom_1(27911) <= 16774422;
srom_1(27912) <= 16739951;
srom_1(27913) <= 16666318;
srom_1(27914) <= 16553868;
srom_1(27915) <= 16403128;
srom_1(27916) <= 16214805;
srom_1(27917) <= 15989783;
srom_1(27918) <= 15729116;
srom_1(27919) <= 15434026;
srom_1(27920) <= 15105899;
srom_1(27921) <= 14746272;
srom_1(27922) <= 14356831;
srom_1(27923) <= 13939403;
srom_1(27924) <= 13495946;
srom_1(27925) <= 13028539;
srom_1(27926) <= 12539373;
srom_1(27927) <= 12030743;
srom_1(27928) <= 11505034;
srom_1(27929) <= 10964711;
srom_1(27930) <= 10412308;
srom_1(27931) <= 9850415;
srom_1(27932) <= 9281666;
srom_1(27933) <= 8708730;
srom_1(27934) <= 8134293;
srom_1(27935) <= 7561049;
srom_1(27936) <= 6991685;
srom_1(27937) <= 6428871;
srom_1(27938) <= 5875248;
srom_1(27939) <= 5333411;
srom_1(27940) <= 4805900;
srom_1(27941) <= 4295190;
srom_1(27942) <= 3803676;
srom_1(27943) <= 3333661;
srom_1(27944) <= 2887352;
srom_1(27945) <= 2466839;
srom_1(27946) <= 2074096;
srom_1(27947) <= 1710963;
srom_1(27948) <= 1379144;
srom_1(27949) <= 1080196;
srom_1(27950) <= 815518;
srom_1(27951) <= 586354;
srom_1(27952) <= 393777;
srom_1(27953) <= 238690;
srom_1(27954) <= 121822;
srom_1(27955) <= 43719;
srom_1(27956) <= 4748;
srom_1(27957) <= 5092;
srom_1(27958) <= 44749;
srom_1(27959) <= 123533;
srom_1(27960) <= 241075;
srom_1(27961) <= 396824;
srom_1(27962) <= 590048;
srom_1(27963) <= 819843;
srom_1(27964) <= 1085131;
srom_1(27965) <= 1384667;
srom_1(27966) <= 1717047;
srom_1(27967) <= 2080712;
srom_1(27968) <= 2473957;
srom_1(27969) <= 2894938;
srom_1(27970) <= 3341680;
srom_1(27971) <= 3812089;
srom_1(27972) <= 4303960;
srom_1(27973) <= 4814984;
srom_1(27974) <= 5342766;
srom_1(27975) <= 5884832;
srom_1(27976) <= 6438638;
srom_1(27977) <= 7001589;
srom_1(27978) <= 7571044;
srom_1(27979) <= 8144332;
srom_1(27980) <= 8718766;
srom_1(27981) <= 9291652;
srom_1(27982) <= 9860303;
srom_1(27983) <= 10422053;
srom_1(27984) <= 10974267;
srom_1(27985) <= 11514357;
srom_1(27986) <= 12039788;
srom_1(27987) <= 12548098;
srom_1(27988) <= 13036903;
srom_1(27989) <= 13503910;
srom_1(27990) <= 13946929;
srom_1(27991) <= 14363884;
srom_1(27992) <= 14752819;
srom_1(27993) <= 15111910;
srom_1(27994) <= 15439473;
srom_1(27995) <= 15733972;
srom_1(27996) <= 15994026;
srom_1(27997) <= 16218415;
srom_1(27998) <= 16406088;
srom_1(27999) <= 16556164;
srom_1(28000) <= 16667940;
srom_1(28001) <= 16740891;
srom_1(28002) <= 16774675;
srom_1(28003) <= 16769135;
srom_1(28004) <= 16724294;
srom_1(28005) <= 16640366;
srom_1(28006) <= 16517741;
srom_1(28007) <= 16356997;
srom_1(28008) <= 16158886;
srom_1(28009) <= 15924337;
srom_1(28010) <= 15654451;
srom_1(28011) <= 15350493;
srom_1(28012) <= 15013888;
srom_1(28013) <= 14646215;
srom_1(28014) <= 14249197;
srom_1(28015) <= 13824698;
srom_1(28016) <= 13374707;
srom_1(28017) <= 12901334;
srom_1(28018) <= 12406799;
srom_1(28019) <= 11893422;
srom_1(28020) <= 11363610;
srom_1(28021) <= 10819846;
srom_1(28022) <= 10264682;
srom_1(28023) <= 9700720;
srom_1(28024) <= 9130606;
srom_1(28025) <= 8557011;
srom_1(28026) <= 7982627;
srom_1(28027) <= 7410147;
srom_1(28028) <= 6842256;
srom_1(28029) <= 6281615;
srom_1(28030) <= 5730855;
srom_1(28031) <= 5192558;
srom_1(28032) <= 4669249;
srom_1(28033) <= 4163380;
srom_1(28034) <= 3677326;
srom_1(28035) <= 3213364;
srom_1(28036) <= 2773670;
srom_1(28037) <= 2360307;
srom_1(28038) <= 1975213;
srom_1(28039) <= 1620194;
srom_1(28040) <= 1296913;
srom_1(28041) <= 1006888;
srom_1(28042) <= 751479;
srom_1(28043) <= 531883;
srom_1(28044) <= 349129;
srom_1(28045) <= 204076;
srom_1(28046) <= 97402;
srom_1(28047) <= 29609;
srom_1(28048) <= 1014;
srom_1(28049) <= 11751;
srom_1(28050) <= 61771;
srom_1(28051) <= 150837;
srom_1(28052) <= 278534;
srom_1(28053) <= 444261;
srom_1(28054) <= 647242;
srom_1(28055) <= 886525;
srom_1(28056) <= 1160988;
srom_1(28057) <= 1469344;
srom_1(28058) <= 1810146;
srom_1(28059) <= 2181797;
srom_1(28060) <= 2582554;
srom_1(28061) <= 3010538;
srom_1(28062) <= 3463741;
srom_1(28063) <= 3940038;
srom_1(28064) <= 4437197;
srom_1(28065) <= 4952885;
srom_1(28066) <= 5484684;
srom_1(28067) <= 6030101;
srom_1(28068) <= 6586577;
srom_1(28069) <= 7151504;
srom_1(28070) <= 7722232;
srom_1(28071) <= 8296085;
srom_1(28072) <= 8870372;
srom_1(28073) <= 9442399;
srom_1(28074) <= 10009485;
srom_1(28075) <= 10568970;
srom_1(28076) <= 11118231;
srom_1(28077) <= 11654692;
srom_1(28078) <= 12175836;
srom_1(28079) <= 12679222;
srom_1(28080) <= 13162487;
srom_1(28081) <= 13623365;
srom_1(28082) <= 14059696;
srom_1(28083) <= 14469433;
srom_1(28084) <= 14850656;
srom_1(28085) <= 15201575;
srom_1(28086) <= 15520546;
srom_1(28087) <= 15806073;
srom_1(28088) <= 16056817;
srom_1(28089) <= 16271602;
srom_1(28090) <= 16449421;
srom_1(28091) <= 16589440;
srom_1(28092) <= 16691003;
srom_1(28093) <= 16753633;
srom_1(28094) <= 16777036;
srom_1(28095) <= 16761103;
srom_1(28096) <= 16705909;
srom_1(28097) <= 16611711;
srom_1(28098) <= 16478953;
srom_1(28099) <= 16308257;
srom_1(28100) <= 16100422;
srom_1(28101) <= 15856424;
srom_1(28102) <= 15577407;
srom_1(28103) <= 15264680;
srom_1(28104) <= 14919708;
srom_1(28105) <= 14544109;
srom_1(28106) <= 14139645;
srom_1(28107) <= 13708213;
srom_1(28108) <= 13251835;
srom_1(28109) <= 12772651;
srom_1(28110) <= 12272910;
srom_1(28111) <= 11754953;
srom_1(28112) <= 11221211;
srom_1(28113) <= 10674186;
srom_1(28114) <= 10116442;
srom_1(28115) <= 9550597;
srom_1(28116) <= 8979302;
srom_1(28117) <= 8405237;
srom_1(28118) <= 7831095;
srom_1(28119) <= 7259566;
srom_1(28120) <= 6693333;
srom_1(28121) <= 6135048;
srom_1(28122) <= 5587332;
srom_1(28123) <= 5052752;
srom_1(28124) <= 4533815;
srom_1(28125) <= 4032954;
srom_1(28126) <= 3552518;
srom_1(28127) <= 3094760;
srom_1(28128) <= 2661827;
srom_1(28129) <= 2255749;
srom_1(28130) <= 1878430;
srom_1(28131) <= 1531640;
srom_1(28132) <= 1217004;
srom_1(28133) <= 935998;
srom_1(28134) <= 689940;
srom_1(28135) <= 479984;
srom_1(28136) <= 307114;
srom_1(28137) <= 172141;
srom_1(28138) <= 75697;
srom_1(28139) <= 18236;
srom_1(28140) <= 27;
srom_1(28141) <= 21154;
srom_1(28142) <= 81519;
srom_1(28143) <= 180839;
srom_1(28144) <= 318648;
srom_1(28145) <= 494300;
srom_1(28146) <= 706971;
srom_1(28147) <= 955663;
srom_1(28148) <= 1239212;
srom_1(28149) <= 1556286;
srom_1(28150) <= 1905399;
srom_1(28151) <= 2284915;
srom_1(28152) <= 2693052;
srom_1(28153) <= 3127899;
srom_1(28154) <= 3587414;
srom_1(28155) <= 4069444;
srom_1(28156) <= 4571728;
srom_1(28157) <= 5091910;
srom_1(28158) <= 5627552;
srom_1(28159) <= 6176141;
srom_1(28160) <= 6735106;
srom_1(28161) <= 7301824;
srom_1(28162) <= 7873639;
srom_1(28163) <= 8447868;
srom_1(28164) <= 9021819;
srom_1(28165) <= 9592802;
srom_1(28166) <= 10158137;
srom_1(28167) <= 10715174;
srom_1(28168) <= 11261301;
srom_1(28169) <= 11793958;
srom_1(28170) <= 12310645;
srom_1(28171) <= 12808940;
srom_1(28172) <= 13286508;
srom_1(28173) <= 13741107;
srom_1(28174) <= 14170606;
srom_1(28175) <= 14572992;
srom_1(28176) <= 14946377;
srom_1(28177) <= 15289010;
srom_1(28178) <= 15599285;
srom_1(28179) <= 15875747;
srom_1(28180) <= 16117098;
srom_1(28181) <= 16322209;
srom_1(28182) <= 16490116;
srom_1(28183) <= 16620032;
srom_1(28184) <= 16711348;
srom_1(28185) <= 16763636;
srom_1(28186) <= 16776650;
srom_1(28187) <= 16750330;
srom_1(28188) <= 16684800;
srom_1(28189) <= 16580365;
srom_1(28190) <= 16437516;
srom_1(28191) <= 16256924;
srom_1(28192) <= 16039434;
srom_1(28193) <= 15786067;
srom_1(28194) <= 15498010;
srom_1(28195) <= 15176615;
srom_1(28196) <= 14823389;
srom_1(28197) <= 14439988;
srom_1(28198) <= 14028210;
srom_1(28199) <= 13589986;
srom_1(28200) <= 13127371;
srom_1(28201) <= 12642534;
srom_1(28202) <= 12137749;
srom_1(28203) <= 11615383;
srom_1(28204) <= 11077885;
srom_1(28205) <= 10527777;
srom_1(28206) <= 9967637;
srom_1(28207) <= 9400092;
srom_1(28208) <= 8827805;
srom_1(28209) <= 8253458;
srom_1(28210) <= 7679744;
srom_1(28211) <= 7109355;
srom_1(28212) <= 6544965;
srom_1(28213) <= 5989220;
srom_1(28214) <= 5444726;
srom_1(28215) <= 4914038;
srom_1(28216) <= 4399643;
srom_1(28217) <= 3903953;
srom_1(28218) <= 3429294;
srom_1(28219) <= 2977890;
srom_1(28220) <= 2551859;
srom_1(28221) <= 2153199;
srom_1(28222) <= 1783779;
srom_1(28223) <= 1445331;
srom_1(28224) <= 1139442;
srom_1(28225) <= 867548;
srom_1(28226) <= 630922;
srom_1(28227) <= 430674;
srom_1(28228) <= 267744;
srom_1(28229) <= 142896;
srom_1(28230) <= 56714;
srom_1(28231) <= 9604;
srom_1(28232) <= 1785;
srom_1(28233) <= 33296;
srom_1(28234) <= 103987;
srom_1(28235) <= 213528;
srom_1(28236) <= 361404;
srom_1(28237) <= 546923;
srom_1(28238) <= 769214;
srom_1(28239) <= 1027235;
srom_1(28240) <= 1319776;
srom_1(28241) <= 1645465;
srom_1(28242) <= 2002775;
srom_1(28243) <= 2390031;
srom_1(28244) <= 2805415;
srom_1(28245) <= 3246982;
srom_1(28246) <= 3712659;
srom_1(28247) <= 4200263;
srom_1(28248) <= 4707508;
srom_1(28249) <= 5232015;
srom_1(28250) <= 5771324;
srom_1(28251) <= 6322907;
srom_1(28252) <= 6884176;
srom_1(28253) <= 7452500;
srom_1(28254) <= 8025214;
srom_1(28255) <= 8599632;
srom_1(28256) <= 9173060;
srom_1(28257) <= 9742810;
srom_1(28258) <= 10306209;
srom_1(28259) <= 10860616;
srom_1(28260) <= 11403431;
srom_1(28261) <= 11932109;
srom_1(28262) <= 12444169;
srom_1(28263) <= 12937212;
srom_1(28264) <= 13408925;
srom_1(28265) <= 13857096;
srom_1(28266) <= 14279623;
srom_1(28267) <= 14674525;
srom_1(28268) <= 15039951;
srom_1(28269) <= 15374186;
srom_1(28270) <= 15675663;
srom_1(28271) <= 15942969;
srom_1(28272) <= 16174849;
srom_1(28273) <= 16370218;
srom_1(28274) <= 16528157;
srom_1(28275) <= 16647928;
srom_1(28276) <= 16728968;
srom_1(28277) <= 16770897;
srom_1(28278) <= 16773518;
srom_1(28279) <= 16736820;
srom_1(28280) <= 16660974;
srom_1(28281) <= 16546337;
srom_1(28282) <= 16393445;
srom_1(28283) <= 16203015;
srom_1(28284) <= 15975941;
srom_1(28285) <= 15713287;
srom_1(28286) <= 15416286;
srom_1(28287) <= 15086329;
srom_1(28288) <= 14724964;
srom_1(28289) <= 14333886;
srom_1(28290) <= 13914928;
srom_1(28291) <= 13470056;
srom_1(28292) <= 13001355;
srom_1(28293) <= 12511023;
srom_1(28294) <= 12001360;
srom_1(28295) <= 11474755;
srom_1(28296) <= 10933679;
srom_1(28297) <= 10380667;
srom_1(28298) <= 9818314;
srom_1(28299) <= 9249257;
srom_1(28300) <= 8676164;
srom_1(28301) <= 8101722;
srom_1(28302) <= 7528626;
srom_1(28303) <= 6959563;
srom_1(28304) <= 6397200;
srom_1(28305) <= 5844176;
srom_1(28306) <= 5303084;
srom_1(28307) <= 4776461;
srom_1(28308) <= 4266777;
srom_1(28309) <= 3776421;
srom_1(28310) <= 3307693;
srom_1(28311) <= 2862792;
srom_1(28312) <= 2443802;
srom_1(28313) <= 2052691;
srom_1(28314) <= 1691290;
srom_1(28315) <= 1361295;
srom_1(28316) <= 1064254;
srom_1(28317) <= 801560;
srom_1(28318) <= 574443;
srom_1(28319) <= 383970;
srom_1(28320) <= 231033;
srom_1(28321) <= 116350;
srom_1(28322) <= 40459;
srom_1(28323) <= 3715;
srom_1(28324) <= 6290;
srom_1(28325) <= 48173;
srom_1(28326) <= 129167;
srom_1(28327) <= 248893;
srom_1(28328) <= 406788;
srom_1(28329) <= 602113;
srom_1(28330) <= 833952;
srom_1(28331) <= 1101216;
srom_1(28332) <= 1402654;
srom_1(28333) <= 1736852;
srom_1(28334) <= 2102242;
srom_1(28335) <= 2497110;
srom_1(28336) <= 2919606;
srom_1(28337) <= 3367748;
srom_1(28338) <= 3839435;
srom_1(28339) <= 4332454;
srom_1(28340) <= 4844494;
srom_1(28341) <= 5373153;
srom_1(28342) <= 5915953;
srom_1(28343) <= 6470348;
srom_1(28344) <= 7033738;
srom_1(28345) <= 7603482;
srom_1(28346) <= 8176908;
srom_1(28347) <= 8751326;
srom_1(28348) <= 9324044;
srom_1(28349) <= 9892374;
srom_1(28350) <= 10453653;
srom_1(28351) <= 11005249;
srom_1(28352) <= 11544574;
srom_1(28353) <= 12069099;
srom_1(28354) <= 12576366;
srom_1(28355) <= 13063995;
srom_1(28356) <= 13529699;
srom_1(28357) <= 13971295;
srom_1(28358) <= 14386711;
srom_1(28359) <= 14774001;
srom_1(28360) <= 15131347;
srom_1(28361) <= 15457074;
srom_1(28362) <= 15749655;
srom_1(28363) <= 16007717;
srom_1(28364) <= 16230051;
srom_1(28365) <= 16415613;
srom_1(28366) <= 16563534;
srom_1(28367) <= 16673120;
srom_1(28368) <= 16743857;
srom_1(28369) <= 16775414;
srom_1(28370) <= 16767641;
srom_1(28371) <= 16720577;
srom_1(28372) <= 16634441;
srom_1(28373) <= 16509638;
srom_1(28374) <= 16346752;
srom_1(28375) <= 16146548;
srom_1(28376) <= 15909964;
srom_1(28377) <= 15638110;
srom_1(28378) <= 15332260;
srom_1(28379) <= 14993849;
srom_1(28380) <= 14624464;
srom_1(28381) <= 14225837;
srom_1(28382) <= 13799838;
srom_1(28383) <= 13348463;
srom_1(28384) <= 12873829;
srom_1(28385) <= 12378163;
srom_1(28386) <= 11863789;
srom_1(28387) <= 11333118;
srom_1(28388) <= 10788639;
srom_1(28389) <= 10232906;
srom_1(28390) <= 9668524;
srom_1(28391) <= 9098140;
srom_1(28392) <= 8524429;
srom_1(28393) <= 7950081;
srom_1(28394) <= 7377789;
srom_1(28395) <= 6810238;
srom_1(28396) <= 6250088;
srom_1(28397) <= 5699966;
srom_1(28398) <= 5162452;
srom_1(28399) <= 4640067;
srom_1(28400) <= 4135260;
srom_1(28401) <= 3650398;
srom_1(28402) <= 3187756;
srom_1(28403) <= 2749502;
srom_1(28404) <= 2337692;
srom_1(28405) <= 1954256;
srom_1(28406) <= 1600994;
srom_1(28407) <= 1279560;
srom_1(28408) <= 991464;
srom_1(28409) <= 738055;
srom_1(28410) <= 520523;
srom_1(28411) <= 339886;
srom_1(28412) <= 196993;
srom_1(28413) <= 92513;
srom_1(28414) <= 26937;
srom_1(28415) <= 571;
srom_1(28416) <= 13539;
srom_1(28417) <= 65781;
srom_1(28418) <= 157052;
srom_1(28419) <= 286923;
srom_1(28420) <= 454786;
srom_1(28421) <= 659853;
srom_1(28422) <= 901163;
srom_1(28423) <= 1177584;
srom_1(28424) <= 1487820;
srom_1(28425) <= 1830416;
srom_1(28426) <= 2203766;
srom_1(28427) <= 2606119;
srom_1(28428) <= 3035588;
srom_1(28429) <= 3490158;
srom_1(28430) <= 3967700;
srom_1(28431) <= 4465973;
srom_1(28432) <= 4982640;
srom_1(28433) <= 5515279;
srom_1(28434) <= 6061392;
srom_1(28435) <= 6618418;
srom_1(28436) <= 7183745;
srom_1(28437) <= 7754722;
srom_1(28438) <= 8328671;
srom_1(28439) <= 8902902;
srom_1(28440) <= 9474721;
srom_1(28441) <= 10041447;
srom_1(28442) <= 10600422;
srom_1(28443) <= 11149025;
srom_1(28444) <= 11684683;
srom_1(28445) <= 12204885;
srom_1(28446) <= 12707192;
srom_1(28447) <= 13189247;
srom_1(28448) <= 13648790;
srom_1(28449) <= 14083666;
srom_1(28450) <= 14491836;
srom_1(28451) <= 14871386;
srom_1(28452) <= 15220536;
srom_1(28453) <= 15537649;
srom_1(28454) <= 15821237;
srom_1(28455) <= 16069972;
srom_1(28456) <= 16282685;
srom_1(28457) <= 16458381;
srom_1(28458) <= 16596235;
srom_1(28459) <= 16695600;
srom_1(28460) <= 16756011;
srom_1(28461) <= 16777185;
srom_1(28462) <= 16759021;
srom_1(28463) <= 16701606;
srom_1(28464) <= 16605208;
srom_1(28465) <= 16470280;
srom_1(28466) <= 16297454;
srom_1(28467) <= 16087540;
srom_1(28468) <= 15841524;
srom_1(28469) <= 15560559;
srom_1(28470) <= 15245961;
srom_1(28471) <= 14899208;
srom_1(28472) <= 14521923;
srom_1(28473) <= 14115878;
srom_1(28474) <= 13682975;
srom_1(28475) <= 13225245;
srom_1(28476) <= 12744835;
srom_1(28477) <= 12243997;
srom_1(28478) <= 11725079;
srom_1(28479) <= 11190516;
srom_1(28480) <= 10642814;
srom_1(28481) <= 10084540;
srom_1(28482) <= 9518314;
srom_1(28483) <= 8946791;
srom_1(28484) <= 8372649;
srom_1(28485) <= 7798583;
srom_1(28486) <= 7227284;
srom_1(28487) <= 6661430;
srom_1(28488) <= 6103676;
srom_1(28489) <= 5556636;
srom_1(28490) <= 5022877;
srom_1(28491) <= 4504900;
srom_1(28492) <= 4005136;
srom_1(28493) <= 3525927;
srom_1(28494) <= 3069521;
srom_1(28495) <= 2638058;
srom_1(28496) <= 2233562;
srom_1(28497) <= 1857928;
srom_1(28498) <= 1512919;
srom_1(28499) <= 1200153;
srom_1(28500) <= 921096;
srom_1(28501) <= 677056;
srom_1(28502) <= 469178;
srom_1(28503) <= 298438;
srom_1(28504) <= 165635;
srom_1(28505) <= 71392;
srom_1(28506) <= 16152;
srom_1(28507) <= 173;
srom_1(28508) <= 23530;
srom_1(28509) <= 86114;
srom_1(28510) <= 187631;
srom_1(28511) <= 327605;
srom_1(28512) <= 505380;
srom_1(28513) <= 720123;
srom_1(28514) <= 970825;
srom_1(28515) <= 1256312;
srom_1(28516) <= 1575245;
srom_1(28517) <= 1926128;
srom_1(28518) <= 2307315;
srom_1(28519) <= 2717020;
srom_1(28520) <= 3153321;
srom_1(28521) <= 3614172;
srom_1(28522) <= 4097412;
srom_1(28523) <= 4600775;
srom_1(28524) <= 5121901;
srom_1(28525) <= 5658345;
srom_1(28526) <= 6207592;
srom_1(28527) <= 6767067;
srom_1(28528) <= 7334145;
srom_1(28529) <= 7906169;
srom_1(28530) <= 8480454;
srom_1(28531) <= 9054309;
srom_1(28532) <= 9625043;
srom_1(28533) <= 10189978;
srom_1(28534) <= 10746466;
srom_1(28535) <= 11291897;
srom_1(28536) <= 11823714;
srom_1(28537) <= 12339422;
srom_1(28538) <= 12836603;
srom_1(28539) <= 13312927;
srom_1(28540) <= 13766158;
srom_1(28541) <= 14194173;
srom_1(28542) <= 14594963;
srom_1(28543) <= 14966649;
srom_1(28544) <= 15307488;
srom_1(28545) <= 15615883;
srom_1(28546) <= 15890386;
srom_1(28547) <= 16129711;
srom_1(28548) <= 16332736;
srom_1(28549) <= 16498507;
srom_1(28550) <= 16626248;
srom_1(28551) <= 16715361;
srom_1(28552) <= 16765426;
srom_1(28553) <= 16776209;
srom_1(28554) <= 16747660;
srom_1(28555) <= 16679913;
srom_1(28556) <= 16573285;
srom_1(28557) <= 16428276;
srom_1(28558) <= 16245566;
srom_1(28559) <= 16026013;
srom_1(28560) <= 15770645;
srom_1(28561) <= 15480660;
srom_1(28562) <= 15157417;
srom_1(28563) <= 14802434;
srom_1(28564) <= 14417374;
srom_1(28565) <= 14004043;
srom_1(28566) <= 13564379;
srom_1(28567) <= 13100445;
srom_1(28568) <= 12614415;
srom_1(28569) <= 12108568;
srom_1(28570) <= 11585278;
srom_1(28571) <= 11046997;
srom_1(28572) <= 10496250;
srom_1(28573) <= 9935620;
srom_1(28574) <= 9367735;
srom_1(28575) <= 8795258;
srom_1(28576) <= 8220875;
srom_1(28577) <= 7647278;
srom_1(28578) <= 7077158;
srom_1(28579) <= 6513188;
srom_1(28580) <= 5958012;
srom_1(28581) <= 5414233;
srom_1(28582) <= 4884403;
srom_1(28583) <= 4371005;
srom_1(28584) <= 3876447;
srom_1(28585) <= 3403048;
srom_1(28586) <= 2953028;
srom_1(28587) <= 2528498;
srom_1(28588) <= 2131447;
srom_1(28589) <= 1763739;
srom_1(28590) <= 1427096;
srom_1(28591) <= 1123099;
srom_1(28592) <= 853172;
srom_1(28593) <= 618581;
srom_1(28594) <= 420427;
srom_1(28595) <= 259638;
srom_1(28596) <= 136969;
srom_1(28597) <= 52994;
srom_1(28598) <= 8108;
srom_1(28599) <= 2521;
srom_1(28600) <= 36259;
srom_1(28601) <= 109165;
srom_1(28602) <= 220895;
srom_1(28603) <= 370927;
srom_1(28604) <= 558556;
srom_1(28605) <= 782903;
srom_1(28606) <= 1042916;
srom_1(28607) <= 1337375;
srom_1(28608) <= 1664900;
srom_1(28609) <= 2023955;
srom_1(28610) <= 2412856;
srom_1(28611) <= 2829779;
srom_1(28612) <= 3272769;
srom_1(28613) <= 3739750;
srom_1(28614) <= 4228530;
srom_1(28615) <= 4736818;
srom_1(28616) <= 5262231;
srom_1(28617) <= 5802305;
srom_1(28618) <= 6354506;
srom_1(28619) <= 6916247;
srom_1(28620) <= 7484891;
srom_1(28621) <= 8057774;
srom_1(28622) <= 8632207;
srom_1(28623) <= 9205499;
srom_1(28624) <= 9774960;
srom_1(28625) <= 10337919;
srom_1(28626) <= 10891738;
srom_1(28627) <= 11433819;
srom_1(28628) <= 11961619;
srom_1(28629) <= 12472665;
srom_1(28630) <= 12964559;
srom_1(28631) <= 13434995;
srom_1(28632) <= 13881766;
srom_1(28633) <= 14302778;
srom_1(28634) <= 14696057;
srom_1(28635) <= 15059758;
srom_1(28636) <= 15392175;
srom_1(28637) <= 15691751;
srom_1(28638) <= 15957079;
srom_1(28639) <= 16186916;
srom_1(28640) <= 16380185;
srom_1(28641) <= 16535978;
srom_1(28642) <= 16653565;
srom_1(28643) <= 16732395;
srom_1(28644) <= 16772098;
srom_1(28645) <= 16772488;
srom_1(28646) <= 16733563;
srom_1(28647) <= 16655506;
srom_1(28648) <= 16538682;
srom_1(28649) <= 16383640;
srom_1(28650) <= 16191107;
srom_1(28651) <= 15961984;
srom_1(28652) <= 15697348;
srom_1(28653) <= 15398439;
srom_1(28654) <= 15066658;
srom_1(28655) <= 14703561;
srom_1(28656) <= 14310851;
srom_1(28657) <= 13890370;
srom_1(28658) <= 13444089;
srom_1(28659) <= 12974102;
srom_1(28660) <= 12482611;
srom_1(28661) <= 11971922;
srom_1(28662) <= 11444430;
srom_1(28663) <= 10902608;
srom_1(28664) <= 10348997;
srom_1(28665) <= 9786193;
srom_1(28666) <= 9216835;
srom_1(28667) <= 8643593;
srom_1(28668) <= 8069156;
srom_1(28669) <= 7496217;
srom_1(28670) <= 6927462;
srom_1(28671) <= 6365559;
srom_1(28672) <= 5813143;
srom_1(28673) <= 5272804;
srom_1(28674) <= 4747077;
srom_1(28675) <= 4238425;
srom_1(28676) <= 3749235;
srom_1(28677) <= 3281801;
srom_1(28678) <= 2838315;
srom_1(28679) <= 2420855;
srom_1(28680) <= 2031381;
srom_1(28681) <= 1671718;
srom_1(28682) <= 1343552;
srom_1(28683) <= 1048423;
srom_1(28684) <= 787715;
srom_1(28685) <= 562650;
srom_1(28686) <= 374284;
srom_1(28687) <= 223499;
srom_1(28688) <= 111004;
srom_1(28689) <= 37325;
srom_1(28690) <= 2808;
srom_1(28691) <= 7615;
srom_1(28692) <= 51723;
srom_1(28693) <= 134926;
srom_1(28694) <= 256833;
srom_1(28695) <= 416873;
srom_1(28696) <= 614295;
srom_1(28697) <= 848174;
srom_1(28698) <= 1117412;
srom_1(28699) <= 1420747;
srom_1(28700) <= 1756757;
srom_1(28701) <= 2123866;
srom_1(28702) <= 2520353;
srom_1(28703) <= 2944357;
srom_1(28704) <= 3393892;
srom_1(28705) <= 3866849;
srom_1(28706) <= 4361009;
srom_1(28707) <= 4874057;
srom_1(28708) <= 5403585;
srom_1(28709) <= 5947112;
srom_1(28710) <= 6502087;
srom_1(28711) <= 7065909;
srom_1(28712) <= 7635933;
srom_1(28713) <= 8209487;
srom_1(28714) <= 8783881;
srom_1(28715) <= 9356421;
srom_1(28716) <= 9924423;
srom_1(28717) <= 10485223;
srom_1(28718) <= 11036191;
srom_1(28719) <= 11574744;
srom_1(28720) <= 12098355;
srom_1(28721) <= 12604571;
srom_1(28722) <= 13091016;
srom_1(28723) <= 13555411;
srom_1(28724) <= 13995576;
srom_1(28725) <= 14409448;
srom_1(28726) <= 14795087;
srom_1(28727) <= 15150683;
srom_1(28728) <= 15474570;
srom_1(28729) <= 15765228;
srom_1(28730) <= 16021294;
srom_1(28731) <= 16241568;
srom_1(28732) <= 16425017;
srom_1(28733) <= 16570781;
srom_1(28734) <= 16678176;
srom_1(28735) <= 16746697;
srom_1(28736) <= 16776025;
srom_1(28737) <= 16766022;
srom_1(28738) <= 16716734;
srom_1(28739) <= 16628392;
srom_1(28740) <= 16501411;
srom_1(28741) <= 16336387;
srom_1(28742) <= 16134092;
srom_1(28743) <= 15895477;
srom_1(28744) <= 15621659;
srom_1(28745) <= 15313923;
srom_1(28746) <= 14973711;
srom_1(28747) <= 14602620;
srom_1(28748) <= 14202389;
srom_1(28749) <= 13774896;
srom_1(28750) <= 13322144;
srom_1(28751) <= 12846257;
srom_1(28752) <= 12349467;
srom_1(28753) <= 11834102;
srom_1(28754) <= 11302581;
srom_1(28755) <= 10757395;
srom_1(28756) <= 10201101;
srom_1(28757) <= 9636308;
srom_1(28758) <= 9065664;
srom_1(28759) <= 8491844;
srom_1(28760) <= 7917541;
srom_1(28761) <= 7345447;
srom_1(28762) <= 6778244;
srom_1(28763) <= 6218593;
srom_1(28764) <= 5669118;
srom_1(28765) <= 5132395;
srom_1(28766) <= 4610942;
srom_1(28767) <= 4107204;
srom_1(28768) <= 3623543;
srom_1(28769) <= 3162226;
srom_1(28770) <= 2725418;
srom_1(28771) <= 2315167;
srom_1(28772) <= 1933396;
srom_1(28773) <= 1581896;
srom_1(28774) <= 1262315;
srom_1(28775) <= 976151;
srom_1(28776) <= 724747;
srom_1(28777) <= 509282;
srom_1(28778) <= 330765;
srom_1(28779) <= 190034;
srom_1(28780) <= 87749;
srom_1(28781) <= 24390;
srom_1(28782) <= 254;
srom_1(28783) <= 15453;
srom_1(28784) <= 69917;
srom_1(28785) <= 163390;
srom_1(28786) <= 295434;
srom_1(28787) <= 465430;
srom_1(28788) <= 672580;
srom_1(28789) <= 915913;
srom_1(28790) <= 1194288;
srom_1(28791) <= 1506400;
srom_1(28792) <= 1850785;
srom_1(28793) <= 2225828;
srom_1(28794) <= 2629771;
srom_1(28795) <= 3060718;
srom_1(28796) <= 3516650;
srom_1(28797) <= 3995428;
srom_1(28798) <= 4494807;
srom_1(28799) <= 5012446;
srom_1(28800) <= 5545917;
srom_1(28801) <= 6092718;
srom_1(28802) <= 6650285;
srom_1(28803) <= 7216004;
srom_1(28804) <= 7787221;
srom_1(28805) <= 8361259;
srom_1(28806) <= 8935425;
srom_1(28807) <= 9507026;
srom_1(28808) <= 10073383;
srom_1(28809) <= 10631840;
srom_1(28810) <= 11179777;
srom_1(28811) <= 11714625;
srom_1(28812) <= 12233877;
srom_1(28813) <= 12735097;
srom_1(28814) <= 13215934;
srom_1(28815) <= 13674135;
srom_1(28816) <= 14107550;
srom_1(28817) <= 14514147;
srom_1(28818) <= 14892019;
srom_1(28819) <= 15239394;
srom_1(28820) <= 15554644;
srom_1(28821) <= 15836289;
srom_1(28822) <= 16083010;
srom_1(28823) <= 16293649;
srom_1(28824) <= 16467219;
srom_1(28825) <= 16602906;
srom_1(28826) <= 16700072;
srom_1(28827) <= 16758264;
srom_1(28828) <= 16777207;
srom_1(28829) <= 16756813;
srom_1(28830) <= 16697178;
srom_1(28831) <= 16598581;
srom_1(28832) <= 16461484;
srom_1(28833) <= 16286531;
srom_1(28834) <= 16074542;
srom_1(28835) <= 15826511;
srom_1(28836) <= 15543602;
srom_1(28837) <= 15227140;
srom_1(28838) <= 14878609;
srom_1(28839) <= 14499645;
srom_1(28840) <= 14092024;
srom_1(28841) <= 13657658;
srom_1(28842) <= 13198583;
srom_1(28843) <= 12716953;
srom_1(28844) <= 12215026;
srom_1(28845) <= 11695155;
srom_1(28846) <= 11159779;
srom_1(28847) <= 10611407;
srom_1(28848) <= 10052613;
srom_1(28849) <= 9486015;
srom_1(28850) <= 8914271;
srom_1(28851) <= 8340062;
srom_1(28852) <= 7766081;
srom_1(28853) <= 7195018;
srom_1(28854) <= 6629554;
srom_1(28855) <= 6072337;
srom_1(28856) <= 5525983;
srom_1(28857) <= 4993052;
srom_1(28858) <= 4476045;
srom_1(28859) <= 3977385;
srom_1(28860) <= 3499410;
srom_1(28861) <= 3044363;
srom_1(28862) <= 2614376;
srom_1(28863) <= 2211467;
srom_1(28864) <= 1837525;
srom_1(28865) <= 1494303;
srom_1(28866) <= 1183410;
srom_1(28867) <= 906306;
srom_1(28868) <= 664288;
srom_1(28869) <= 458492;
srom_1(28870) <= 289884;
srom_1(28871) <= 159253;
srom_1(28872) <= 67212;
srom_1(28873) <= 14194;
srom_1(28874) <= 445;
srom_1(28875) <= 26032;
srom_1(28876) <= 90834;
srom_1(28877) <= 194547;
srom_1(28878) <= 336684;
srom_1(28879) <= 516580;
srom_1(28880) <= 733390;
srom_1(28881) <= 986099;
srom_1(28882) <= 1273520;
srom_1(28883) <= 1594306;
srom_1(28884) <= 1946954;
srom_1(28885) <= 2329808;
srom_1(28886) <= 2741074;
srom_1(28887) <= 3178823;
srom_1(28888) <= 3641003;
srom_1(28889) <= 4125446;
srom_1(28890) <= 4629880;
srom_1(28891) <= 5151941;
srom_1(28892) <= 5689179;
srom_1(28893) <= 6239075;
srom_1(28894) <= 6799052;
srom_1(28895) <= 7366483;
srom_1(28896) <= 7938706;
srom_1(28897) <= 8513040;
srom_1(28898) <= 9086789;
srom_1(28899) <= 9657265;
srom_1(28900) <= 10221792;
srom_1(28901) <= 10777722;
srom_1(28902) <= 11322449;
srom_1(28903) <= 11853418;
srom_1(28904) <= 12368139;
srom_1(28905) <= 12864199;
srom_1(28906) <= 13339272;
srom_1(28907) <= 13791129;
srom_1(28908) <= 14217651;
srom_1(28909) <= 14616840;
srom_1(28910) <= 14986822;
srom_1(28911) <= 15325862;
srom_1(28912) <= 15632372;
srom_1(28913) <= 15904913;
srom_1(28914) <= 16142207;
srom_1(28915) <= 16343142;
srom_1(28916) <= 16506776;
srom_1(28917) <= 16632341;
srom_1(28918) <= 16719248;
srom_1(28919) <= 16767090;
srom_1(28920) <= 16775642;
srom_1(28921) <= 16744864;
srom_1(28922) <= 16674902;
srom_1(28923) <= 16566081;
srom_1(28924) <= 16418914;
srom_1(28925) <= 16234090;
srom_1(28926) <= 16012476;
srom_1(28927) <= 15755111;
srom_1(28928) <= 15463202;
srom_1(28929) <= 15138117;
srom_1(28930) <= 14781382;
srom_1(28931) <= 14394669;
srom_1(28932) <= 13979792;
srom_1(28933) <= 13538695;
srom_1(28934) <= 13073448;
srom_1(28935) <= 12586232;
srom_1(28936) <= 12079332;
srom_1(28937) <= 11555125;
srom_1(28938) <= 11016069;
srom_1(28939) <= 10464692;
srom_1(28940) <= 9903579;
srom_1(28941) <= 9335362;
srom_1(28942) <= 8762706;
srom_1(28943) <= 8188295;
srom_1(28944) <= 7614824;
srom_1(28945) <= 7044981;
srom_1(28946) <= 6481439;
srom_1(28947) <= 5926840;
srom_1(28948) <= 5383785;
srom_1(28949) <= 4854821;
srom_1(28950) <= 4342428;
srom_1(28951) <= 3849009;
srom_1(28952) <= 3376878;
srom_1(28953) <= 2928248;
srom_1(28954) <= 2505224;
srom_1(28955) <= 2109789;
srom_1(28956) <= 1743798;
srom_1(28957) <= 1408967;
srom_1(28958) <= 1106865;
srom_1(28959) <= 838910;
srom_1(28960) <= 606358;
srom_1(28961) <= 410300;
srom_1(28962) <= 251654;
srom_1(28963) <= 131166;
srom_1(28964) <= 49400;
srom_1(28965) <= 6739;
srom_1(28966) <= 3383;
srom_1(28967) <= 39349;
srom_1(28968) <= 114467;
srom_1(28969) <= 228386;
srom_1(28970) <= 380571;
srom_1(28971) <= 570308;
srom_1(28972) <= 796707;
srom_1(28973) <= 1058708;
srom_1(28974) <= 1355081;
srom_1(28975) <= 1684437;
srom_1(28976) <= 2045231;
srom_1(28977) <= 2435771;
srom_1(28978) <= 2854226;
srom_1(28979) <= 3298634;
srom_1(28980) <= 3766910;
srom_1(28981) <= 4256860;
srom_1(28982) <= 4766184;
srom_1(28983) <= 5292495;
srom_1(28984) <= 5833325;
srom_1(28985) <= 6386137;
srom_1(28986) <= 6948340;
srom_1(28987) <= 7517296;
srom_1(28988) <= 8090339;
srom_1(28989) <= 8664780;
srom_1(28990) <= 9237926;
srom_1(28991) <= 9807089;
srom_1(28992) <= 10369600;
srom_1(28993) <= 10922822;
srom_1(28994) <= 11464161;
srom_1(28995) <= 11991076;
srom_1(28996) <= 12501099;
srom_1(28997) <= 12991837;
srom_1(28998) <= 13460988;
srom_1(28999) <= 13906354;
srom_1(29000) <= 14325845;
srom_1(29001) <= 14717494;
srom_1(29002) <= 15079464;
srom_1(29003) <= 15410059;
srom_1(29004) <= 15707728;
srom_1(29005) <= 15971076;
srom_1(29006) <= 16198866;
srom_1(29007) <= 16390031;
srom_1(29008) <= 16543675;
srom_1(29009) <= 16659077;
srom_1(29010) <= 16735696;
srom_1(29011) <= 16773173;
srom_1(29012) <= 16771331;
srom_1(29013) <= 16730180;
srom_1(29014) <= 16649912;
srom_1(29015) <= 16530905;
srom_1(29016) <= 16373715;
srom_1(29017) <= 16179081;
srom_1(29018) <= 15947914;
srom_1(29019) <= 15681299;
srom_1(29020) <= 15380486;
srom_1(29021) <= 15046886;
srom_1(29022) <= 14682062;
srom_1(29023) <= 14287727;
srom_1(29024) <= 13865729;
srom_1(29025) <= 13418046;
srom_1(29026) <= 12946779;
srom_1(29027) <= 12454137;
srom_1(29028) <= 11942430;
srom_1(29029) <= 11414058;
srom_1(29030) <= 10871499;
srom_1(29031) <= 10317296;
srom_1(29032) <= 9754050;
srom_1(29033) <= 9184400;
srom_1(29034) <= 8611019;
srom_1(29035) <= 8036594;
srom_1(29036) <= 7463820;
srom_1(29037) <= 6895383;
srom_1(29038) <= 6333949;
srom_1(29039) <= 5782149;
srom_1(29040) <= 5242571;
srom_1(29041) <= 4717747;
srom_1(29042) <= 4210136;
srom_1(29043) <= 3722120;
srom_1(29044) <= 3255987;
srom_1(29045) <= 2813922;
srom_1(29046) <= 2397999;
srom_1(29047) <= 2010167;
srom_1(29048) <= 1652247;
srom_1(29049) <= 1325915;
srom_1(29050) <= 1032703;
srom_1(29051) <= 773986;
srom_1(29052) <= 550976;
srom_1(29053) <= 364719;
srom_1(29054) <= 216089;
srom_1(29055) <= 105783;
srom_1(29056) <= 34317;
srom_1(29057) <= 2028;
srom_1(29058) <= 9067;
srom_1(29059) <= 55400;
srom_1(29060) <= 140810;
srom_1(29061) <= 264897;
srom_1(29062) <= 427079;
srom_1(29063) <= 626595;
srom_1(29064) <= 862510;
srom_1(29065) <= 1133717;
srom_1(29066) <= 1438945;
srom_1(29067) <= 1776763;
srom_1(29068) <= 2145585;
srom_1(29069) <= 2543684;
srom_1(29070) <= 2969191;
srom_1(29071) <= 3420111;
srom_1(29072) <= 3894331;
srom_1(29073) <= 4389626;
srom_1(29074) <= 4903673;
srom_1(29075) <= 5434063;
srom_1(29076) <= 5978307;
srom_1(29077) <= 6533854;
srom_1(29078) <= 7098099;
srom_1(29079) <= 7668395;
srom_1(29080) <= 8242069;
srom_1(29081) <= 8816429;
srom_1(29082) <= 9388784;
srom_1(29083) <= 9956448;
srom_1(29084) <= 10516760;
srom_1(29085) <= 11067093;
srom_1(29086) <= 11604865;
srom_1(29087) <= 12127555;
srom_1(29088) <= 12632712;
srom_1(29089) <= 13117967;
srom_1(29090) <= 13581044;
srom_1(29091) <= 14019772;
srom_1(29092) <= 14432094;
srom_1(29093) <= 14816076;
srom_1(29094) <= 15169917;
srom_1(29095) <= 15491958;
srom_1(29096) <= 15780689;
srom_1(29097) <= 16034756;
srom_1(29098) <= 16252967;
srom_1(29099) <= 16434300;
srom_1(29100) <= 16577904;
srom_1(29101) <= 16683106;
srom_1(29102) <= 16749412;
srom_1(29103) <= 16776511;
srom_1(29104) <= 16764276;
srom_1(29105) <= 16712765;
srom_1(29106) <= 16622219;
srom_1(29107) <= 16493063;
srom_1(29108) <= 16325902;
srom_1(29109) <= 16121520;
srom_1(29110) <= 15880877;
srom_1(29111) <= 15605099;
srom_1(29112) <= 15295481;
srom_1(29113) <= 14953474;
srom_1(29114) <= 14580682;
srom_1(29115) <= 14178854;
srom_1(29116) <= 13749872;
srom_1(29117) <= 13295751;
srom_1(29118) <= 12818617;
srom_1(29119) <= 12320710;
srom_1(29120) <= 11804364;
srom_1(29121) <= 11272001;
srom_1(29122) <= 10726116;
srom_1(29123) <= 10169270;
srom_1(29124) <= 9604073;
srom_1(29125) <= 9033177;
srom_1(29126) <= 8459258;
srom_1(29127) <= 7885008;
srom_1(29128) <= 7313120;
srom_1(29129) <= 6746275;
srom_1(29130) <= 6187131;
srom_1(29131) <= 5638311;
srom_1(29132) <= 5102387;
srom_1(29133) <= 4581874;
srom_1(29134) <= 4079213;
srom_1(29135) <= 3596759;
srom_1(29136) <= 3136776;
srom_1(29137) <= 2701420;
srom_1(29138) <= 2292734;
srom_1(29139) <= 1912634;
srom_1(29140) <= 1562901;
srom_1(29141) <= 1245177;
srom_1(29142) <= 960950;
srom_1(29143) <= 711555;
srom_1(29144) <= 498159;
srom_1(29145) <= 321765;
srom_1(29146) <= 183199;
srom_1(29147) <= 83111;
srom_1(29148) <= 21970;
srom_1(29149) <= 63;
srom_1(29150) <= 17493;
srom_1(29151) <= 74178;
srom_1(29152) <= 169853;
srom_1(29153) <= 304067;
srom_1(29154) <= 476193;
srom_1(29155) <= 685423;
srom_1(29156) <= 930776;
srom_1(29157) <= 1211101;
srom_1(29158) <= 1525084;
srom_1(29159) <= 1871253;
srom_1(29160) <= 2247983;
srom_1(29161) <= 2653509;
srom_1(29162) <= 3085929;
srom_1(29163) <= 3543215;
srom_1(29164) <= 4023223;
srom_1(29165) <= 4523701;
srom_1(29166) <= 5042304;
srom_1(29167) <= 5576598;
srom_1(29168) <= 6124078;
srom_1(29169) <= 6682178;
srom_1(29170) <= 7248280;
srom_1(29171) <= 7819730;
srom_1(29172) <= 8393846;
srom_1(29173) <= 8967939;
srom_1(29174) <= 9539315;
srom_1(29175) <= 10105294;
srom_1(29176) <= 10663224;
srom_1(29177) <= 11210487;
srom_1(29178) <= 11744517;
srom_1(29179) <= 12262810;
srom_1(29180) <= 12762936;
srom_1(29181) <= 13242549;
srom_1(29182) <= 13699400;
srom_1(29183) <= 14131347;
srom_1(29184) <= 14536365;
srom_1(29185) <= 14912553;
srom_1(29186) <= 15258149;
srom_1(29187) <= 15571530;
srom_1(29188) <= 15851229;
srom_1(29189) <= 16095933;
srom_1(29190) <= 16304494;
srom_1(29191) <= 16475935;
srom_1(29192) <= 16609452;
srom_1(29193) <= 16704419;
srom_1(29194) <= 16760390;
srom_1(29195) <= 16777102;
srom_1(29196) <= 16754478;
srom_1(29197) <= 16692624;
srom_1(29198) <= 16591829;
srom_1(29199) <= 16452567;
srom_1(29200) <= 16275490;
srom_1(29201) <= 16061428;
srom_1(29202) <= 15811387;
srom_1(29203) <= 15526537;
srom_1(29204) <= 15208215;
srom_1(29205) <= 14857913;
srom_1(29206) <= 14477275;
srom_1(29207) <= 14068084;
srom_1(29208) <= 13632261;
srom_1(29209) <= 13171848;
srom_1(29210) <= 12689006;
srom_1(29211) <= 12185997;
srom_1(29212) <= 11665181;
srom_1(29213) <= 11129000;
srom_1(29214) <= 10579968;
srom_1(29215) <= 10020660;
srom_1(29216) <= 9453699;
srom_1(29217) <= 8881743;
srom_1(29218) <= 8307475;
srom_1(29219) <= 7733587;
srom_1(29220) <= 7162771;
srom_1(29221) <= 6597704;
srom_1(29222) <= 6041034;
srom_1(29223) <= 5495373;
srom_1(29224) <= 4963279;
srom_1(29225) <= 4447248;
srom_1(29226) <= 3949700;
srom_1(29227) <= 3472966;
srom_1(29228) <= 3019284;
srom_1(29229) <= 2590781;
srom_1(29230) <= 2189466;
srom_1(29231) <= 1817220;
srom_1(29232) <= 1475790;
srom_1(29233) <= 1166777;
srom_1(29234) <= 891629;
srom_1(29235) <= 651637;
srom_1(29236) <= 447926;
srom_1(29237) <= 281452;
srom_1(29238) <= 152995;
srom_1(29239) <= 63158;
srom_1(29240) <= 12362;
srom_1(29241) <= 845;
srom_1(29242) <= 28661;
srom_1(29243) <= 95679;
srom_1(29244) <= 201586;
srom_1(29245) <= 345885;
srom_1(29246) <= 527898;
srom_1(29247) <= 746774;
srom_1(29248) <= 1001484;
srom_1(29249) <= 1290836;
srom_1(29250) <= 1613471;
srom_1(29251) <= 1967877;
srom_1(29252) <= 2352392;
srom_1(29253) <= 2765213;
srom_1(29254) <= 3204404;
srom_1(29255) <= 3667905;
srom_1(29256) <= 4153544;
srom_1(29257) <= 4659042;
srom_1(29258) <= 5182029;
srom_1(29259) <= 5720053;
srom_1(29260) <= 6270591;
srom_1(29261) <= 6831061;
srom_1(29262) <= 7398835;
srom_1(29263) <= 7971250;
srom_1(29264) <= 8545623;
srom_1(29265) <= 9119259;
srom_1(29266) <= 9689469;
srom_1(29267) <= 10253578;
srom_1(29268) <= 10808942;
srom_1(29269) <= 11352956;
srom_1(29270) <= 11883070;
srom_1(29271) <= 12396797;
srom_1(29272) <= 12891728;
srom_1(29273) <= 13365542;
srom_1(29274) <= 13816017;
srom_1(29275) <= 14241042;
srom_1(29276) <= 14638623;
srom_1(29277) <= 15006895;
srom_1(29278) <= 15344132;
srom_1(29279) <= 15648751;
srom_1(29280) <= 15919326;
srom_1(29281) <= 16154586;
srom_1(29282) <= 16353429;
srom_1(29283) <= 16514923;
srom_1(29284) <= 16638309;
srom_1(29285) <= 16723009;
srom_1(29286) <= 16768627;
srom_1(29287) <= 16774948;
srom_1(29288) <= 16741942;
srom_1(29289) <= 16669765;
srom_1(29290) <= 16558754;
srom_1(29291) <= 16409431;
srom_1(29292) <= 16222496;
srom_1(29293) <= 15998824;
srom_1(29294) <= 15739466;
srom_1(29295) <= 15445637;
srom_1(29296) <= 15118716;
srom_1(29297) <= 14760234;
srom_1(29298) <= 14371874;
srom_1(29299) <= 13955456;
srom_1(29300) <= 13512933;
srom_1(29301) <= 13046380;
srom_1(29302) <= 12557986;
srom_1(29303) <= 12050040;
srom_1(29304) <= 11524924;
srom_1(29305) <= 10985101;
srom_1(29306) <= 10433102;
srom_1(29307) <= 9871516;
srom_1(29308) <= 9302976;
srom_1(29309) <= 8730148;
srom_1(29310) <= 8155718;
srom_1(29311) <= 7582381;
srom_1(29312) <= 7012824;
srom_1(29313) <= 6449719;
srom_1(29314) <= 5895706;
srom_1(29315) <= 5353383;
srom_1(29316) <= 4825293;
srom_1(29317) <= 4313913;
srom_1(29318) <= 3821640;
srom_1(29319) <= 3350783;
srom_1(29320) <= 2903551;
srom_1(29321) <= 2482040;
srom_1(29322) <= 2088226;
srom_1(29323) <= 1723958;
srom_1(29324) <= 1390942;
srom_1(29325) <= 1090741;
srom_1(29326) <= 824762;
srom_1(29327) <= 594252;
srom_1(29328) <= 400293;
srom_1(29329) <= 243794;
srom_1(29330) <= 125488;
srom_1(29331) <= 45931;
srom_1(29332) <= 5496;
srom_1(29333) <= 4372;
srom_1(29334) <= 42565;
srom_1(29335) <= 119895;
srom_1(29336) <= 236000;
srom_1(29337) <= 390335;
srom_1(29338) <= 582177;
srom_1(29339) <= 810626;
srom_1(29340) <= 1074611;
srom_1(29341) <= 1372893;
srom_1(29342) <= 1704075;
srom_1(29343) <= 2066603;
srom_1(29344) <= 2458777;
srom_1(29345) <= 2878757;
srom_1(29346) <= 3324576;
srom_1(29347) <= 3794141;
srom_1(29348) <= 4285251;
srom_1(29349) <= 4795604;
srom_1(29350) <= 5322805;
srom_1(29351) <= 5864383;
srom_1(29352) <= 6417798;
srom_1(29353) <= 6980454;
srom_1(29354) <= 7549714;
srom_1(29355) <= 8122908;
srom_1(29356) <= 8697348;
srom_1(29357) <= 9270340;
srom_1(29358) <= 9839197;
srom_1(29359) <= 10401251;
srom_1(29360) <= 10953868;
srom_1(29361) <= 11494456;
srom_1(29362) <= 12020479;
srom_1(29363) <= 12529471;
srom_1(29364) <= 13019045;
srom_1(29365) <= 13486905;
srom_1(29366) <= 13930858;
srom_1(29367) <= 14348821;
srom_1(29368) <= 14738835;
srom_1(29369) <= 15099070;
srom_1(29370) <= 15427837;
srom_1(29371) <= 15723596;
srom_1(29372) <= 15984957;
srom_1(29373) <= 16210697;
srom_1(29374) <= 16399757;
srom_1(29375) <= 16551249;
srom_1(29376) <= 16664465;
srom_1(29377) <= 16738871;
srom_1(29378) <= 16774121;
srom_1(29379) <= 16770048;
srom_1(29380) <= 16726671;
srom_1(29381) <= 16644194;
srom_1(29382) <= 16523005;
srom_1(29383) <= 16363670;
srom_1(29384) <= 16166937;
srom_1(29385) <= 15933729;
srom_1(29386) <= 15665139;
srom_1(29387) <= 15362428;
srom_1(29388) <= 15027013;
srom_1(29389) <= 14660469;
srom_1(29390) <= 14264514;
srom_1(29391) <= 13841005;
srom_1(29392) <= 13391927;
srom_1(29393) <= 12919387;
srom_1(29394) <= 12425601;
srom_1(29395) <= 11912884;
srom_1(29396) <= 11383641;
srom_1(29397) <= 10840353;
srom_1(29398) <= 10285567;
srom_1(29399) <= 9721886;
srom_1(29400) <= 9151953;
srom_1(29401) <= 8578441;
srom_1(29402) <= 8004038;
srom_1(29403) <= 7431438;
srom_1(29404) <= 6863327;
srom_1(29405) <= 6302369;
srom_1(29406) <= 5751194;
srom_1(29407) <= 5212386;
srom_1(29408) <= 4688473;
srom_1(29409) <= 4181911;
srom_1(29410) <= 3695075;
srom_1(29411) <= 3230250;
srom_1(29412) <= 2789613;
srom_1(29413) <= 2375232;
srom_1(29414) <= 1989050;
srom_1(29415) <= 1632878;
srom_1(29416) <= 1308385;
srom_1(29417) <= 1017094;
srom_1(29418) <= 760371;
srom_1(29419) <= 539419;
srom_1(29420) <= 355275;
srom_1(29421) <= 208802;
srom_1(29422) <= 100686;
srom_1(29423) <= 31436;
srom_1(29424) <= 1375;
srom_1(29425) <= 10645;
srom_1(29426) <= 59202;
srom_1(29427) <= 146818;
srom_1(29428) <= 273083;
srom_1(29429) <= 437404;
srom_1(29430) <= 639012;
srom_1(29431) <= 876959;
srom_1(29432) <= 1150132;
srom_1(29433) <= 1457248;
srom_1(29434) <= 1796868;
srom_1(29435) <= 2167399;
srom_1(29436) <= 2567103;
srom_1(29437) <= 2994106;
srom_1(29438) <= 3446406;
srom_1(29439) <= 3921881;
srom_1(29440) <= 4418302;
srom_1(29441) <= 4933342;
srom_1(29442) <= 5464584;
srom_1(29443) <= 6009539;
srom_1(29444) <= 6565649;
srom_1(29445) <= 7130308;
srom_1(29446) <= 7700868;
srom_1(29447) <= 8274652;
srom_1(29448) <= 8848971;
srom_1(29449) <= 9421132;
srom_1(29450) <= 9988450;
srom_1(29451) <= 10548266;
srom_1(29452) <= 11097955;
srom_1(29453) <= 11634938;
srom_1(29454) <= 12156699;
srom_1(29455) <= 12660789;
srom_1(29456) <= 13144846;
srom_1(29457) <= 13606599;
srom_1(29458) <= 14043884;
srom_1(29459) <= 14454648;
srom_1(29460) <= 14836967;
srom_1(29461) <= 15189048;
srom_1(29462) <= 15509239;
srom_1(29463) <= 15796038;
srom_1(29464) <= 16048102;
srom_1(29465) <= 16264248;
srom_1(29466) <= 16443462;
srom_1(29467) <= 16584904;
srom_1(29468) <= 16687911;
srom_1(29469) <= 16751999;
srom_1(29470) <= 16776869;
srom_1(29471) <= 16762403;
srom_1(29472) <= 16708670;
srom_1(29473) <= 16615921;
srom_1(29474) <= 16484592;
srom_1(29475) <= 16315297;
srom_1(29476) <= 16108832;
srom_1(29477) <= 15866163;
srom_1(29478) <= 15588430;
srom_1(29479) <= 15276935;
srom_1(29480) <= 14933137;
srom_1(29481) <= 14558651;
srom_1(29482) <= 14155230;
srom_1(29483) <= 13724768;
srom_1(29484) <= 13269283;
srom_1(29485) <= 12790911;
srom_1(29486) <= 12291895;
srom_1(29487) <= 11774575;
srom_1(29488) <= 11241377;
srom_1(29489) <= 10694801;
srom_1(29490) <= 10137411;
srom_1(29491) <= 9571820;
srom_1(29492) <= 9000681;
srom_1(29493) <= 8426671;
srom_1(29494) <= 7852483;
srom_1(29495) <= 7280809;
srom_1(29496) <= 6714330;
srom_1(29497) <= 6155702;
srom_1(29498) <= 5607545;
srom_1(29499) <= 5072429;
srom_1(29500) <= 4552864;
srom_1(29501) <= 4051286;
srom_1(29502) <= 3570047;
srom_1(29503) <= 3111405;
srom_1(29504) <= 2677508;
srom_1(29505) <= 2270393;
srom_1(29506) <= 1891969;
srom_1(29507) <= 1544009;
srom_1(29508) <= 1228146;
srom_1(29509) <= 945861;
srom_1(29510) <= 698478;
srom_1(29511) <= 487156;
srom_1(29512) <= 312887;
srom_1(29513) <= 176487;
srom_1(29514) <= 78598;
srom_1(29515) <= 19676;
srom_1(29516) <= 0;
srom_1(29517) <= 19660;
srom_1(29518) <= 78565;
srom_1(29519) <= 176439;
srom_1(29520) <= 312823;
srom_1(29521) <= 487076;
srom_1(29522) <= 698383;
srom_1(29523) <= 945752;
srom_1(29524) <= 1228023;
srom_1(29525) <= 1543872;
srom_1(29526) <= 1891819;
srom_1(29527) <= 2270231;
srom_1(29528) <= 2677335;
srom_1(29529) <= 3111220;
srom_1(29530) <= 3569853;
srom_1(29531) <= 4051083;
srom_1(29532) <= 4552653;
srom_1(29533) <= 5072211;
srom_1(29534) <= 5607321;
srom_1(29535) <= 6155473;
srom_1(29536) <= 6714098;
srom_1(29537) <= 7280574;
srom_1(29538) <= 7852247;
srom_1(29539) <= 8426434;
srom_1(29540) <= 9000444;
srom_1(29541) <= 9571586;
srom_1(29542) <= 10137179;
srom_1(29543) <= 10694573;
srom_1(29544) <= 11241154;
srom_1(29545) <= 11774358;
srom_1(29546) <= 12291685;
srom_1(29547) <= 12790709;
srom_1(29548) <= 13269090;
srom_1(29549) <= 13724585;
srom_1(29550) <= 14155058;
srom_1(29551) <= 14558490;
srom_1(29552) <= 14932989;
srom_1(29553) <= 15276799;
srom_1(29554) <= 15588309;
srom_1(29555) <= 15866056;
srom_1(29556) <= 16108739;
srom_1(29557) <= 16315219;
srom_1(29558) <= 16484529;
srom_1(29559) <= 16615875;
srom_1(29560) <= 16708640;
srom_1(29561) <= 16762389;
srom_1(29562) <= 16776871;
srom_1(29563) <= 16752018;
srom_1(29564) <= 16687945;
srom_1(29565) <= 16584954;
srom_1(29566) <= 16443528;
srom_1(29567) <= 16264329;
srom_1(29568) <= 16048199;
srom_1(29569) <= 15796150;
srom_1(29570) <= 15509364;
srom_1(29571) <= 15189187;
srom_1(29572) <= 14837119;
srom_1(29573) <= 14454812;
srom_1(29574) <= 14044059;
srom_1(29575) <= 13606785;
srom_1(29576) <= 13145042;
srom_1(29577) <= 12660993;
srom_1(29578) <= 12156911;
srom_1(29579) <= 11635157;
srom_1(29580) <= 11098179;
srom_1(29581) <= 10548495;
srom_1(29582) <= 9988683;
srom_1(29583) <= 9421367;
srom_1(29584) <= 8849208;
srom_1(29585) <= 8274889;
srom_1(29586) <= 7701104;
srom_1(29587) <= 7130543;
srom_1(29588) <= 6565881;
srom_1(29589) <= 6009766;
srom_1(29590) <= 5464807;
srom_1(29591) <= 4933558;
srom_1(29592) <= 4418511;
srom_1(29593) <= 3922082;
srom_1(29594) <= 3446597;
srom_1(29595) <= 2994287;
srom_1(29596) <= 2567273;
srom_1(29597) <= 2167558;
srom_1(29598) <= 1797015;
srom_1(29599) <= 1457382;
srom_1(29600) <= 1150252;
srom_1(29601) <= 877065;
srom_1(29602) <= 639102;
srom_1(29603) <= 437480;
srom_1(29604) <= 273143;
srom_1(29605) <= 146862;
srom_1(29606) <= 59230;
srom_1(29607) <= 10657;
srom_1(29608) <= 1371;
srom_1(29609) <= 31415;
srom_1(29610) <= 100650;
srom_1(29611) <= 208749;
srom_1(29612) <= 355207;
srom_1(29613) <= 539336;
srom_1(29614) <= 760272;
srom_1(29615) <= 1016981;
srom_1(29616) <= 1308258;
srom_1(29617) <= 1632737;
srom_1(29618) <= 1988897;
srom_1(29619) <= 2375067;
srom_1(29620) <= 2789437;
srom_1(29621) <= 3230063;
srom_1(29622) <= 3694879;
srom_1(29623) <= 4181706;
srom_1(29624) <= 4688260;
srom_1(29625) <= 5212167;
srom_1(29626) <= 5750969;
srom_1(29627) <= 6302139;
srom_1(29628) <= 6863094;
srom_1(29629) <= 7431203;
srom_1(29630) <= 8003801;
srom_1(29631) <= 8578204;
srom_1(29632) <= 9151717;
srom_1(29633) <= 9721652;
srom_1(29634) <= 10285336;
srom_1(29635) <= 10840126;
srom_1(29636) <= 11383419;
srom_1(29637) <= 11912669;
srom_1(29638) <= 12425393;
srom_1(29639) <= 12919188;
srom_1(29640) <= 13391737;
srom_1(29641) <= 13840824;
srom_1(29642) <= 14264345;
srom_1(29643) <= 14660312;
srom_1(29644) <= 15026868;
srom_1(29645) <= 15362296;
srom_1(29646) <= 15665021;
srom_1(29647) <= 15933625;
srom_1(29648) <= 16166848;
srom_1(29649) <= 16363596;
srom_1(29650) <= 16522947;
srom_1(29651) <= 16644152;
srom_1(29652) <= 16726645;
srom_1(29653) <= 16770038;
srom_1(29654) <= 16774127;
srom_1(29655) <= 16738894;
srom_1(29656) <= 16664503;
srom_1(29657) <= 16551304;
srom_1(29658) <= 16399827;
srom_1(29659) <= 16210783;
srom_1(29660) <= 15985058;
srom_1(29661) <= 15723711;
srom_1(29662) <= 15427966;
srom_1(29663) <= 15099212;
srom_1(29664) <= 14738989;
srom_1(29665) <= 14348988;
srom_1(29666) <= 13931036;
srom_1(29667) <= 13487093;
srom_1(29668) <= 13019243;
srom_1(29669) <= 12529677;
srom_1(29670) <= 12020693;
srom_1(29671) <= 11494676;
srom_1(29672) <= 10954094;
srom_1(29673) <= 10401482;
srom_1(29674) <= 9839430;
srom_1(29675) <= 9270575;
srom_1(29676) <= 8697585;
srom_1(29677) <= 8123145;
srom_1(29678) <= 7549950;
srom_1(29679) <= 6980688;
srom_1(29680) <= 6418028;
srom_1(29681) <= 5864609;
srom_1(29682) <= 5323026;
srom_1(29683) <= 4795818;
srom_1(29684) <= 4285458;
srom_1(29685) <= 3794339;
srom_1(29686) <= 3324765;
srom_1(29687) <= 2878936;
srom_1(29688) <= 2458944;
srom_1(29689) <= 2066759;
srom_1(29690) <= 1704218;
srom_1(29691) <= 1373023;
srom_1(29692) <= 1074727;
srom_1(29693) <= 810728;
srom_1(29694) <= 582264;
srom_1(29695) <= 390407;
srom_1(29696) <= 236056;
srom_1(29697) <= 119935;
srom_1(29698) <= 42589;
srom_1(29699) <= 4380;
srom_1(29700) <= 5487;
srom_1(29701) <= 45906;
srom_1(29702) <= 125447;
srom_1(29703) <= 243737;
srom_1(29704) <= 400221;
srom_1(29705) <= 594164;
srom_1(29706) <= 824659;
srom_1(29707) <= 1090624;
srom_1(29708) <= 1390811;
srom_1(29709) <= 1723814;
srom_1(29710) <= 2088070;
srom_1(29711) <= 2481871;
srom_1(29712) <= 2903372;
srom_1(29713) <= 3350594;
srom_1(29714) <= 3821441;
srom_1(29715) <= 4313705;
srom_1(29716) <= 4825078;
srom_1(29717) <= 5353162;
srom_1(29718) <= 5895479;
srom_1(29719) <= 6449488;
srom_1(29720) <= 7012590;
srom_1(29721) <= 7582145;
srom_1(29722) <= 8155481;
srom_1(29723) <= 8729911;
srom_1(29724) <= 9302740;
srom_1(29725) <= 9871283;
srom_1(29726) <= 10432872;
srom_1(29727) <= 10984876;
srom_1(29728) <= 11524704;
srom_1(29729) <= 12049827;
srom_1(29730) <= 12557780;
srom_1(29731) <= 13046183;
srom_1(29732) <= 13512745;
srom_1(29733) <= 13955278;
srom_1(29734) <= 14371707;
srom_1(29735) <= 14760080;
srom_1(29736) <= 15118574;
srom_1(29737) <= 15445509;
srom_1(29738) <= 15739352;
srom_1(29739) <= 15998725;
srom_1(29740) <= 16222411;
srom_1(29741) <= 16409362;
srom_1(29742) <= 16558701;
srom_1(29743) <= 16669727;
srom_1(29744) <= 16741920;
srom_1(29745) <= 16774942;
srom_1(29746) <= 16768638;
srom_1(29747) <= 16723036;
srom_1(29748) <= 16638352;
srom_1(29749) <= 16514982;
srom_1(29750) <= 16353504;
srom_1(29751) <= 16154676;
srom_1(29752) <= 15919430;
srom_1(29753) <= 15648870;
srom_1(29754) <= 15344264;
srom_1(29755) <= 15007041;
srom_1(29756) <= 14638781;
srom_1(29757) <= 14241212;
srom_1(29758) <= 13816198;
srom_1(29759) <= 13365733;
srom_1(29760) <= 12891928;
srom_1(29761) <= 12397005;
srom_1(29762) <= 11883285;
srom_1(29763) <= 11353178;
srom_1(29764) <= 10809169;
srom_1(29765) <= 10253809;
srom_1(29766) <= 9689703;
srom_1(29767) <= 9119495;
srom_1(29768) <= 8545860;
srom_1(29769) <= 7971487;
srom_1(29770) <= 7399071;
srom_1(29771) <= 6831294;
srom_1(29772) <= 6270821;
srom_1(29773) <= 5720278;
srom_1(29774) <= 5182248;
srom_1(29775) <= 4659254;
srom_1(29776) <= 4153749;
srom_1(29777) <= 3668101;
srom_1(29778) <= 3204590;
srom_1(29779) <= 2765389;
srom_1(29780) <= 2352557;
srom_1(29781) <= 1968029;
srom_1(29782) <= 1613610;
srom_1(29783) <= 1290962;
srom_1(29784) <= 1001597;
srom_1(29785) <= 746872;
srom_1(29786) <= 527981;
srom_1(29787) <= 345952;
srom_1(29788) <= 201638;
srom_1(29789) <= 95715;
srom_1(29790) <= 28680;
srom_1(29791) <= 848;
srom_1(29792) <= 12349;
srom_1(29793) <= 63129;
srom_1(29794) <= 152950;
srom_1(29795) <= 281391;
srom_1(29796) <= 447850;
srom_1(29797) <= 651545;
srom_1(29798) <= 891522;
srom_1(29799) <= 1166656;
srom_1(29800) <= 1475656;
srom_1(29801) <= 1817073;
srom_1(29802) <= 2189306;
srom_1(29803) <= 2590610;
srom_1(29804) <= 3019102;
srom_1(29805) <= 3472774;
srom_1(29806) <= 3949498;
srom_1(29807) <= 4447039;
srom_1(29808) <= 4963063;
srom_1(29809) <= 5495150;
srom_1(29810) <= 6040806;
srom_1(29811) <= 6597472;
srom_1(29812) <= 7162537;
srom_1(29813) <= 7733351;
srom_1(29814) <= 8307238;
srom_1(29815) <= 8881507;
srom_1(29816) <= 9453464;
srom_1(29817) <= 10020427;
srom_1(29818) <= 10579739;
srom_1(29819) <= 11128775;
srom_1(29820) <= 11664962;
srom_1(29821) <= 12185785;
srom_1(29822) <= 12688802;
srom_1(29823) <= 13171654;
srom_1(29824) <= 13632076;
srom_1(29825) <= 14067910;
srom_1(29826) <= 14477111;
srom_1(29827) <= 14857762;
srom_1(29828) <= 15208076;
srom_1(29829) <= 15526412;
srom_1(29830) <= 15811276;
srom_1(29831) <= 16061333;
srom_1(29832) <= 16275409;
srom_1(29833) <= 16452502;
srom_1(29834) <= 16591780;
srom_1(29835) <= 16692591;
srom_1(29836) <= 16754461;
srom_1(29837) <= 16777101;
srom_1(29838) <= 16760405;
srom_1(29839) <= 16704450;
srom_1(29840) <= 16609499;
srom_1(29841) <= 16475998;
srom_1(29842) <= 16304573;
srom_1(29843) <= 16096026;
srom_1(29844) <= 15851337;
srom_1(29845) <= 15571653;
srom_1(29846) <= 15258285;
srom_1(29847) <= 14912702;
srom_1(29848) <= 14536526;
srom_1(29849) <= 14131520;
srom_1(29850) <= 13699584;
srom_1(29851) <= 13242742;
srom_1(29852) <= 12763138;
srom_1(29853) <= 12263020;
srom_1(29854) <= 11744734;
srom_1(29855) <= 11210710;
srom_1(29856) <= 10663452;
srom_1(29857) <= 10105526;
srom_1(29858) <= 9539549;
srom_1(29859) <= 8968175;
srom_1(29860) <= 8394084;
srom_1(29861) <= 7819966;
srom_1(29862) <= 7248515;
srom_1(29863) <= 6682410;
srom_1(29864) <= 6124307;
srom_1(29865) <= 5576821;
srom_1(29866) <= 5042521;
srom_1(29867) <= 4523912;
srom_1(29868) <= 4023425;
srom_1(29869) <= 3543409;
srom_1(29870) <= 3086113;
srom_1(29871) <= 2653682;
srom_1(29872) <= 2248145;
srom_1(29873) <= 1871402;
srom_1(29874) <= 1525221;
srom_1(29875) <= 1211224;
srom_1(29876) <= 930885;
srom_1(29877) <= 685517;
srom_1(29878) <= 476272;
srom_1(29879) <= 304131;
srom_1(29880) <= 169900;
srom_1(29881) <= 74210;
srom_1(29882) <= 17509;
srom_1(29883) <= 62;
srom_1(29884) <= 21953;
srom_1(29885) <= 83078;
srom_1(29886) <= 183150;
srom_1(29887) <= 321700;
srom_1(29888) <= 498079;
srom_1(29889) <= 711459;
srom_1(29890) <= 960840;
srom_1(29891) <= 1245052;
srom_1(29892) <= 1562763;
srom_1(29893) <= 1912483;
srom_1(29894) <= 2292571;
srom_1(29895) <= 2701246;
srom_1(29896) <= 3136591;
srom_1(29897) <= 3596564;
srom_1(29898) <= 4079009;
srom_1(29899) <= 4581663;
srom_1(29900) <= 5102169;
srom_1(29901) <= 5638087;
srom_1(29902) <= 6186902;
srom_1(29903) <= 6746042;
srom_1(29904) <= 7312885;
srom_1(29905) <= 7884772;
srom_1(29906) <= 8459021;
srom_1(29907) <= 9032941;
srom_1(29908) <= 9603839;
srom_1(29909) <= 10169038;
srom_1(29910) <= 10725888;
srom_1(29911) <= 11271778;
srom_1(29912) <= 11804148;
srom_1(29913) <= 12320501;
srom_1(29914) <= 12818416;
srom_1(29915) <= 13295558;
srom_1(29916) <= 13749690;
srom_1(29917) <= 14178682;
srom_1(29918) <= 14580522;
srom_1(29919) <= 14953326;
srom_1(29920) <= 15295346;
srom_1(29921) <= 15604978;
srom_1(29922) <= 15880770;
srom_1(29923) <= 16121428;
srom_1(29924) <= 16325825;
srom_1(29925) <= 16493001;
srom_1(29926) <= 16622173;
srom_1(29927) <= 16712735;
srom_1(29928) <= 16764263;
srom_1(29929) <= 16776514;
srom_1(29930) <= 16749431;
srom_1(29931) <= 16683141;
srom_1(29932) <= 16577956;
srom_1(29933) <= 16434367;
srom_1(29934) <= 16253050;
srom_1(29935) <= 16034853;
srom_1(29936) <= 15780801;
srom_1(29937) <= 15492084;
srom_1(29938) <= 15170056;
srom_1(29939) <= 14816228;
srom_1(29940) <= 14432258;
srom_1(29941) <= 14019948;
srom_1(29942) <= 13581230;
srom_1(29943) <= 13118163;
srom_1(29944) <= 12632917;
srom_1(29945) <= 12127768;
srom_1(29946) <= 11605084;
srom_1(29947) <= 11067318;
srom_1(29948) <= 10516990;
srom_1(29949) <= 9956681;
srom_1(29950) <= 9389019;
srom_1(29951) <= 8816666;
srom_1(29952) <= 8242306;
srom_1(29953) <= 7668631;
srom_1(29954) <= 7098333;
srom_1(29955) <= 6534085;
srom_1(29956) <= 5978534;
srom_1(29957) <= 5434285;
srom_1(29958) <= 4903889;
srom_1(29959) <= 4389834;
srom_1(29960) <= 3894531;
srom_1(29961) <= 3420302;
srom_1(29962) <= 2969372;
srom_1(29963) <= 2543854;
srom_1(29964) <= 2145744;
srom_1(29965) <= 1776909;
srom_1(29966) <= 1439078;
srom_1(29967) <= 1133836;
srom_1(29968) <= 862615;
srom_1(29969) <= 626685;
srom_1(29970) <= 427153;
srom_1(29971) <= 264956;
srom_1(29972) <= 140853;
srom_1(29973) <= 55427;
srom_1(29974) <= 9078;
srom_1(29975) <= 2023;
srom_1(29976) <= 34296;
srom_1(29977) <= 105745;
srom_1(29978) <= 216035;
srom_1(29979) <= 364650;
srom_1(29980) <= 550891;
srom_1(29981) <= 773886;
srom_1(29982) <= 1032589;
srom_1(29983) <= 1325788;
srom_1(29984) <= 1652106;
srom_1(29985) <= 2010013;
srom_1(29986) <= 2397833;
srom_1(29987) <= 2813745;
srom_1(29988) <= 3255799;
srom_1(29989) <= 3721923;
srom_1(29990) <= 4209931;
srom_1(29991) <= 4717534;
srom_1(29992) <= 5242352;
srom_1(29993) <= 5781923;
srom_1(29994) <= 6333719;
srom_1(29995) <= 6895150;
srom_1(29996) <= 7463585;
srom_1(29997) <= 8036357;
srom_1(29998) <= 8610782;
srom_1(29999) <= 9184164;
srom_1(30000) <= 9753816;
srom_1(30001) <= 10317066;
srom_1(30002) <= 10871272;
srom_1(30003) <= 11413837;
srom_1(30004) <= 11942215;
srom_1(30005) <= 12453929;
srom_1(30006) <= 12946580;
srom_1(30007) <= 13417856;
srom_1(30008) <= 13865549;
srom_1(30009) <= 14287558;
srom_1(30010) <= 14681906;
srom_1(30011) <= 15046741;
srom_1(30012) <= 15380355;
srom_1(30013) <= 15681182;
srom_1(30014) <= 15947811;
srom_1(30015) <= 16178993;
srom_1(30016) <= 16373643;
srom_1(30017) <= 16530848;
srom_1(30018) <= 16649871;
srom_1(30019) <= 16730155;
srom_1(30020) <= 16771322;
srom_1(30021) <= 16773180;
srom_1(30022) <= 16735720;
srom_1(30023) <= 16659117;
srom_1(30024) <= 16543731;
srom_1(30025) <= 16390102;
srom_1(30026) <= 16198952;
srom_1(30027) <= 15971177;
srom_1(30028) <= 15707844;
srom_1(30029) <= 15410189;
srom_1(30030) <= 15079607;
srom_1(30031) <= 14717649;
srom_1(30032) <= 14326012;
srom_1(30033) <= 13906532;
srom_1(30034) <= 13461177;
srom_1(30035) <= 12992035;
srom_1(30036) <= 12501306;
srom_1(30037) <= 11991290;
srom_1(30038) <= 11464381;
srom_1(30039) <= 10923048;
srom_1(30040) <= 10369831;
srom_1(30041) <= 9807323;
srom_1(30042) <= 9238161;
srom_1(30043) <= 8665017;
srom_1(30044) <= 8090575;
srom_1(30045) <= 7517532;
srom_1(30046) <= 6948573;
srom_1(30047) <= 6386367;
srom_1(30048) <= 5833550;
srom_1(30049) <= 5292715;
srom_1(30050) <= 4766398;
srom_1(30051) <= 4257066;
srom_1(30052) <= 3767108;
srom_1(30053) <= 3298823;
srom_1(30054) <= 2854405;
srom_1(30055) <= 2435938;
srom_1(30056) <= 2045386;
srom_1(30057) <= 1684580;
srom_1(30058) <= 1355211;
srom_1(30059) <= 1058823;
srom_1(30060) <= 796808;
srom_1(30061) <= 570394;
srom_1(30062) <= 380641;
srom_1(30063) <= 228441;
srom_1(30064) <= 114506;
srom_1(30065) <= 39372;
srom_1(30066) <= 3390;
srom_1(30067) <= 6729;
srom_1(30068) <= 49374;
srom_1(30069) <= 131124;
srom_1(30070) <= 251597;
srom_1(30071) <= 410226;
srom_1(30072) <= 606269;
srom_1(30073) <= 838807;
srom_1(30074) <= 1106747;
srom_1(30075) <= 1408835;
srom_1(30076) <= 1743653;
srom_1(30077) <= 2109632;
srom_1(30078) <= 2505055;
srom_1(30079) <= 2928068;
srom_1(30080) <= 3376688;
srom_1(30081) <= 3848810;
srom_1(30082) <= 4342221;
srom_1(30083) <= 4854606;
srom_1(30084) <= 5383564;
srom_1(30085) <= 5926613;
srom_1(30086) <= 6481208;
srom_1(30087) <= 7044747;
srom_1(30088) <= 7614588;
srom_1(30089) <= 8188058;
srom_1(30090) <= 8762469;
srom_1(30091) <= 9335127;
srom_1(30092) <= 9903346;
srom_1(30093) <= 10464462;
srom_1(30094) <= 11015844;
srom_1(30095) <= 11554905;
srom_1(30096) <= 12079119;
srom_1(30097) <= 12586027;
srom_1(30098) <= 13073251;
srom_1(30099) <= 13538508;
srom_1(30100) <= 13979615;
srom_1(30101) <= 14394504;
srom_1(30102) <= 14781229;
srom_1(30103) <= 15137977;
srom_1(30104) <= 15463074;
srom_1(30105) <= 15754998;
srom_1(30106) <= 16012377;
srom_1(30107) <= 16234006;
srom_1(30108) <= 16418846;
srom_1(30109) <= 16566029;
srom_1(30110) <= 16674865;
srom_1(30111) <= 16744844;
srom_1(30112) <= 16775637;
srom_1(30113) <= 16767101;
srom_1(30114) <= 16719276;
srom_1(30115) <= 16632385;
srom_1(30116) <= 16506836;
srom_1(30117) <= 16343218;
srom_1(30118) <= 16142298;
srom_1(30119) <= 15905018;
srom_1(30120) <= 15632491;
srom_1(30121) <= 15325996;
srom_1(30122) <= 14986968;
srom_1(30123) <= 14616998;
srom_1(30124) <= 14217822;
srom_1(30125) <= 13791310;
srom_1(30126) <= 13339463;
srom_1(30127) <= 12864400;
srom_1(30128) <= 12368348;
srom_1(30129) <= 11853634;
srom_1(30130) <= 11322671;
srom_1(30131) <= 10777949;
srom_1(30132) <= 10222023;
srom_1(30133) <= 9657500;
srom_1(30134) <= 9087026;
srom_1(30135) <= 8513277;
srom_1(30136) <= 7938943;
srom_1(30137) <= 7366718;
srom_1(30138) <= 6799285;
srom_1(30139) <= 6239305;
srom_1(30140) <= 5689403;
srom_1(30141) <= 5152159;
srom_1(30142) <= 4630092;
srom_1(30143) <= 4125650;
srom_1(30144) <= 3641199;
srom_1(30145) <= 3179009;
srom_1(30146) <= 2741249;
srom_1(30147) <= 2329972;
srom_1(30148) <= 1947106;
srom_1(30149) <= 1594446;
srom_1(30150) <= 1273646;
srom_1(30151) <= 986210;
srom_1(30152) <= 733487;
srom_1(30153) <= 516662;
srom_1(30154) <= 336751;
srom_1(30155) <= 194597;
srom_1(30156) <= 90869;
srom_1(30157) <= 26051;
srom_1(30158) <= 448;
srom_1(30159) <= 14180;
srom_1(30160) <= 67182;
srom_1(30161) <= 159207;
srom_1(30162) <= 289822;
srom_1(30163) <= 458415;
srom_1(30164) <= 664196;
srom_1(30165) <= 906198;
srom_1(30166) <= 1183289;
srom_1(30167) <= 1494168;
srom_1(30168) <= 1837377;
srom_1(30169) <= 2211307;
srom_1(30170) <= 2614204;
srom_1(30171) <= 3044180;
srom_1(30172) <= 3499217;
srom_1(30173) <= 3977183;
srom_1(30174) <= 4475835;
srom_1(30175) <= 4992836;
srom_1(30176) <= 5525760;
srom_1(30177) <= 6072109;
srom_1(30178) <= 6629322;
srom_1(30179) <= 7194784;
srom_1(30180) <= 7765844;
srom_1(30181) <= 8339825;
srom_1(30182) <= 8914034;
srom_1(30183) <= 9485780;
srom_1(30184) <= 10052380;
srom_1(30185) <= 10611179;
srom_1(30186) <= 11159555;
srom_1(30187) <= 11694937;
srom_1(30188) <= 12214815;
srom_1(30189) <= 12716750;
srom_1(30190) <= 13198389;
srom_1(30191) <= 13657473;
srom_1(30192) <= 14091850;
srom_1(30193) <= 14499483;
srom_1(30194) <= 14878459;
srom_1(30195) <= 15227002;
srom_1(30196) <= 15543478;
srom_1(30197) <= 15826402;
srom_1(30198) <= 16074447;
srom_1(30199) <= 16286452;
srom_1(30200) <= 16461420;
srom_1(30201) <= 16598532;
srom_1(30202) <= 16697145;
srom_1(30203) <= 16756796;
srom_1(30204) <= 16777207;
srom_1(30205) <= 16758280;
srom_1(30206) <= 16700104;
srom_1(30207) <= 16602954;
srom_1(30208) <= 16467283;
srom_1(30209) <= 16293729;
srom_1(30210) <= 16083105;
srom_1(30211) <= 15836398;
srom_1(30212) <= 15554767;
srom_1(30213) <= 15239531;
srom_1(30214) <= 14892168;
srom_1(30215) <= 14514309;
srom_1(30216) <= 14107723;
srom_1(30217) <= 13674319;
srom_1(30218) <= 13216128;
srom_1(30219) <= 12735299;
srom_1(30220) <= 12234088;
srom_1(30221) <= 11714843;
srom_1(30222) <= 11180000;
srom_1(30223) <= 10632068;
srom_1(30224) <= 10073615;
srom_1(30225) <= 9507261;
srom_1(30226) <= 8935661;
srom_1(30227) <= 8361496;
srom_1(30228) <= 7787458;
srom_1(30229) <= 7216238;
srom_1(30230) <= 6650517;
srom_1(30231) <= 6092946;
srom_1(30232) <= 5546140;
srom_1(30233) <= 5012663;
srom_1(30234) <= 4495017;
srom_1(30235) <= 3995630;
srom_1(30236) <= 3516843;
srom_1(30237) <= 3060901;
srom_1(30238) <= 2629943;
srom_1(30239) <= 2225989;
srom_1(30240) <= 1850934;
srom_1(30241) <= 1506536;
srom_1(30242) <= 1194410;
srom_1(30243) <= 916021;
srom_1(30244) <= 672673;
srom_1(30245) <= 465508;
srom_1(30246) <= 295496;
srom_1(30247) <= 163437;
srom_1(30248) <= 69947;
srom_1(30249) <= 15467;
srom_1(30250) <= 252;
srom_1(30251) <= 24372;
srom_1(30252) <= 87715;
srom_1(30253) <= 189984;
srom_1(30254) <= 330699;
srom_1(30255) <= 509200;
srom_1(30256) <= 724651;
srom_1(30257) <= 976040;
srom_1(30258) <= 1262190;
srom_1(30259) <= 1581757;
srom_1(30260) <= 1933245;
srom_1(30261) <= 2315004;
srom_1(30262) <= 2725244;
srom_1(30263) <= 3162041;
srom_1(30264) <= 3623348;
srom_1(30265) <= 4107000;
srom_1(30266) <= 4610731;
srom_1(30267) <= 5132177;
srom_1(30268) <= 5668894;
srom_1(30269) <= 6218364;
srom_1(30270) <= 6778011;
srom_1(30271) <= 7345211;
srom_1(30272) <= 7917304;
srom_1(30273) <= 8491607;
srom_1(30274) <= 9065427;
srom_1(30275) <= 9636074;
srom_1(30276) <= 10200870;
srom_1(30277) <= 10757168;
srom_1(30278) <= 11302359;
srom_1(30279) <= 11833886;
srom_1(30280) <= 12349258;
srom_1(30281) <= 12846056;
srom_1(30282) <= 13321952;
srom_1(30283) <= 13774714;
srom_1(30284) <= 14202218;
srom_1(30285) <= 14602461;
srom_1(30286) <= 14973564;
srom_1(30287) <= 15313789;
srom_1(30288) <= 15621539;
srom_1(30289) <= 15895371;
srom_1(30290) <= 16134001;
srom_1(30291) <= 16336311;
srom_1(30292) <= 16501351;
srom_1(30293) <= 16628348;
srom_1(30294) <= 16716705;
srom_1(30295) <= 16766010;
srom_1(30296) <= 16776029;
srom_1(30297) <= 16746718;
srom_1(30298) <= 16678212;
srom_1(30299) <= 16570833;
srom_1(30300) <= 16425085;
srom_1(30301) <= 16241652;
srom_1(30302) <= 16021393;
srom_1(30303) <= 15765340;
srom_1(30304) <= 15474696;
srom_1(30305) <= 15150823;
srom_1(30306) <= 14795240;
srom_1(30307) <= 14409613;
srom_1(30308) <= 13995752;
srom_1(30309) <= 13555597;
srom_1(30310) <= 13091213;
srom_1(30311) <= 12604776;
srom_1(30312) <= 12098568;
srom_1(30313) <= 11574963;
srom_1(30314) <= 11036416;
srom_1(30315) <= 10485452;
srom_1(30316) <= 9924656;
srom_1(30317) <= 9356656;
srom_1(30318) <= 8784118;
srom_1(30319) <= 8209724;
srom_1(30320) <= 7636169;
srom_1(30321) <= 7066143;
srom_1(30322) <= 6502318;
srom_1(30323) <= 5947338;
srom_1(30324) <= 5403807;
srom_1(30325) <= 4874272;
srom_1(30326) <= 4361217;
srom_1(30327) <= 3867048;
srom_1(30328) <= 3394083;
srom_1(30329) <= 2944538;
srom_1(30330) <= 2520522;
srom_1(30331) <= 2124024;
srom_1(30332) <= 1756902;
srom_1(30333) <= 1420879;
srom_1(30334) <= 1117530;
srom_1(30335) <= 848278;
srom_1(30336) <= 614384;
srom_1(30337) <= 416947;
srom_1(30338) <= 256892;
srom_1(30339) <= 134969;
srom_1(30340) <= 51750;
srom_1(30341) <= 7625;
srom_1(30342) <= 2802;
srom_1(30343) <= 37303;
srom_1(30344) <= 110966;
srom_1(30345) <= 223445;
srom_1(30346) <= 374214;
srom_1(30347) <= 562565;
srom_1(30348) <= 787615;
srom_1(30349) <= 1048309;
srom_1(30350) <= 1343424;
srom_1(30351) <= 1671576;
srom_1(30352) <= 2031226;
srom_1(30353) <= 2420689;
srom_1(30354) <= 2838137;
srom_1(30355) <= 3281613;
srom_1(30356) <= 3749038;
srom_1(30357) <= 4238219;
srom_1(30358) <= 4746863;
srom_1(30359) <= 5272584;
srom_1(30360) <= 5812917;
srom_1(30361) <= 6365329;
srom_1(30362) <= 6927228;
srom_1(30363) <= 7495981;
srom_1(30364) <= 8068919;
srom_1(30365) <= 8643356;
srom_1(30366) <= 9216599;
srom_1(30367) <= 9785959;
srom_1(30368) <= 10348766;
srom_1(30369) <= 10902382;
srom_1(30370) <= 11444209;
srom_1(30371) <= 11971708;
srom_1(30372) <= 12482404;
srom_1(30373) <= 12973903;
srom_1(30374) <= 13443900;
srom_1(30375) <= 13890191;
srom_1(30376) <= 14310683;
srom_1(30377) <= 14703405;
srom_1(30378) <= 15066514;
srom_1(30379) <= 15398308;
srom_1(30380) <= 15697232;
srom_1(30381) <= 15961883;
srom_1(30382) <= 16191020;
srom_1(30383) <= 16383568;
srom_1(30384) <= 16538626;
srom_1(30385) <= 16655466;
srom_1(30386) <= 16733539;
srom_1(30387) <= 16772480;
srom_1(30388) <= 16772106;
srom_1(30389) <= 16732419;
srom_1(30390) <= 16653605;
srom_1(30391) <= 16536034;
srom_1(30392) <= 16380257;
srom_1(30393) <= 16187004;
srom_1(30394) <= 15957181;
srom_1(30395) <= 15691867;
srom_1(30396) <= 15392306;
srom_1(30397) <= 15059902;
srom_1(30398) <= 14696213;
srom_1(30399) <= 14302947;
srom_1(30400) <= 13881945;
srom_1(30401) <= 13435184;
srom_1(30402) <= 12964758;
srom_1(30403) <= 12472872;
srom_1(30404) <= 11961834;
srom_1(30405) <= 11434040;
srom_1(30406) <= 10891964;
srom_1(30407) <= 10338150;
srom_1(30408) <= 9775194;
srom_1(30409) <= 9205735;
srom_1(30410) <= 8632444;
srom_1(30411) <= 8058011;
srom_1(30412) <= 7485127;
srom_1(30413) <= 6916480;
srom_1(30414) <= 6354736;
srom_1(30415) <= 5802530;
srom_1(30416) <= 5262451;
srom_1(30417) <= 4737032;
srom_1(30418) <= 4228736;
srom_1(30419) <= 3739947;
srom_1(30420) <= 3272957;
srom_1(30421) <= 2829956;
srom_1(30422) <= 2413022;
srom_1(30423) <= 2024109;
srom_1(30424) <= 1665042;
srom_1(30425) <= 1337504;
srom_1(30426) <= 1043031;
srom_1(30427) <= 783003;
srom_1(30428) <= 558641;
srom_1(30429) <= 370996;
srom_1(30430) <= 220949;
srom_1(30431) <= 109203;
srom_1(30432) <= 36281;
srom_1(30433) <= 2527;
srom_1(30434) <= 8098;
srom_1(30435) <= 52967;
srom_1(30436) <= 136926;
srom_1(30437) <= 259579;
srom_1(30438) <= 420353;
srom_1(30439) <= 618492;
srom_1(30440) <= 853068;
srom_1(30441) <= 1122980;
srom_1(30442) <= 1426964;
srom_1(30443) <= 1763593;
srom_1(30444) <= 2131289;
srom_1(30445) <= 2528328;
srom_1(30446) <= 2952848;
srom_1(30447) <= 3402858;
srom_1(30448) <= 3876247;
srom_1(30449) <= 4370797;
srom_1(30450) <= 4884188;
srom_1(30451) <= 5414012;
srom_1(30452) <= 5957785;
srom_1(30453) <= 6512956;
srom_1(30454) <= 7076924;
srom_1(30455) <= 7647042;
srom_1(30456) <= 8220638;
srom_1(30457) <= 8795022;
srom_1(30458) <= 9367499;
srom_1(30459) <= 9935387;
srom_1(30460) <= 10496021;
srom_1(30461) <= 11046772;
srom_1(30462) <= 11585059;
srom_1(30463) <= 12108356;
srom_1(30464) <= 12614210;
srom_1(30465) <= 13100249;
srom_1(30466) <= 13564193;
srom_1(30467) <= 14003867;
srom_1(30468) <= 14417209;
srom_1(30469) <= 14802281;
srom_1(30470) <= 15157277;
srom_1(30471) <= 15480533;
srom_1(30472) <= 15770532;
srom_1(30473) <= 16025915;
srom_1(30474) <= 16245483;
srom_1(30475) <= 16428208;
srom_1(30476) <= 16573233;
srom_1(30477) <= 16679877;
srom_1(30478) <= 16747641;
srom_1(30479) <= 16776206;
srom_1(30480) <= 16765438;
srom_1(30481) <= 16715389;
srom_1(30482) <= 16626293;
srom_1(30483) <= 16498568;
srom_1(30484) <= 16332812;
srom_1(30485) <= 16129803;
srom_1(30486) <= 15890492;
srom_1(30487) <= 15616003;
srom_1(30488) <= 15307622;
srom_1(30489) <= 14966796;
srom_1(30490) <= 14595122;
srom_1(30491) <= 14194344;
srom_1(30492) <= 13766340;
srom_1(30493) <= 13313119;
srom_1(30494) <= 12836804;
srom_1(30495) <= 12339631;
srom_1(30496) <= 11823930;
srom_1(30497) <= 11292119;
srom_1(30498) <= 10746693;
srom_1(30499) <= 10190209;
srom_1(30500) <= 9625277;
srom_1(30501) <= 9054546;
srom_1(30502) <= 8480691;
srom_1(30503) <= 7906405;
srom_1(30504) <= 7334381;
srom_1(30505) <= 6767299;
srom_1(30506) <= 6207821;
srom_1(30507) <= 5658569;
srom_1(30508) <= 5122119;
srom_1(30509) <= 4600987;
srom_1(30510) <= 4097616;
srom_1(30511) <= 3614367;
srom_1(30512) <= 3153507;
srom_1(30513) <= 2717195;
srom_1(30514) <= 2307479;
srom_1(30515) <= 1926279;
srom_1(30516) <= 1575383;
srom_1(30517) <= 1256437;
srom_1(30518) <= 970936;
srom_1(30519) <= 720219;
srom_1(30520) <= 505461;
srom_1(30521) <= 327671;
srom_1(30522) <= 187681;
srom_1(30523) <= 86148;
srom_1(30524) <= 23548;
srom_1(30525) <= 174;
srom_1(30526) <= 16137;
srom_1(30527) <= 71361;
srom_1(30528) <= 165588;
srom_1(30529) <= 298375;
srom_1(30530) <= 469100;
srom_1(30531) <= 676963;
srom_1(30532) <= 920988;
srom_1(30533) <= 1200031;
srom_1(30534) <= 1512784;
srom_1(30535) <= 1857779;
srom_1(30536) <= 2233401;
srom_1(30537) <= 2637886;
srom_1(30538) <= 3069338;
srom_1(30539) <= 3525734;
srom_1(30540) <= 4004934;
srom_1(30541) <= 4504690;
srom_1(30542) <= 5022660;
srom_1(30543) <= 5556413;
srom_1(30544) <= 6103448;
srom_1(30545) <= 6661198;
srom_1(30546) <= 7227049;
srom_1(30547) <= 7798347;
srom_1(30548) <= 8372412;
srom_1(30549) <= 8946554;
srom_1(30550) <= 9518079;
srom_1(30551) <= 10084308;
srom_1(30552) <= 10642585;
srom_1(30553) <= 11190293;
srom_1(30554) <= 11724862;
srom_1(30555) <= 12243786;
srom_1(30556) <= 12744632;
srom_1(30557) <= 13225052;
srom_1(30558) <= 13682791;
srom_1(30559) <= 14115705;
srom_1(30560) <= 14521762;
srom_1(30561) <= 14899058;
srom_1(30562) <= 15245825;
srom_1(30563) <= 15560436;
srom_1(30564) <= 15841415;
srom_1(30565) <= 16087446;
srom_1(30566) <= 16297375;
srom_1(30567) <= 16470216;
srom_1(30568) <= 16605160;
srom_1(30569) <= 16701574;
srom_1(30570) <= 16759006;
srom_1(30571) <= 16777185;
srom_1(30572) <= 16756028;
srom_1(30573) <= 16695633;
srom_1(30574) <= 16596284;
srom_1(30575) <= 16458446;
srom_1(30576) <= 16282766;
srom_1(30577) <= 16070067;
srom_1(30578) <= 15821347;
srom_1(30579) <= 15537773;
srom_1(30580) <= 15220674;
srom_1(30581) <= 14871537;
srom_1(30582) <= 14491999;
srom_1(30583) <= 14083840;
srom_1(30584) <= 13648974;
srom_1(30585) <= 13189441;
srom_1(30586) <= 12707395;
srom_1(30587) <= 12205097;
srom_1(30588) <= 11684901;
srom_1(30589) <= 11149249;
srom_1(30590) <= 10600650;
srom_1(30591) <= 10041679;
srom_1(30592) <= 9474956;
srom_1(30593) <= 8903139;
srom_1(30594) <= 8328908;
srom_1(30595) <= 7754958;
srom_1(30596) <= 7183979;
srom_1(30597) <= 6618649;
srom_1(30598) <= 6061619;
srom_1(30599) <= 5515501;
srom_1(30600) <= 4982856;
srom_1(30601) <= 4466182;
srom_1(30602) <= 3967901;
srom_1(30603) <= 3490351;
srom_1(30604) <= 3035770;
srom_1(30605) <= 2606291;
srom_1(30606) <= 2203926;
srom_1(30607) <= 1830564;
srom_1(30608) <= 1487955;
srom_1(30609) <= 1177705;
srom_1(30610) <= 901270;
srom_1(30611) <= 659945;
srom_1(30612) <= 454863;
srom_1(30613) <= 286984;
srom_1(30614) <= 157097;
srom_1(30615) <= 65811;
srom_1(30616) <= 13552;
srom_1(30617) <= 568;
srom_1(30618) <= 26918;
srom_1(30619) <= 92478;
srom_1(30620) <= 196942;
srom_1(30621) <= 339820;
srom_1(30622) <= 520441;
srom_1(30623) <= 737958;
srom_1(30624) <= 991352;
srom_1(30625) <= 1279435;
srom_1(30626) <= 1600854;
srom_1(30627) <= 1954104;
srom_1(30628) <= 2337527;
srom_1(30629) <= 2749326;
srom_1(30630) <= 3187570;
srom_1(30631) <= 3650203;
srom_1(30632) <= 4135056;
srom_1(30633) <= 4639855;
srom_1(30634) <= 5162234;
srom_1(30635) <= 5699742;
srom_1(30636) <= 6249859;
srom_1(30637) <= 6810005;
srom_1(30638) <= 7377554;
srom_1(30639) <= 7949844;
srom_1(30640) <= 8524192;
srom_1(30641) <= 9097904;
srom_1(30642) <= 9668290;
srom_1(30643) <= 10232674;
srom_1(30644) <= 10788412;
srom_1(30645) <= 11332896;
srom_1(30646) <= 11863573;
srom_1(30647) <= 12377955;
srom_1(30648) <= 12873629;
srom_1(30649) <= 13348271;
srom_1(30650) <= 13799656;
srom_1(30651) <= 14225667;
srom_1(30652) <= 14624306;
srom_1(30653) <= 14993703;
srom_1(30654) <= 15332127;
srom_1(30655) <= 15637990;
srom_1(30656) <= 15909859;
srom_1(30657) <= 16146457;
srom_1(30658) <= 16346677;
srom_1(30659) <= 16509578;
srom_1(30660) <= 16634398;
srom_1(30661) <= 16720549;
srom_1(30662) <= 16767630;
srom_1(30663) <= 16775419;
srom_1(30664) <= 16743878;
srom_1(30665) <= 16673158;
srom_1(30666) <= 16563588;
srom_1(30667) <= 16415682;
srom_1(30668) <= 16230135;
srom_1(30669) <= 16007817;
srom_1(30670) <= 15749769;
srom_1(30671) <= 15457202;
srom_1(30672) <= 15131488;
srom_1(30673) <= 14774155;
srom_1(30674) <= 14386877;
srom_1(30675) <= 13971472;
srom_1(30676) <= 13529886;
srom_1(30677) <= 13064192;
srom_1(30678) <= 12576571;
srom_1(30679) <= 12069313;
srom_1(30680) <= 11544794;
srom_1(30681) <= 11005474;
srom_1(30682) <= 10453883;
srom_1(30683) <= 9892608;
srom_1(30684) <= 9324279;
srom_1(30685) <= 8751563;
srom_1(30686) <= 8177145;
srom_1(30687) <= 7603718;
srom_1(30688) <= 7033972;
srom_1(30689) <= 6470579;
srom_1(30690) <= 5916180;
srom_1(30691) <= 5373374;
srom_1(30692) <= 4844709;
srom_1(30693) <= 4332661;
srom_1(30694) <= 3839634;
srom_1(30695) <= 3367938;
srom_1(30696) <= 2919786;
srom_1(30697) <= 2497279;
srom_1(30698) <= 2102398;
srom_1(30699) <= 1736996;
srom_1(30700) <= 1402786;
srom_1(30701) <= 1101334;
srom_1(30702) <= 834055;
srom_1(30703) <= 602201;
srom_1(30704) <= 406861;
srom_1(30705) <= 248950;
srom_1(30706) <= 129209;
srom_1(30707) <= 48198;
srom_1(30708) <= 6299;
srom_1(30709) <= 3708;
srom_1(30710) <= 40436;
srom_1(30711) <= 116311;
srom_1(30712) <= 230978;
srom_1(30713) <= 383899;
srom_1(30714) <= 574357;
srom_1(30715) <= 801458;
srom_1(30716) <= 1064139;
srom_1(30717) <= 1361166;
srom_1(30718) <= 1691147;
srom_1(30719) <= 2052535;
srom_1(30720) <= 2443635;
srom_1(30721) <= 2862613;
srom_1(30722) <= 3307504;
srom_1(30723) <= 3776223;
srom_1(30724) <= 4266570;
srom_1(30725) <= 4776247;
srom_1(30726) <= 5302864;
srom_1(30727) <= 5843950;
srom_1(30728) <= 6396970;
srom_1(30729) <= 6959329;
srom_1(30730) <= 7528390;
srom_1(30731) <= 8101485;
srom_1(30732) <= 8675927;
srom_1(30733) <= 9249021;
srom_1(30734) <= 9818081;
srom_1(30735) <= 10380437;
srom_1(30736) <= 10933453;
srom_1(30737) <= 11474535;
srom_1(30738) <= 12001146;
srom_1(30739) <= 12510817;
srom_1(30740) <= 13001157;
srom_1(30741) <= 13469867;
srom_1(30742) <= 13914750;
srom_1(30743) <= 14333719;
srom_1(30744) <= 14724809;
srom_1(30745) <= 15086186;
srom_1(30746) <= 15416156;
srom_1(30747) <= 15713172;
srom_1(30748) <= 15975840;
srom_1(30749) <= 16202929;
srom_1(30750) <= 16393374;
srom_1(30751) <= 16546281;
srom_1(30752) <= 16660935;
srom_1(30753) <= 16736797;
srom_1(30754) <= 16773511;
srom_1(30755) <= 16770906;
srom_1(30756) <= 16728993;
srom_1(30757) <= 16647969;
srom_1(30758) <= 16528215;
srom_1(30759) <= 16370290;
srom_1(30760) <= 16174937;
srom_1(30761) <= 15943072;
srom_1(30762) <= 15675780;
srom_1(30763) <= 15374317;
srom_1(30764) <= 15040095;
srom_1(30765) <= 14674682;
srom_1(30766) <= 14279792;
srom_1(30767) <= 13857276;
srom_1(30768) <= 13409115;
srom_1(30769) <= 12937411;
srom_1(30770) <= 12444377;
srom_1(30771) <= 11932323;
srom_1(30772) <= 11403652;
srom_1(30773) <= 10860843;
srom_1(30774) <= 10306440;
srom_1(30775) <= 9743044;
srom_1(30776) <= 9173296;
srom_1(30777) <= 8599869;
srom_1(30778) <= 8025451;
srom_1(30779) <= 7452736;
srom_1(30780) <= 6884409;
srom_1(30781) <= 6323136;
srom_1(30782) <= 5771549;
srom_1(30783) <= 5232235;
srom_1(30784) <= 4707721;
srom_1(30785) <= 4200469;
srom_1(30786) <= 3712856;
srom_1(30787) <= 3247169;
srom_1(30788) <= 2805592;
srom_1(30789) <= 2390196;
srom_1(30790) <= 2002929;
srom_1(30791) <= 1645606;
srom_1(30792) <= 1319903;
srom_1(30793) <= 1027348;
srom_1(30794) <= 769313;
srom_1(30795) <= 547007;
srom_1(30796) <= 361473;
srom_1(30797) <= 213581;
srom_1(30798) <= 104024;
srom_1(30799) <= 33317;
srom_1(30800) <= 1790;
srom_1(30801) <= 9592;
srom_1(30802) <= 56687;
srom_1(30803) <= 142852;
srom_1(30804) <= 267685;
srom_1(30805) <= 430599;
srom_1(30806) <= 630832;
srom_1(30807) <= 867443;
srom_1(30808) <= 1139323;
srom_1(30809) <= 1445198;
srom_1(30810) <= 1783633;
srom_1(30811) <= 2153041;
srom_1(30812) <= 2551689;
srom_1(30813) <= 2977709;
srom_1(30814) <= 3429103;
srom_1(30815) <= 3903753;
srom_1(30816) <= 4399434;
srom_1(30817) <= 4913822;
srom_1(30818) <= 5444504;
srom_1(30819) <= 5988992;
srom_1(30820) <= 6544733;
srom_1(30821) <= 7109121;
srom_1(30822) <= 7679508;
srom_1(30823) <= 8253221;
srom_1(30824) <= 8827568;
srom_1(30825) <= 9399857;
srom_1(30826) <= 9967404;
srom_1(30827) <= 10527547;
srom_1(30828) <= 11077660;
srom_1(30829) <= 11615164;
srom_1(30830) <= 12137537;
srom_1(30831) <= 12642329;
srom_1(30832) <= 13127175;
srom_1(30833) <= 13589800;
srom_1(30834) <= 14028034;
srom_1(30835) <= 14439824;
srom_1(30836) <= 14823237;
srom_1(30837) <= 15176476;
srom_1(30838) <= 15497884;
srom_1(30839) <= 15785955;
srom_1(30840) <= 16039337;
srom_1(30841) <= 16256842;
srom_1(30842) <= 16437450;
srom_1(30843) <= 16580314;
srom_1(30844) <= 16684764;
srom_1(30845) <= 16750311;
srom_1(30846) <= 16776648;
srom_1(30847) <= 16763649;
srom_1(30848) <= 16711377;
srom_1(30849) <= 16620077;
srom_1(30850) <= 16490177;
srom_1(30851) <= 16322286;
srom_1(30852) <= 16117191;
srom_1(30853) <= 15875853;
srom_1(30854) <= 15599406;
srom_1(30855) <= 15289145;
srom_1(30856) <= 14946525;
srom_1(30857) <= 14573152;
srom_1(30858) <= 14170778;
srom_1(30859) <= 13741289;
srom_1(30860) <= 13286700;
srom_1(30861) <= 12809142;
srom_1(30862) <= 12310854;
srom_1(30863) <= 11794174;
srom_1(30864) <= 11261524;
srom_1(30865) <= 10715402;
srom_1(30866) <= 10158369;
srom_1(30867) <= 9593036;
srom_1(30868) <= 9022056;
srom_1(30869) <= 8448105;
srom_1(30870) <= 7873875;
srom_1(30871) <= 7302059;
srom_1(30872) <= 6735338;
srom_1(30873) <= 6176370;
srom_1(30874) <= 5627776;
srom_1(30875) <= 5092128;
srom_1(30876) <= 4571939;
srom_1(30877) <= 4069647;
srom_1(30878) <= 3587608;
srom_1(30879) <= 3128083;
srom_1(30880) <= 2693226;
srom_1(30881) <= 2285077;
srom_1(30882) <= 1905550;
srom_1(30883) <= 1556423;
srom_1(30884) <= 1239336;
srom_1(30885) <= 955773;
srom_1(30886) <= 707066;
srom_1(30887) <= 494380;
srom_1(30888) <= 318713;
srom_1(30889) <= 180888;
srom_1(30890) <= 81552;
srom_1(30891) <= 21171;
srom_1(30892) <= 27;
srom_1(30893) <= 18221;
srom_1(30894) <= 75666;
srom_1(30895) <= 172093;
srom_1(30896) <= 307050;
srom_1(30897) <= 479905;
srom_1(30898) <= 689846;
srom_1(30899) <= 935889;
srom_1(30900) <= 1216881;
srom_1(30901) <= 1531503;
srom_1(30902) <= 1878281;
srom_1(30903) <= 2255588;
srom_1(30904) <= 2661654;
srom_1(30905) <= 3094577;
srom_1(30906) <= 3552324;
srom_1(30907) <= 4032751;
srom_1(30908) <= 4533604;
srom_1(30909) <= 5052534;
srom_1(30910) <= 5587109;
srom_1(30911) <= 6134820;
srom_1(30912) <= 6693100;
srom_1(30913) <= 7259331;
srom_1(30914) <= 7830858;
srom_1(30915) <= 8405000;
srom_1(30916) <= 8979065;
srom_1(30917) <= 9550362;
srom_1(30918) <= 10116210;
srom_1(30919) <= 10673957;
srom_1(30920) <= 11220988;
srom_1(30921) <= 11754736;
srom_1(30922) <= 12272700;
srom_1(30923) <= 12772449;
srom_1(30924) <= 13251641;
srom_1(30925) <= 13708029;
srom_1(30926) <= 14139472;
srom_1(30927) <= 14543948;
srom_1(30928) <= 14919559;
srom_1(30929) <= 15264544;
srom_1(30930) <= 15577285;
srom_1(30931) <= 15856316;
srom_1(30932) <= 16100329;
srom_1(30933) <= 16308179;
srom_1(30934) <= 16478891;
srom_1(30935) <= 16611665;
srom_1(30936) <= 16705878;
srom_1(30937) <= 16761088;
srom_1(30938) <= 16777037;
srom_1(30939) <= 16753650;
srom_1(30940) <= 16691037;
srom_1(30941) <= 16589490;
srom_1(30942) <= 16449487;
srom_1(30943) <= 16271683;
srom_1(30944) <= 16056913;
srom_1(30945) <= 15806184;
srom_1(30946) <= 15520671;
srom_1(30947) <= 15201713;
srom_1(30948) <= 14850807;
srom_1(30949) <= 14469597;
srom_1(30950) <= 14059871;
srom_1(30951) <= 13623550;
srom_1(30952) <= 13162681;
srom_1(30953) <= 12679425;
srom_1(30954) <= 12176048;
srom_1(30955) <= 11654910;
srom_1(30956) <= 11118455;
srom_1(30957) <= 10569199;
srom_1(30958) <= 10009718;
srom_1(30959) <= 9442634;
srom_1(30960) <= 8870608;
srom_1(30961) <= 8296322;
srom_1(30962) <= 7722468;
srom_1(30963) <= 7151738;
srom_1(30964) <= 6586809;
srom_1(30965) <= 6030328;
srom_1(30966) <= 5484906;
srom_1(30967) <= 4953101;
srom_1(30968) <= 4437406;
srom_1(30969) <= 3940239;
srom_1(30970) <= 3463933;
srom_1(30971) <= 3010720;
srom_1(30972) <= 2582725;
srom_1(30973) <= 2181957;
srom_1(30974) <= 1810293;
srom_1(30975) <= 1469478;
srom_1(30976) <= 1161108;
srom_1(30977) <= 886631;
srom_1(30978) <= 647334;
srom_1(30979) <= 444337;
srom_1(30980) <= 278594;
srom_1(30981) <= 150882;
srom_1(30982) <= 61799;
srom_1(30983) <= 11764;
srom_1(30984) <= 1010;
srom_1(30985) <= 29589;
srom_1(30986) <= 97366;
srom_1(30987) <= 204024;
srom_1(30988) <= 349062;
srom_1(30989) <= 531800;
srom_1(30990) <= 751381;
srom_1(30991) <= 1006776;
srom_1(30992) <= 1296787;
srom_1(30993) <= 1620053;
srom_1(30994) <= 1975060;
srom_1(30995) <= 2360143;
srom_1(30996) <= 2773494;
srom_1(30997) <= 3213177;
srom_1(30998) <= 3677129;
srom_1(30999) <= 4163176;
srom_1(31000) <= 4669036;
srom_1(31001) <= 5192339;
srom_1(31002) <= 5730630;
srom_1(31003) <= 6281386;
srom_1(31004) <= 6842022;
srom_1(31005) <= 7409912;
srom_1(31006) <= 7982391;
srom_1(31007) <= 8556774;
srom_1(31008) <= 9130369;
srom_1(31009) <= 9700486;
srom_1(31010) <= 10264451;
srom_1(31011) <= 10819619;
srom_1(31012) <= 11363388;
srom_1(31013) <= 11893207;
srom_1(31014) <= 12406591;
srom_1(31015) <= 12901134;
srom_1(31016) <= 13374516;
srom_1(31017) <= 13824517;
srom_1(31018) <= 14249028;
srom_1(31019) <= 14646057;
srom_1(31020) <= 15013742;
srom_1(31021) <= 15350360;
srom_1(31022) <= 15654332;
srom_1(31023) <= 15924233;
srom_1(31024) <= 16158796;
srom_1(31025) <= 16356923;
srom_1(31026) <= 16517683;
srom_1(31027) <= 16640323;
srom_1(31028) <= 16724268;
srom_1(31029) <= 16769124;
srom_1(31030) <= 16774681;
srom_1(31031) <= 16740913;
srom_1(31032) <= 16667978;
srom_1(31033) <= 16556218;
srom_1(31034) <= 16406158;
srom_1(31035) <= 16218500;
srom_1(31036) <= 15994126;
srom_1(31037) <= 15734086;
srom_1(31038) <= 15439601;
srom_1(31039) <= 15112052;
srom_1(31040) <= 14752974;
srom_1(31041) <= 14364051;
srom_1(31042) <= 13947107;
srom_1(31043) <= 13504098;
srom_1(31044) <= 13037100;
srom_1(31045) <= 12548304;
srom_1(31046) <= 12040002;
srom_1(31047) <= 11514577;
srom_1(31048) <= 10974493;
srom_1(31049) <= 10422283;
srom_1(31050) <= 9860537;
srom_1(31051) <= 9291888;
srom_1(31052) <= 8719003;
srom_1(31053) <= 8144569;
srom_1(31054) <= 7571279;
srom_1(31055) <= 7001823;
srom_1(31056) <= 6438869;
srom_1(31057) <= 5885058;
srom_1(31058) <= 5342987;
srom_1(31059) <= 4815198;
srom_1(31060) <= 4304167;
srom_1(31061) <= 3812288;
srom_1(31062) <= 3341869;
srom_1(31063) <= 2895117;
srom_1(31064) <= 2474125;
srom_1(31065) <= 2080868;
srom_1(31066) <= 1717190;
srom_1(31067) <= 1384797;
srom_1(31068) <= 1085247;
srom_1(31069) <= 819946;
srom_1(31070) <= 590136;
srom_1(31071) <= 396896;
srom_1(31072) <= 241131;
srom_1(31073) <= 123573;
srom_1(31074) <= 44773;
srom_1(31075) <= 5100;
srom_1(31076) <= 4740;
srom_1(31077) <= 43694;
srom_1(31078) <= 121781;
srom_1(31079) <= 238634;
srom_1(31080) <= 393705;
srom_1(31081) <= 586267;
srom_1(31082) <= 815416;
srom_1(31083) <= 1080079;
srom_1(31084) <= 1379014;
srom_1(31085) <= 1710820;
srom_1(31086) <= 2073940;
srom_1(31087) <= 2466671;
srom_1(31088) <= 2887173;
srom_1(31089) <= 3333472;
srom_1(31090) <= 3803477;
srom_1(31091) <= 4294983;
srom_1(31092) <= 4805686;
srom_1(31093) <= 5333190;
srom_1(31094) <= 5875022;
srom_1(31095) <= 6428641;
srom_1(31096) <= 6991451;
srom_1(31097) <= 7560813;
srom_1(31098) <= 8134056;
srom_1(31099) <= 8708493;
srom_1(31100) <= 9281431;
srom_1(31101) <= 9850181;
srom_1(31102) <= 10412078;
srom_1(31103) <= 10964485;
srom_1(31104) <= 11504814;
srom_1(31105) <= 12030530;
srom_1(31106) <= 12539167;
srom_1(31107) <= 13028341;
srom_1(31108) <= 13495758;
srom_1(31109) <= 13939226;
srom_1(31110) <= 14356664;
srom_1(31111) <= 14746117;
srom_1(31112) <= 15105757;
srom_1(31113) <= 15433898;
srom_1(31114) <= 15729001;
srom_1(31115) <= 15989682;
srom_1(31116) <= 16214720;
srom_1(31117) <= 16403058;
srom_1(31118) <= 16553814;
srom_1(31119) <= 16666280;
srom_1(31120) <= 16739929;
srom_1(31121) <= 16774416;
srom_1(31122) <= 16769579;
srom_1(31123) <= 16725441;
srom_1(31124) <= 16642209;
srom_1(31125) <= 16520272;
srom_1(31126) <= 16360204;
srom_1(31127) <= 16162754;
srom_1(31128) <= 15928848;
srom_1(31129) <= 15659583;
srom_1(31130) <= 15356223;
srom_1(31131) <= 15020188;
srom_1(31132) <= 14653056;
srom_1(31133) <= 14256548;
srom_1(31134) <= 13832523;
srom_1(31135) <= 13382970;
srom_1(31136) <= 12909996;
srom_1(31137) <= 12415821;
srom_1(31138) <= 11902760;
srom_1(31139) <= 11373220;
srom_1(31140) <= 10829684;
srom_1(31141) <= 10274701;
srom_1(31142) <= 9710873;
srom_1(31143) <= 9140845;
srom_1(31144) <= 8567290;
srom_1(31145) <= 7992896;
srom_1(31146) <= 7420358;
srom_1(31147) <= 6852361;
srom_1(31148) <= 6291567;
srom_1(31149) <= 5740608;
srom_1(31150) <= 5202065;
srom_1(31151) <= 4678466;
srom_1(31152) <= 4172265;
srom_1(31153) <= 3685835;
srom_1(31154) <= 3221458;
srom_1(31155) <= 2781312;
srom_1(31156) <= 2367461;
srom_1(31157) <= 1981845;
srom_1(31158) <= 1626272;
srom_1(31159) <= 1302410;
srom_1(31160) <= 1011777;
srom_1(31161) <= 755738;
srom_1(31162) <= 535491;
srom_1(31163) <= 352070;
srom_1(31164) <= 206336;
srom_1(31165) <= 98971;
srom_1(31166) <= 30478;
srom_1(31167) <= 1180;
srom_1(31168) <= 11214;
srom_1(31169) <= 60532;
srom_1(31170) <= 148903;
srom_1(31171) <= 275913;
srom_1(31172) <= 440966;
srom_1(31173) <= 643288;
srom_1(31174) <= 881931;
srom_1(31175) <= 1155775;
srom_1(31176) <= 1463537;
srom_1(31177) <= 1803772;
srom_1(31178) <= 2174886;
srom_1(31179) <= 2575138;
srom_1(31180) <= 3002652;
srom_1(31181) <= 3455422;
srom_1(31182) <= 3931326;
srom_1(31183) <= 4428131;
srom_1(31184) <= 4943509;
srom_1(31185) <= 5475041;
srom_1(31186) <= 6020237;
srom_1(31187) <= 6576538;
srom_1(31188) <= 7141337;
srom_1(31189) <= 7711985;
srom_1(31190) <= 8285805;
srom_1(31191) <= 8860108;
srom_1(31192) <= 9432200;
srom_1(31193) <= 9999397;
srom_1(31194) <= 10559042;
srom_1(31195) <= 11108508;
srom_1(31196) <= 11645220;
srom_1(31197) <= 12166661;
srom_1(31198) <= 12670384;
srom_1(31199) <= 13154030;
srom_1(31200) <= 13615328;
srom_1(31201) <= 14052117;
srom_1(31202) <= 14462347;
srom_1(31203) <= 14844096;
srom_1(31204) <= 15195572;
srom_1(31205) <= 15515129;
srom_1(31206) <= 15801266;
srom_1(31207) <= 16052643;
srom_1(31208) <= 16268081;
srom_1(31209) <= 16446570;
srom_1(31210) <= 16587271;
srom_1(31211) <= 16689527;
srom_1(31212) <= 16752856;
srom_1(31213) <= 16776963;
srom_1(31214) <= 16761734;
srom_1(31215) <= 16707240;
srom_1(31216) <= 16613737;
srom_1(31217) <= 16481664;
srom_1(31218) <= 16311640;
srom_1(31219) <= 16104462;
srom_1(31220) <= 15861102;
srom_1(31221) <= 15582700;
srom_1(31222) <= 15270563;
srom_1(31223) <= 14926154;
srom_1(31224) <= 14551089;
srom_1(31225) <= 14147125;
srom_1(31226) <= 13716158;
srom_1(31227) <= 13260207;
srom_1(31228) <= 12781413;
srom_1(31229) <= 12282019;
srom_1(31230) <= 11764367;
srom_1(31231) <= 11230885;
srom_1(31232) <= 10684075;
srom_1(31233) <= 10126501;
srom_1(31234) <= 9560777;
srom_1(31235) <= 8989556;
srom_1(31236) <= 8415518;
srom_1(31237) <= 7841353;
srom_1(31238) <= 7269754;
srom_1(31239) <= 6703402;
srom_1(31240) <= 6144953;
srom_1(31241) <= 5597024;
srom_1(31242) <= 5062187;
srom_1(31243) <= 4542948;
srom_1(31244) <= 4041743;
srom_1(31245) <= 3560922;
srom_1(31246) <= 3102739;
srom_1(31247) <= 2669344;
srom_1(31248) <= 2262768;
srom_1(31249) <= 1884918;
srom_1(31250) <= 1537567;
srom_1(31251) <= 1222342;
srom_1(31252) <= 940723;
srom_1(31253) <= 694029;
srom_1(31254) <= 483417;
srom_1(31255) <= 309876;
srom_1(31256) <= 174219;
srom_1(31257) <= 77082;
srom_1(31258) <= 18920;
srom_1(31259) <= 7;
srom_1(31260) <= 20431;
srom_1(31261) <= 80096;
srom_1(31262) <= 178722;
srom_1(31263) <= 315847;
srom_1(31264) <= 490829;
srom_1(31265) <= 702846;
srom_1(31266) <= 950903;
srom_1(31267) <= 1233839;
srom_1(31268) <= 1550326;
srom_1(31269) <= 1898880;
srom_1(31270) <= 2277867;
srom_1(31271) <= 2685509;
srom_1(31272) <= 3119895;
srom_1(31273) <= 3578987;
srom_1(31274) <= 4060634;
srom_1(31275) <= 4562576;
srom_1(31276) <= 5082459;
srom_1(31277) <= 5617846;
srom_1(31278) <= 6166227;
srom_1(31279) <= 6725028;
srom_1(31280) <= 7291631;
srom_1(31281) <= 7863378;
srom_1(31282) <= 8437588;
srom_1(31283) <= 9011568;
srom_1(31284) <= 9582627;
srom_1(31285) <= 10148086;
srom_1(31286) <= 10705295;
srom_1(31287) <= 11251640;
srom_1(31288) <= 11784560;
srom_1(31289) <= 12301554;
srom_1(31290) <= 12800200;
srom_1(31291) <= 13278158;
srom_1(31292) <= 13733187;
srom_1(31293) <= 14163154;
srom_1(31294) <= 14566041;
srom_1(31295) <= 14939961;
srom_1(31296) <= 15283159;
srom_1(31297) <= 15594026;
srom_1(31298) <= 15871105;
srom_1(31299) <= 16113095;
srom_1(31300) <= 16318863;
srom_1(31301) <= 16487443;
srom_1(31302) <= 16618045;
srom_1(31303) <= 16710056;
srom_1(31304) <= 16763045;
srom_1(31305) <= 16776763;
srom_1(31306) <= 16751147;
srom_1(31307) <= 16686315;
srom_1(31308) <= 16582573;
srom_1(31309) <= 16440406;
srom_1(31310) <= 16260482;
srom_1(31311) <= 16043644;
srom_1(31312) <= 15790909;
srom_1(31313) <= 15503462;
srom_1(31314) <= 15182650;
srom_1(31315) <= 14829980;
srom_1(31316) <= 14447103;
srom_1(31317) <= 14035816;
srom_1(31318) <= 13598047;
srom_1(31319) <= 13135850;
srom_1(31320) <= 12651391;
srom_1(31321) <= 12146942;
srom_1(31322) <= 11624870;
srom_1(31323) <= 11087621;
srom_1(31324) <= 10537715;
srom_1(31325) <= 9977732;
srom_1(31326) <= 9410297;
srom_1(31327) <= 8838071;
srom_1(31328) <= 8263737;
srom_1(31329) <= 7689988;
srom_1(31330) <= 7119516;
srom_1(31331) <= 6554995;
srom_1(31332) <= 5999072;
srom_1(31333) <= 5454355;
srom_1(31334) <= 4923397;
srom_1(31335) <= 4408689;
srom_1(31336) <= 3912644;
srom_1(31337) <= 3437589;
srom_1(31338) <= 2985750;
srom_1(31339) <= 2559248;
srom_1(31340) <= 2160081;
srom_1(31341) <= 1790122;
srom_1(31342) <= 1451105;
srom_1(31343) <= 1144621;
srom_1(31344) <= 872106;
srom_1(31345) <= 634839;
srom_1(31346) <= 433932;
srom_1(31347) <= 270327;
srom_1(31348) <= 144791;
srom_1(31349) <= 57914;
srom_1(31350) <= 10102;
srom_1(31351) <= 1580;
srom_1(31352) <= 32387;
srom_1(31353) <= 102379;
srom_1(31354) <= 211229;
srom_1(31355) <= 358425;
srom_1(31356) <= 543277;
srom_1(31357) <= 764919;
srom_1(31358) <= 1022311;
srom_1(31359) <= 1314246;
srom_1(31360) <= 1639355;
srom_1(31361) <= 1996113;
srom_1(31362) <= 2382849;
srom_1(31363) <= 2797747;
srom_1(31364) <= 3238863;
srom_1(31365) <= 3704127;
srom_1(31366) <= 4191359;
srom_1(31367) <= 4698273;
srom_1(31368) <= 5222492;
srom_1(31369) <= 5761559;
srom_1(31370) <= 6312944;
srom_1(31371) <= 6874063;
srom_1(31372) <= 7442284;
srom_1(31373) <= 8014943;
srom_1(31374) <= 8589354;
srom_1(31375) <= 9162824;
srom_1(31376) <= 9732663;
srom_1(31377) <= 10296199;
srom_1(31378) <= 10850790;
srom_1(31379) <= 11393835;
srom_1(31380) <= 11922788;
srom_1(31381) <= 12435167;
srom_1(31382) <= 12928571;
srom_1(31383) <= 13400685;
srom_1(31384) <= 13849296;
srom_1(31385) <= 14272300;
srom_1(31386) <= 14667713;
srom_1(31387) <= 15033681;
srom_1(31388) <= 15368489;
srom_1(31389) <= 15670565;
srom_1(31390) <= 15938493;
srom_1(31391) <= 16171018;
srom_1(31392) <= 16367048;
srom_1(31393) <= 16525665;
srom_1(31394) <= 16646124;
srom_1(31395) <= 16727861;
srom_1(31396) <= 16770492;
srom_1(31397) <= 16773817;
srom_1(31398) <= 16737822;
srom_1(31399) <= 16662674;
srom_1(31400) <= 16548726;
srom_1(31401) <= 16396512;
srom_1(31402) <= 16206747;
srom_1(31403) <= 15980320;
srom_1(31404) <= 15718293;
srom_1(31405) <= 15421894;
srom_1(31406) <= 15092513;
srom_1(31407) <= 14731696;
srom_1(31408) <= 14341134;
srom_1(31409) <= 13922658;
srom_1(31410) <= 13478232;
srom_1(31411) <= 13009938;
srom_1(31412) <= 12519973;
srom_1(31413) <= 12010635;
srom_1(31414) <= 11484312;
srom_1(31415) <= 10943473;
srom_1(31416) <= 10390652;
srom_1(31417) <= 9828443;
srom_1(31418) <= 9259483;
srom_1(31419) <= 8686438;
srom_1(31420) <= 8111997;
srom_1(31421) <= 7538853;
srom_1(31422) <= 6969694;
srom_1(31423) <= 6407188;
srom_1(31424) <= 5853974;
srom_1(31425) <= 5312646;
srom_1(31426) <= 4785742;
srom_1(31427) <= 4275733;
srom_1(31428) <= 3785011;
srom_1(31429) <= 3315877;
srom_1(31430) <= 2870530;
srom_1(31431) <= 2451060;
srom_1(31432) <= 2059433;
srom_1(31433) <= 1697485;
srom_1(31434) <= 1366915;
srom_1(31435) <= 1069271;
srom_1(31436) <= 805951;
srom_1(31437) <= 578188;
srom_1(31438) <= 387051;
srom_1(31439) <= 233436;
srom_1(31440) <= 118063;
srom_1(31441) <= 41474;
srom_1(31442) <= 4027;
srom_1(31443) <= 5898;
srom_1(31444) <= 47079;
srom_1(31445) <= 127376;
srom_1(31446) <= 246413;
srom_1(31447) <= 403632;
srom_1(31448) <= 598294;
srom_1(31449) <= 829489;
srom_1(31450) <= 1096130;
srom_1(31451) <= 1396968;
srom_1(31452) <= 1730593;
srom_1(31453) <= 2095439;
srom_1(31454) <= 2489796;
srom_1(31455) <= 2911815;
srom_1(31456) <= 3359516;
srom_1(31457) <= 3830801;
srom_1(31458) <= 4323458;
srom_1(31459) <= 4835179;
srom_1(31460) <= 5363562;
srom_1(31461) <= 5906131;
srom_1(31462) <= 6460342;
srom_1(31463) <= 7023594;
srom_1(31464) <= 7593248;
srom_1(31465) <= 8166631;
srom_1(31466) <= 8741055;
srom_1(31467) <= 9313827;
srom_1(31468) <= 9882259;
srom_1(31469) <= 10443688;
srom_1(31470) <= 10995479;
srom_1(31471) <= 11535046;
srom_1(31472) <= 12059859;
srom_1(31473) <= 12567455;
srom_1(31474) <= 13055456;
srom_1(31475) <= 13521572;
srom_1(31476) <= 13963617;
srom_1(31477) <= 14379520;
srom_1(31478) <= 14767329;
srom_1(31479) <= 15125226;
srom_1(31480) <= 15451533;
srom_1(31481) <= 15744719;
srom_1(31482) <= 16003410;
srom_1(31483) <= 16226393;
srom_1(31484) <= 16412622;
srom_1(31485) <= 16561223;
srom_1(31486) <= 16671500;
srom_1(31487) <= 16742935;
srom_1(31488) <= 16775194;
srom_1(31489) <= 16768126;
srom_1(31490) <= 16721763;
srom_1(31491) <= 16636323;
srom_1(31492) <= 16512207;
srom_1(31493) <= 16349997;
srom_1(31494) <= 16150453;
srom_1(31495) <= 15914510;
srom_1(31496) <= 15643277;
srom_1(31497) <= 15338023;
srom_1(31498) <= 15000182;
srom_1(31499) <= 14631336;
srom_1(31500) <= 14233216;
srom_1(31501) <= 13807689;
srom_1(31502) <= 13356750;
srom_1(31503) <= 12882513;
srom_1(31504) <= 12387203;
srom_1(31505) <= 11873143;
srom_1(31506) <= 11342742;
srom_1(31507) <= 10798488;
srom_1(31508) <= 10242933;
srom_1(31509) <= 9678683;
srom_1(31510) <= 9108383;
srom_1(31511) <= 8534708;
srom_1(31512) <= 7960348;
srom_1(31513) <= 7387996;
srom_1(31514) <= 6820336;
srom_1(31515) <= 6260030;
srom_1(31516) <= 5709706;
srom_1(31517) <= 5171945;
srom_1(31518) <= 4649267;
srom_1(31519) <= 4144124;
srom_1(31520) <= 3658885;
srom_1(31521) <= 3195826;
srom_1(31522) <= 2757117;
srom_1(31523) <= 2344816;
srom_1(31524) <= 1960857;
srom_1(31525) <= 1607039;
srom_1(31526) <= 1285023;
srom_1(31527) <= 996318;
srom_1(31528) <= 742278;
srom_1(31529) <= 524094;
srom_1(31530) <= 342789;
srom_1(31531) <= 199214;
srom_1(31532) <= 94042;
srom_1(31533) <= 27766;
srom_1(31534) <= 697;
srom_1(31535) <= 12961;
srom_1(31536) <= 64502;
srom_1(31537) <= 155078;
srom_1(31538) <= 284263;
srom_1(31539) <= 451452;
srom_1(31540) <= 655862;
srom_1(31541) <= 896533;
srom_1(31542) <= 1172337;
srom_1(31543) <= 1481980;
srom_1(31544) <= 1824011;
srom_1(31545) <= 2196825;
srom_1(31546) <= 2598675;
srom_1(31547) <= 3027676;
srom_1(31548) <= 3481817;
srom_1(31549) <= 3958966;
srom_1(31550) <= 4456888;
srom_1(31551) <= 4973247;
srom_1(31552) <= 5505622;
srom_1(31553) <= 6051516;
srom_1(31554) <= 6608370;
srom_1(31555) <= 7173572;
srom_1(31556) <= 7744471;
srom_1(31557) <= 8318391;
srom_1(31558) <= 8892641;
srom_1(31559) <= 9464526;
srom_1(31560) <= 10031367;
srom_1(31561) <= 10590503;
srom_1(31562) <= 11139315;
srom_1(31563) <= 11675227;
srom_1(31564) <= 12195728;
srom_1(31565) <= 12698375;
srom_1(31566) <= 13180812;
srom_1(31567) <= 13640778;
srom_1(31568) <= 14076114;
srom_1(31569) <= 14484779;
srom_1(31570) <= 14864857;
srom_1(31571) <= 15214566;
srom_1(31572) <= 15532265;
srom_1(31573) <= 15816466;
srom_1(31574) <= 16065834;
srom_1(31575) <= 16279202;
srom_1(31576) <= 16455568;
srom_1(31577) <= 16594105;
srom_1(31578) <= 16694164;
srom_1(31579) <= 16755275;
srom_1(31580) <= 16777151;
srom_1(31581) <= 16759692;
srom_1(31582) <= 16702977;
srom_1(31583) <= 16607273;
srom_1(31584) <= 16473029;
srom_1(31585) <= 16300875;
srom_1(31586) <= 16091617;
srom_1(31587) <= 15846237;
srom_1(31588) <= 15565886;
srom_1(31589) <= 15251877;
srom_1(31590) <= 14905685;
srom_1(31591) <= 14528932;
srom_1(31592) <= 14123385;
srom_1(31593) <= 13690945;
srom_1(31594) <= 13233641;
srom_1(31595) <= 12753617;
srom_1(31596) <= 12253124;
srom_1(31597) <= 11734509;
srom_1(31598) <= 11200204;
srom_1(31599) <= 10652714;
srom_1(31600) <= 10094607;
srom_1(31601) <= 9528500;
srom_1(31602) <= 8957048;
srom_1(31603) <= 8382930;
srom_1(31604) <= 7808839;
srom_1(31605) <= 7237466;
srom_1(31606) <= 6671491;
srom_1(31607) <= 6113569;
srom_1(31608) <= 5566315;
srom_1(31609) <= 5032296;
srom_1(31610) <= 4514016;
srom_1(31611) <= 4013904;
srom_1(31612) <= 3534308;
srom_1(31613) <= 3077475;
srom_1(31614) <= 2645547;
srom_1(31615) <= 2240551;
srom_1(31616) <= 1864385;
srom_1(31617) <= 1518814;
srom_1(31618) <= 1205457;
srom_1(31619) <= 925785;
srom_1(31620) <= 681108;
srom_1(31621) <= 472574;
srom_1(31622) <= 301162;
srom_1(31623) <= 167674;
srom_1(31624) <= 72737;
srom_1(31625) <= 16796;
srom_1(31626) <= 113;
srom_1(31627) <= 22767;
srom_1(31628) <= 84651;
srom_1(31629) <= 185475;
srom_1(31630) <= 324766;
srom_1(31631) <= 501872;
srom_1(31632) <= 715961;
srom_1(31633) <= 966030;
srom_1(31634) <= 1250906;
srom_1(31635) <= 1569253;
srom_1(31636) <= 1919578;
srom_1(31637) <= 2300239;
srom_1(31638) <= 2709450;
srom_1(31639) <= 3145293;
srom_1(31640) <= 3605723;
srom_1(31641) <= 4088582;
srom_1(31642) <= 4591606;
srom_1(31643) <= 5112434;
srom_1(31644) <= 5648626;
srom_1(31645) <= 6197667;
srom_1(31646) <= 6756981;
srom_1(31647) <= 7323947;
srom_1(31648) <= 7895906;
srom_1(31649) <= 8470175;
srom_1(31650) <= 9044061;
srom_1(31651) <= 9614874;
srom_1(31652) <= 10179936;
srom_1(31653) <= 10736598;
srom_1(31654) <= 11282250;
srom_1(31655) <= 11814332;
srom_1(31656) <= 12330350;
srom_1(31657) <= 12827884;
srom_1(31658) <= 13304600;
srom_1(31659) <= 13758264;
srom_1(31660) <= 14186748;
srom_1(31661) <= 14588042;
srom_1(31662) <= 14960264;
srom_1(31663) <= 15301670;
srom_1(31664) <= 15610659;
srom_1(31665) <= 15885780;
srom_1(31666) <= 16125745;
srom_1(31667) <= 16329428;
srom_1(31668) <= 16495873;
srom_1(31669) <= 16624301;
srom_1(31670) <= 16714108;
srom_1(31671) <= 16764875;
srom_1(31672) <= 16776362;
srom_1(31673) <= 16748516;
srom_1(31674) <= 16681468;
srom_1(31675) <= 16575532;
srom_1(31676) <= 16431204;
srom_1(31677) <= 16249162;
srom_1(31678) <= 16030259;
srom_1(31679) <= 15775522;
srom_1(31680) <= 15486145;
srom_1(31681) <= 15163485;
srom_1(31682) <= 14809055;
srom_1(31683) <= 14424518;
srom_1(31684) <= 14011676;
srom_1(31685) <= 13572466;
srom_1(31686) <= 13108947;
srom_1(31687) <= 12623292;
srom_1(31688) <= 12117780;
srom_1(31689) <= 11594780;
srom_1(31690) <= 11056746;
srom_1(31691) <= 10506199;
srom_1(31692) <= 9945723;
srom_1(31693) <= 9377944;
srom_1(31694) <= 8805526;
srom_1(31695) <= 8231154;
srom_1(31696) <= 7657519;
srom_1(31697) <= 7087313;
srom_1(31698) <= 6523209;
srom_1(31699) <= 5967853;
srom_1(31700) <= 5423848;
srom_1(31701) <= 4893746;
srom_1(31702) <= 4380033;
srom_1(31703) <= 3885117;
srom_1(31704) <= 3411320;
srom_1(31705) <= 2960863;
srom_1(31706) <= 2535858;
srom_1(31707) <= 2138299;
srom_1(31708) <= 1770050;
srom_1(31709) <= 1432837;
srom_1(31710) <= 1128243;
srom_1(31711) <= 857695;
srom_1(31712) <= 622462;
srom_1(31713) <= 423647;
srom_1(31714) <= 262182;
srom_1(31715) <= 138825;
srom_1(31716) <= 54154;
srom_1(31717) <= 8566;
srom_1(31718) <= 2275;
srom_1(31719) <= 35311;
srom_1(31720) <= 107518;
srom_1(31721) <= 218558;
srom_1(31722) <= 367910;
srom_1(31723) <= 554873;
srom_1(31724) <= 778572;
srom_1(31725) <= 1037957;
srom_1(31726) <= 1331812;
srom_1(31727) <= 1658758;
srom_1(31728) <= 2017263;
srom_1(31729) <= 2405645;
srom_1(31730) <= 2822084;
srom_1(31731) <= 3264626;
srom_1(31732) <= 3731196;
srom_1(31733) <= 4219606;
srom_1(31734) <= 4727566;
srom_1(31735) <= 5252694;
srom_1(31736) <= 5792527;
srom_1(31737) <= 6344534;
srom_1(31738) <= 6906127;
srom_1(31739) <= 7474671;
srom_1(31740) <= 8047501;
srom_1(31741) <= 8621931;
srom_1(31742) <= 9195267;
srom_1(31743) <= 9764820;
srom_1(31744) <= 10327919;
srom_1(31745) <= 10881924;
srom_1(31746) <= 11424237;
srom_1(31747) <= 11952316;
srom_1(31748) <= 12463682;
srom_1(31749) <= 12955939;
srom_1(31750) <= 13426779;
srom_1(31751) <= 13873992;
srom_1(31752) <= 14295483;
srom_1(31753) <= 14689275;
srom_1(31754) <= 15053520;
srom_1(31755) <= 15386512;
srom_1(31756) <= 15686687;
srom_1(31757) <= 15952640;
srom_1(31758) <= 16183122;
srom_1(31759) <= 16377053;
srom_1(31760) <= 16533524;
srom_1(31761) <= 16651800;
srom_1(31762) <= 16731327;
srom_1(31763) <= 16771733;
srom_1(31764) <= 16772827;
srom_1(31765) <= 16734604;
srom_1(31766) <= 16657244;
srom_1(31767) <= 16541110;
srom_1(31768) <= 16386746;
srom_1(31769) <= 16194876;
srom_1(31770) <= 15966400;
srom_1(31771) <= 15702388;
srom_1(31772) <= 15404080;
srom_1(31773) <= 15072874;
srom_1(31774) <= 14710323;
srom_1(31775) <= 14318128;
srom_1(31776) <= 13898126;
srom_1(31777) <= 13452289;
srom_1(31778) <= 12982707;
srom_1(31779) <= 12491581;
srom_1(31780) <= 11981215;
srom_1(31781) <= 11454001;
srom_1(31782) <= 10912414;
srom_1(31783) <= 10358991;
srom_1(31784) <= 9796328;
srom_1(31785) <= 9227064;
srom_1(31786) <= 8653869;
srom_1(31787) <= 8079429;
srom_1(31788) <= 7506439;
srom_1(31789) <= 6937586;
srom_1(31790) <= 6375538;
srom_1(31791) <= 5822929;
srom_1(31792) <= 5282352;
srom_1(31793) <= 4756341;
srom_1(31794) <= 4247362;
srom_1(31795) <= 3757804;
srom_1(31796) <= 3289961;
srom_1(31797) <= 2846027;
srom_1(31798) <= 2428085;
srom_1(31799) <= 2038093;
srom_1(31800) <= 1677881;
srom_1(31801) <= 1349138;
srom_1(31802) <= 1053406;
srom_1(31803) <= 792070;
srom_1(31804) <= 566358;
srom_1(31805) <= 377326;
srom_1(31806) <= 225863;
srom_1(31807) <= 112677;
srom_1(31808) <= 38300;
srom_1(31809) <= 3080;
srom_1(31810) <= 7183;
srom_1(31811) <= 50590;
srom_1(31812) <= 133096;
srom_1(31813) <= 254315;
srom_1(31814) <= 413679;
srom_1(31815) <= 610440;
srom_1(31816) <= 843675;
srom_1(31817) <= 1112291;
srom_1(31818) <= 1415028;
srom_1(31819) <= 1750467;
srom_1(31820) <= 2117034;
srom_1(31821) <= 2513011;
srom_1(31822) <= 2936540;
srom_1(31823) <= 3385636;
srom_1(31824) <= 3858193;
srom_1(31825) <= 4351995;
srom_1(31826) <= 4864725;
srom_1(31827) <= 5393980;
srom_1(31828) <= 5937278;
srom_1(31829) <= 6492071;
srom_1(31830) <= 7055758;
srom_1(31831) <= 7625695;
srom_1(31832) <= 8199209;
srom_1(31833) <= 8773611;
srom_1(31834) <= 9346209;
srom_1(31835) <= 9914315;
srom_1(31836) <= 10475267;
srom_1(31837) <= 11026434;
srom_1(31838) <= 11565231;
srom_1(31839) <= 12089132;
srom_1(31840) <= 12595680;
srom_1(31841) <= 13082500;
srom_1(31842) <= 13547308;
srom_1(31843) <= 13987925;
srom_1(31844) <= 14402285;
srom_1(31845) <= 14788445;
srom_1(31846) <= 15144594;
srom_1(31847) <= 15469062;
srom_1(31848) <= 15760327;
srom_1(31849) <= 16017024;
srom_1(31850) <= 16237948;
srom_1(31851) <= 16422064;
srom_1(31852) <= 16568508;
srom_1(31853) <= 16676594;
srom_1(31854) <= 16745815;
srom_1(31855) <= 16775846;
srom_1(31856) <= 16766546;
srom_1(31857) <= 16717960;
srom_1(31858) <= 16630314;
srom_1(31859) <= 16504020;
srom_1(31860) <= 16339670;
srom_1(31861) <= 16138034;
srom_1(31862) <= 15900059;
srom_1(31863) <= 15626860;
srom_1(31864) <= 15319719;
srom_1(31865) <= 14980075;
srom_1(31866) <= 14609521;
srom_1(31867) <= 14209796;
srom_1(31868) <= 13782773;
srom_1(31869) <= 13330455;
srom_1(31870) <= 12854962;
srom_1(31871) <= 12358526;
srom_1(31872) <= 11843473;
srom_1(31873) <= 11312219;
srom_1(31874) <= 10767256;
srom_1(31875) <= 10211138;
srom_1(31876) <= 9646473;
srom_1(31877) <= 9075910;
srom_1(31878) <= 8502124;
srom_1(31879) <= 7927806;
srom_1(31880) <= 7355648;
srom_1(31881) <= 6788334;
srom_1(31882) <= 6228525;
srom_1(31883) <= 5678845;
srom_1(31884) <= 5141872;
srom_1(31885) <= 4620124;
srom_1(31886) <= 4116048;
srom_1(31887) <= 3632007;
srom_1(31888) <= 3170272;
srom_1(31889) <= 2733007;
srom_1(31890) <= 2322263;
srom_1(31891) <= 1939966;
srom_1(31892) <= 1587910;
srom_1(31893) <= 1267744;
srom_1(31894) <= 980970;
srom_1(31895) <= 728933;
srom_1(31896) <= 512815;
srom_1(31897) <= 333629;
srom_1(31898) <= 192216;
srom_1(31899) <= 89239;
srom_1(31900) <= 25180;
srom_1(31901) <= 340;
srom_1(31902) <= 14836;
srom_1(31903) <= 68599;
srom_1(31904) <= 161377;
srom_1(31905) <= 292736;
srom_1(31906) <= 462059;
srom_1(31907) <= 668552;
srom_1(31908) <= 911248;
srom_1(31909) <= 1189007;
srom_1(31910) <= 1500528;
srom_1(31911) <= 1844349;
srom_1(31912) <= 2218858;
srom_1(31913) <= 2622300;
srom_1(31914) <= 3052782;
srom_1(31915) <= 3508285;
srom_1(31916) <= 3986674;
srom_1(31917) <= 4485705;
srom_1(31918) <= 5003038;
srom_1(31919) <= 5536247;
srom_1(31920) <= 6082832;
srom_1(31921) <= 6640229;
srom_1(31922) <= 7205825;
srom_1(31923) <= 7776968;
srom_1(31924) <= 8350978;
srom_1(31925) <= 8925166;
srom_1(31926) <= 9496837;
srom_1(31927) <= 10063311;
srom_1(31928) <= 10621932;
srom_1(31929) <= 11170080;
srom_1(31930) <= 11705185;
srom_1(31931) <= 12224737;
srom_1(31932) <= 12726301;
srom_1(31933) <= 13207523;
srom_1(31934) <= 13666148;
srom_1(31935) <= 14100024;
srom_1(31936) <= 14507118;
srom_1(31937) <= 14885520;
srom_1(31938) <= 15233456;
srom_1(31939) <= 15549294;
srom_1(31940) <= 15831553;
srom_1(31941) <= 16078910;
srom_1(31942) <= 16290204;
srom_1(31943) <= 16464444;
srom_1(31944) <= 16600815;
srom_1(31945) <= 16698675;
srom_1(31946) <= 16757567;
srom_1(31947) <= 16777213;
srom_1(31948) <= 16757523;
srom_1(31949) <= 16698588;
srom_1(31950) <= 16600685;
srom_1(31951) <= 16464272;
srom_1(31952) <= 16289990;
srom_1(31953) <= 16078655;
srom_1(31954) <= 15831260;
srom_1(31955) <= 15548963;
srom_1(31956) <= 15233088;
srom_1(31957) <= 14885118;
srom_1(31958) <= 14506683;
srom_1(31959) <= 14099558;
srom_1(31960) <= 13665653;
srom_1(31961) <= 13207002;
srom_1(31962) <= 12725756;
srom_1(31963) <= 12224171;
srom_1(31964) <= 11704601;
srom_1(31965) <= 11169480;
srom_1(31966) <= 10621319;
srom_1(31967) <= 10062688;
srom_1(31968) <= 9496206;
srom_1(31969) <= 8924531;
srom_1(31970) <= 8350342;
srom_1(31971) <= 7776333;
srom_1(31972) <= 7205195;
srom_1(31973) <= 6639607;
srom_1(31974) <= 6082220;
srom_1(31975) <= 5535648;
srom_1(31976) <= 5002456;
srom_1(31977) <= 4485141;
srom_1(31978) <= 3986132;
srom_1(31979) <= 3507767;
srom_1(31980) <= 3052291;
srom_1(31981) <= 2621838;
srom_1(31982) <= 2218427;
srom_1(31983) <= 1843951;
srom_1(31984) <= 1500164;
srom_1(31985) <= 1188680;
srom_1(31986) <= 910959;
srom_1(31987) <= 668303;
srom_1(31988) <= 461851;
srom_1(31989) <= 292569;
srom_1(31990) <= 161253;
srom_1(31991) <= 68517;
srom_1(31992) <= 14798;
srom_1(31993) <= 346;
srom_1(31994) <= 25229;
srom_1(31995) <= 89331;
srom_1(31996) <= 192352;
srom_1(31997) <= 333807;
srom_1(31998) <= 513034;
srom_1(31999) <= 729192;
srom_1(32000) <= 981268;
srom_1(32001) <= 1268080;
srom_1(32002) <= 1588282;
srom_1(32003) <= 1940373;
srom_1(32004) <= 2322702;
srom_1(32005) <= 2733477;
srom_1(32006) <= 3170770;
srom_1(32007) <= 3632531;
srom_1(32008) <= 4116595;
srom_1(32009) <= 4620693;
srom_1(32010) <= 5142459;
srom_1(32011) <= 5679447;
srom_1(32012) <= 6229140;
srom_1(32013) <= 6788959;
srom_1(32014) <= 7356280;
srom_1(32015) <= 7928441;
srom_1(32016) <= 8502760;
srom_1(32017) <= 9076544;
srom_1(32018) <= 9647102;
srom_1(32019) <= 10211759;
srom_1(32020) <= 10767866;
srom_1(32021) <= 11312816;
srom_1(32022) <= 11844053;
srom_1(32023) <= 12359086;
srom_1(32024) <= 12855501;
srom_1(32025) <= 13330969;
srom_1(32026) <= 13783260;
srom_1(32027) <= 14210254;
srom_1(32028) <= 14609948;
srom_1(32029) <= 14980469;
srom_1(32030) <= 15320077;
srom_1(32031) <= 15627182;
srom_1(32032) <= 15900342;
srom_1(32033) <= 16138278;
srom_1(32034) <= 16339872;
srom_1(32035) <= 16504181;
srom_1(32036) <= 16630432;
srom_1(32037) <= 16718035;
srom_1(32038) <= 16766578;
srom_1(32039) <= 16775835;
srom_1(32040) <= 16745760;
srom_1(32041) <= 16676496;
srom_1(32042) <= 16568367;
srom_1(32043) <= 16421881;
srom_1(32044) <= 16237723;
srom_1(32045) <= 16016759;
srom_1(32046) <= 15760023;
srom_1(32047) <= 15468721;
srom_1(32048) <= 15144217;
srom_1(32049) <= 14788034;
srom_1(32050) <= 14401842;
srom_1(32051) <= 13987451;
srom_1(32052) <= 13546806;
srom_1(32053) <= 13081972;
srom_1(32054) <= 12595130;
srom_1(32055) <= 12088561;
srom_1(32056) <= 11564642;
srom_1(32057) <= 11025830;
srom_1(32058) <= 10474651;
srom_1(32059) <= 9913689;
srom_1(32060) <= 9345576;
srom_1(32061) <= 8772976;
srom_1(32062) <= 8198573;
srom_1(32063) <= 7625061;
srom_1(32064) <= 7055130;
srom_1(32065) <= 6491451;
srom_1(32066) <= 5936670;
srom_1(32067) <= 5393386;
srom_1(32068) <= 4864148;
srom_1(32069) <= 4351437;
srom_1(32070) <= 3857658;
srom_1(32071) <= 3385126;
srom_1(32072) <= 2936057;
srom_1(32073) <= 2512557;
srom_1(32074) <= 2116612;
srom_1(32075) <= 1750078;
srom_1(32076) <= 1414674;
srom_1(32077) <= 1111974;
srom_1(32078) <= 843397;
srom_1(32079) <= 610201;
srom_1(32080) <= 413481;
srom_1(32081) <= 254160;
srom_1(32082) <= 132983;
srom_1(32083) <= 50520;
srom_1(32084) <= 7157;
srom_1(32085) <= 3098;
srom_1(32086) <= 38361;
srom_1(32087) <= 112781;
srom_1(32088) <= 226010;
srom_1(32089) <= 377515;
srom_1(32090) <= 566588;
srom_1(32091) <= 792340;
srom_1(32092) <= 1053714;
srom_1(32093) <= 1349484;
srom_1(32094) <= 1678263;
srom_1(32095) <= 2038509;
srom_1(32096) <= 2428532;
srom_1(32097) <= 2846505;
srom_1(32098) <= 3290466;
srom_1(32099) <= 3758335;
srom_1(32100) <= 4247916;
srom_1(32101) <= 4756914;
srom_1(32102) <= 5282943;
srom_1(32103) <= 5823535;
srom_1(32104) <= 6376155;
srom_1(32105) <= 6938213;
srom_1(32106) <= 7507072;
srom_1(32107) <= 8080065;
srom_1(32108) <= 8654505;
srom_1(32109) <= 9227697;
srom_1(32110) <= 9796955;
srom_1(32111) <= 10359609;
srom_1(32112) <= 10913020;
srom_1(32113) <= 11454594;
srom_1(32114) <= 11981790;
srom_1(32115) <= 12492136;
srom_1(32116) <= 12983239;
srom_1(32117) <= 13452796;
srom_1(32118) <= 13898606;
srom_1(32119) <= 14318578;
srom_1(32120) <= 14710741;
srom_1(32121) <= 15073258;
srom_1(32122) <= 15404429;
srom_1(32123) <= 15702700;
srom_1(32124) <= 15966672;
srom_1(32125) <= 16195109;
srom_1(32126) <= 16386938;
srom_1(32127) <= 16541260;
srom_1(32128) <= 16657352;
srom_1(32129) <= 16734668;
srom_1(32130) <= 16772847;
srom_1(32131) <= 16771710;
srom_1(32132) <= 16731261;
srom_1(32133) <= 16651690;
srom_1(32134) <= 16533372;
srom_1(32135) <= 16376859;
srom_1(32136) <= 16182887;
srom_1(32137) <= 15952365;
srom_1(32138) <= 15686374;
srom_1(32139) <= 15386161;
srom_1(32140) <= 15053134;
srom_1(32141) <= 14688855;
srom_1(32142) <= 14295032;
srom_1(32143) <= 13873511;
srom_1(32144) <= 13426270;
srom_1(32145) <= 12955406;
srom_1(32146) <= 12463126;
srom_1(32147) <= 11951740;
srom_1(32148) <= 11423644;
srom_1(32149) <= 10881317;
srom_1(32150) <= 10327300;
srom_1(32151) <= 9764192;
srom_1(32152) <= 9194633;
srom_1(32153) <= 8621295;
srom_1(32154) <= 8046866;
srom_1(32155) <= 7474039;
srom_1(32156) <= 6905501;
srom_1(32157) <= 6343917;
srom_1(32158) <= 5791922;
srom_1(32159) <= 5252104;
srom_1(32160) <= 4726994;
srom_1(32161) <= 4219054;
srom_1(32162) <= 3730667;
srom_1(32163) <= 3264122;
srom_1(32164) <= 2821608;
srom_1(32165) <= 2405199;
srom_1(32166) <= 2016849;
srom_1(32167) <= 1658378;
srom_1(32168) <= 1331468;
srom_1(32169) <= 1037651;
srom_1(32170) <= 778305;
srom_1(32171) <= 554646;
srom_1(32172) <= 367723;
srom_1(32173) <= 218413;
srom_1(32174) <= 107416;
srom_1(32175) <= 35253;
srom_1(32176) <= 2261;
srom_1(32177) <= 8595;
srom_1(32178) <= 54226;
srom_1(32179) <= 138940;
srom_1(32180) <= 262340;
srom_1(32181) <= 423846;
srom_1(32182) <= 622702;
srom_1(32183) <= 857975;
srom_1(32184) <= 1128562;
srom_1(32185) <= 1433193;
srom_1(32186) <= 1770441;
srom_1(32187) <= 2138723;
srom_1(32188) <= 2536314;
srom_1(32189) <= 2961348;
srom_1(32190) <= 3411832;
srom_1(32191) <= 3885654;
srom_1(32192) <= 4380592;
srom_1(32193) <= 4894325;
srom_1(32194) <= 5424443;
srom_1(32195) <= 5968462;
srom_1(32196) <= 6523829;
srom_1(32197) <= 7087942;
srom_1(32198) <= 7658153;
srom_1(32199) <= 8231790;
srom_1(32200) <= 8806162;
srom_1(32201) <= 9378576;
srom_1(32202) <= 9946348;
srom_1(32203) <= 10506815;
srom_1(32204) <= 11057349;
srom_1(32205) <= 11595368;
srom_1(32206) <= 12118350;
srom_1(32207) <= 12623841;
srom_1(32208) <= 13109473;
srom_1(32209) <= 13572966;
srom_1(32210) <= 14012148;
srom_1(32211) <= 14424960;
srom_1(32212) <= 14809465;
srom_1(32213) <= 15163860;
srom_1(32214) <= 15486484;
srom_1(32215) <= 15775823;
srom_1(32216) <= 16030522;
srom_1(32217) <= 16249384;
srom_1(32218) <= 16431385;
srom_1(32219) <= 16575670;
srom_1(32220) <= 16681564;
srom_1(32221) <= 16748569;
srom_1(32222) <= 16776371;
srom_1(32223) <= 16764840;
srom_1(32224) <= 16714030;
srom_1(32225) <= 16624180;
srom_1(32226) <= 16495710;
srom_1(32227) <= 16329222;
srom_1(32228) <= 16125499;
srom_1(32229) <= 15885495;
srom_1(32230) <= 15610335;
srom_1(32231) <= 15301310;
srom_1(32232) <= 14959869;
srom_1(32233) <= 14587613;
srom_1(32234) <= 14186288;
srom_1(32235) <= 13757775;
srom_1(32236) <= 13304085;
srom_1(32237) <= 12827344;
srom_1(32238) <= 12329789;
srom_1(32239) <= 11813751;
srom_1(32240) <= 11281653;
srom_1(32241) <= 10735987;
srom_1(32242) <= 10179314;
srom_1(32243) <= 9614244;
srom_1(32244) <= 9043427;
srom_1(32245) <= 8469538;
srom_1(32246) <= 7895271;
srom_1(32247) <= 7323316;
srom_1(32248) <= 6756357;
srom_1(32249) <= 6197053;
srom_1(32250) <= 5648025;
srom_1(32251) <= 5111849;
srom_1(32252) <= 4591038;
srom_1(32253) <= 4088036;
srom_1(32254) <= 3605201;
srom_1(32255) <= 3144796;
srom_1(32256) <= 2708982;
srom_1(32257) <= 2299801;
srom_1(32258) <= 1919173;
srom_1(32259) <= 1568882;
srom_1(32260) <= 1250572;
srom_1(32261) <= 965734;
srom_1(32262) <= 715704;
srom_1(32263) <= 501655;
srom_1(32264) <= 324591;
srom_1(32265) <= 185342;
srom_1(32266) <= 84561;
srom_1(32267) <= 22720;
srom_1(32268) <= 110;
srom_1(32269) <= 16836;
srom_1(32270) <= 72820;
srom_1(32271) <= 167800;
srom_1(32272) <= 301331;
srom_1(32273) <= 472785;
srom_1(32274) <= 681359;
srom_1(32275) <= 926075;
srom_1(32276) <= 1205786;
srom_1(32277) <= 1519179;
srom_1(32278) <= 1864785;
srom_1(32279) <= 2240984;
srom_1(32280) <= 2646011;
srom_1(32281) <= 3077967;
srom_1(32282) <= 3534827;
srom_1(32283) <= 4014447;
srom_1(32284) <= 4514580;
srom_1(32285) <= 5032879;
srom_1(32286) <= 5566914;
srom_1(32287) <= 6114181;
srom_1(32288) <= 6672114;
srom_1(32289) <= 7238096;
srom_1(32290) <= 7809473;
srom_1(32291) <= 8383566;
srom_1(32292) <= 8957683;
srom_1(32293) <= 9529130;
srom_1(32294) <= 10095230;
srom_1(32295) <= 10653327;
srom_1(32296) <= 11200803;
srom_1(32297) <= 11735093;
srom_1(32298) <= 12253689;
srom_1(32299) <= 12754161;
srom_1(32300) <= 13234161;
srom_1(32301) <= 13691438;
srom_1(32302) <= 14123849;
srom_1(32303) <= 14529366;
srom_1(32304) <= 14906086;
srom_1(32305) <= 15252243;
srom_1(32306) <= 15566215;
srom_1(32307) <= 15846528;
srom_1(32308) <= 16091869;
srom_1(32309) <= 16301086;
srom_1(32310) <= 16473199;
srom_1(32311) <= 16607400;
srom_1(32312) <= 16703061;
srom_1(32313) <= 16759733;
srom_1(32314) <= 16777149;
srom_1(32315) <= 16755229;
srom_1(32316) <= 16694074;
srom_1(32317) <= 16593973;
srom_1(32318) <= 16455393;
srom_1(32319) <= 16278986;
srom_1(32320) <= 16065578;
srom_1(32321) <= 15816170;
srom_1(32322) <= 15531932;
srom_1(32323) <= 15214196;
srom_1(32324) <= 14864452;
srom_1(32325) <= 14484342;
srom_1(32326) <= 14075646;
srom_1(32327) <= 13640281;
srom_1(32328) <= 13180290;
srom_1(32329) <= 12697829;
srom_1(32330) <= 12195161;
srom_1(32331) <= 11674642;
srom_1(32332) <= 11138714;
srom_1(32333) <= 10589890;
srom_1(32334) <= 10030743;
srom_1(32335) <= 9463895;
srom_1(32336) <= 8892005;
srom_1(32337) <= 8317755;
srom_1(32338) <= 7743837;
srom_1(32339) <= 7172942;
srom_1(32340) <= 6607748;
srom_1(32341) <= 6050905;
srom_1(32342) <= 5505025;
srom_1(32343) <= 4972666;
srom_1(32344) <= 4456326;
srom_1(32345) <= 3958426;
srom_1(32346) <= 3481301;
srom_1(32347) <= 3027187;
srom_1(32348) <= 2598215;
srom_1(32349) <= 2196396;
srom_1(32350) <= 1823615;
srom_1(32351) <= 1481619;
srom_1(32352) <= 1172012;
srom_1(32353) <= 896247;
srom_1(32354) <= 655615;
srom_1(32355) <= 451247;
srom_1(32356) <= 284099;
srom_1(32357) <= 154956;
srom_1(32358) <= 64424;
srom_1(32359) <= 12926;
srom_1(32360) <= 705;
srom_1(32361) <= 27818;
srom_1(32362) <= 94137;
srom_1(32363) <= 199352;
srom_1(32364) <= 342969;
srom_1(32365) <= 524315;
srom_1(32366) <= 742539;
srom_1(32367) <= 996619;
srom_1(32368) <= 1285362;
srom_1(32369) <= 1607414;
srom_1(32370) <= 1961266;
srom_1(32371) <= 2345258;
srom_1(32372) <= 2757589;
srom_1(32373) <= 3196326;
srom_1(32374) <= 3659411;
srom_1(32375) <= 4144673;
srom_1(32376) <= 4649836;
srom_1(32377) <= 5172532;
srom_1(32378) <= 5710309;
srom_1(32379) <= 6260646;
srom_1(32380) <= 6820961;
srom_1(32381) <= 7388627;
srom_1(32382) <= 7960983;
srom_1(32383) <= 8535344;
srom_1(32384) <= 9109017;
srom_1(32385) <= 9679312;
srom_1(32386) <= 10243554;
srom_1(32387) <= 10799097;
srom_1(32388) <= 11343337;
srom_1(32389) <= 11873721;
srom_1(32390) <= 12387763;
srom_1(32391) <= 12883051;
srom_1(32392) <= 13357262;
srom_1(32393) <= 13808175;
srom_1(32394) <= 14233673;
srom_1(32395) <= 14631761;
srom_1(32396) <= 15000573;
srom_1(32397) <= 15338380;
srom_1(32398) <= 15643596;
srom_1(32399) <= 15914791;
srom_1(32400) <= 16150694;
srom_1(32401) <= 16350197;
srom_1(32402) <= 16512366;
srom_1(32403) <= 16636440;
srom_1(32404) <= 16721836;
srom_1(32405) <= 16768156;
srom_1(32406) <= 16775180;
srom_1(32407) <= 16742878;
srom_1(32408) <= 16671399;
srom_1(32409) <= 16561079;
srom_1(32410) <= 16412436;
srom_1(32411) <= 16226166;
srom_1(32412) <= 16003144;
srom_1(32413) <= 15744414;
srom_1(32414) <= 15451190;
srom_1(32415) <= 15124847;
srom_1(32416) <= 14766916;
srom_1(32417) <= 14379075;
srom_1(32418) <= 13963142;
srom_1(32419) <= 13521068;
srom_1(32420) <= 13054927;
srom_1(32421) <= 12566903;
srom_1(32422) <= 12059287;
srom_1(32423) <= 11534457;
srom_1(32424) <= 10994875;
srom_1(32425) <= 10443071;
srom_1(32426) <= 9881633;
srom_1(32427) <= 9313194;
srom_1(32428) <= 8740419;
srom_1(32429) <= 8165995;
srom_1(32430) <= 7592614;
srom_1(32431) <= 7022966;
srom_1(32432) <= 6459722;
srom_1(32433) <= 5905524;
srom_1(32434) <= 5362969;
srom_1(32435) <= 4834602;
srom_1(32436) <= 4322902;
srom_1(32437) <= 3830267;
srom_1(32438) <= 3359007;
srom_1(32439) <= 2911333;
srom_1(32440) <= 2489344;
srom_1(32441) <= 2095019;
srom_1(32442) <= 1730206;
srom_1(32443) <= 1396617;
srom_1(32444) <= 1095816;
srom_1(32445) <= 829213;
srom_1(32446) <= 598058;
srom_1(32447) <= 403437;
srom_1(32448) <= 246260;
srom_1(32449) <= 127266;
srom_1(32450) <= 47012;
srom_1(32451) <= 5874;
srom_1(32452) <= 4047;
srom_1(32453) <= 41537;
srom_1(32454) <= 118169;
srom_1(32455) <= 233585;
srom_1(32456) <= 387242;
srom_1(32457) <= 578420;
srom_1(32458) <= 806223;
srom_1(32459) <= 1069582;
srom_1(32460) <= 1367263;
srom_1(32461) <= 1697869;
srom_1(32462) <= 2059850;
srom_1(32463) <= 2451509;
srom_1(32464) <= 2871010;
srom_1(32465) <= 3316384;
srom_1(32466) <= 3785543;
srom_1(32467) <= 4276288;
srom_1(32468) <= 4786317;
srom_1(32469) <= 5313238;
srom_1(32470) <= 5854581;
srom_1(32471) <= 6407807;
srom_1(32472) <= 6970321;
srom_1(32473) <= 7539486;
srom_1(32474) <= 8112633;
srom_1(32475) <= 8687074;
srom_1(32476) <= 9260115;
srom_1(32477) <= 9829070;
srom_1(32478) <= 10391270;
srom_1(32479) <= 10944079;
srom_1(32480) <= 11484904;
srom_1(32481) <= 12011209;
srom_1(32482) <= 12520527;
srom_1(32483) <= 13010469;
srom_1(32484) <= 13478738;
srom_1(32485) <= 13923137;
srom_1(32486) <= 14341582;
srom_1(32487) <= 14732113;
srom_1(32488) <= 15092896;
srom_1(32489) <= 15422240;
srom_1(32490) <= 15718602;
srom_1(32491) <= 15980591;
srom_1(32492) <= 16206978;
srom_1(32493) <= 16396702;
srom_1(32494) <= 16548873;
srom_1(32495) <= 16662778;
srom_1(32496) <= 16737883;
srom_1(32497) <= 16773835;
srom_1(32498) <= 16770466;
srom_1(32499) <= 16727792;
srom_1(32500) <= 16646012;
srom_1(32501) <= 16525510;
srom_1(32502) <= 16366852;
srom_1(32503) <= 16170781;
srom_1(32504) <= 15938216;
srom_1(32505) <= 15670249;
srom_1(32506) <= 15368136;
srom_1(32507) <= 15033293;
srom_1(32508) <= 14667291;
srom_1(32509) <= 14271846;
srom_1(32510) <= 13848813;
srom_1(32511) <= 13400175;
srom_1(32512) <= 12928036;
srom_1(32513) <= 12434610;
srom_1(32514) <= 11922211;
srom_1(32515) <= 11393241;
srom_1(32516) <= 10850182;
srom_1(32517) <= 10295580;
srom_1(32518) <= 9732035;
srom_1(32519) <= 9162190;
srom_1(32520) <= 8588718;
srom_1(32521) <= 8014308;
srom_1(32522) <= 7441652;
srom_1(32523) <= 6873437;
srom_1(32524) <= 6312328;
srom_1(32525) <= 5760955;
srom_1(32526) <= 5221903;
srom_1(32527) <= 4697702;
srom_1(32528) <= 4190808;
srom_1(32529) <= 3703599;
srom_1(32530) <= 3238360;
srom_1(32531) <= 2797273;
srom_1(32532) <= 2382404;
srom_1(32533) <= 1995701;
srom_1(32534) <= 1638977;
srom_1(32535) <= 1313904;
srom_1(32536) <= 1022007;
srom_1(32537) <= 764654;
srom_1(32538) <= 543052;
srom_1(32539) <= 358241;
srom_1(32540) <= 211087;
srom_1(32541) <= 102280;
srom_1(32542) <= 32331;
srom_1(32543) <= 1567;
srom_1(32544) <= 10133;
srom_1(32545) <= 57989;
srom_1(32546) <= 144909;
srom_1(32547) <= 270487;
srom_1(32548) <= 434134;
srom_1(32549) <= 635082;
srom_1(32550) <= 872389;
srom_1(32551) <= 1144942;
srom_1(32552) <= 1451463;
srom_1(32553) <= 1790515;
srom_1(32554) <= 2160507;
srom_1(32555) <= 2559705;
srom_1(32556) <= 2986237;
srom_1(32557) <= 3438103;
srom_1(32558) <= 3913183;
srom_1(32559) <= 4409249;
srom_1(32560) <= 4923977;
srom_1(32561) <= 5454951;
srom_1(32562) <= 5999682;
srom_1(32563) <= 6555616;
srom_1(32564) <= 7120145;
srom_1(32565) <= 7690623;
srom_1(32566) <= 8264373;
srom_1(32567) <= 8838706;
srom_1(32568) <= 9410929;
srom_1(32569) <= 9978357;
srom_1(32570) <= 10538330;
srom_1(32571) <= 11088223;
srom_1(32572) <= 11625456;
srom_1(32573) <= 12147511;
srom_1(32574) <= 12651939;
srom_1(32575) <= 13136374;
srom_1(32576) <= 13598546;
srom_1(32577) <= 14036287;
srom_1(32578) <= 14447543;
srom_1(32579) <= 14830387;
srom_1(32580) <= 15183024;
srom_1(32581) <= 15503799;
srom_1(32582) <= 15791208;
srom_1(32583) <= 16043904;
srom_1(32584) <= 16260702;
srom_1(32585) <= 16440585;
srom_1(32586) <= 16582709;
srom_1(32587) <= 16686408;
srom_1(32588) <= 16751197;
srom_1(32589) <= 16776770;
srom_1(32590) <= 16763008;
srom_1(32591) <= 16709975;
srom_1(32592) <= 16617921;
srom_1(32593) <= 16487277;
srom_1(32594) <= 16318655;
srom_1(32595) <= 16112847;
srom_1(32596) <= 15870817;
srom_1(32597) <= 15593700;
srom_1(32598) <= 15282797;
srom_1(32599) <= 14939564;
srom_1(32600) <= 14565611;
srom_1(32601) <= 14162692;
srom_1(32602) <= 13732697;
srom_1(32603) <= 13277641;
srom_1(32604) <= 12799659;
srom_1(32605) <= 12300992;
srom_1(32606) <= 11783978;
srom_1(32607) <= 11251042;
srom_1(32608) <= 10704684;
srom_1(32609) <= 10147464;
srom_1(32610) <= 9581997;
srom_1(32611) <= 9010933;
srom_1(32612) <= 8436952;
srom_1(32613) <= 7862743;
srom_1(32614) <= 7291000;
srom_1(32615) <= 6724405;
srom_1(32616) <= 6165613;
srom_1(32617) <= 5617246;
srom_1(32618) <= 5081875;
srom_1(32619) <= 4562010;
srom_1(32620) <= 4060089;
srom_1(32621) <= 3578466;
srom_1(32622) <= 3119400;
srom_1(32623) <= 2685043;
srom_1(32624) <= 2277431;
srom_1(32625) <= 1898477;
srom_1(32626) <= 1549958;
srom_1(32627) <= 1233507;
srom_1(32628) <= 950609;
srom_1(32629) <= 702591;
srom_1(32630) <= 490614;
srom_1(32631) <= 315674;
srom_1(32632) <= 178591;
srom_1(32633) <= 80008;
srom_1(32634) <= 20386;
srom_1(32635) <= 6;
srom_1(32636) <= 18963;
srom_1(32637) <= 77168;
srom_1(32638) <= 174348;
srom_1(32639) <= 310048;
srom_1(32640) <= 483630;
srom_1(32641) <= 694282;
srom_1(32642) <= 941015;
srom_1(32643) <= 1222673;
srom_1(32644) <= 1537934;
srom_1(32645) <= 1885320;
srom_1(32646) <= 2263203;
srom_1(32647) <= 2669809;
srom_1(32648) <= 3103233;
srom_1(32649) <= 3561442;
srom_1(32650) <= 4042287;
srom_1(32651) <= 4543514;
srom_1(32652) <= 5062771;
srom_1(32653) <= 5597624;
srom_1(32654) <= 6145566;
srom_1(32655) <= 6704025;
srom_1(32656) <= 7270385;
srom_1(32657) <= 7841988;
srom_1(32658) <= 8416154;
srom_1(32659) <= 8990191;
srom_1(32660) <= 9561407;
srom_1(32661) <= 10127123;
srom_1(32662) <= 10684687;
srom_1(32663) <= 11231484;
srom_1(32664) <= 11764950;
srom_1(32665) <= 12282582;
srom_1(32666) <= 12781955;
srom_1(32667) <= 13260725;
srom_1(32668) <= 13716649;
srom_1(32669) <= 14147588;
srom_1(32670) <= 14551520;
srom_1(32671) <= 14926553;
srom_1(32672) <= 15270927;
srom_1(32673) <= 15583027;
srom_1(32674) <= 15861391;
srom_1(32675) <= 16104712;
srom_1(32676) <= 16311849;
srom_1(32677) <= 16481832;
srom_1(32678) <= 16613862;
srom_1(32679) <= 16707322;
srom_1(32680) <= 16761772;
srom_1(32681) <= 16776958;
srom_1(32682) <= 16752808;
srom_1(32683) <= 16689435;
srom_1(32684) <= 16587137;
srom_1(32685) <= 16446393;
srom_1(32686) <= 16267863;
srom_1(32687) <= 16052385;
srom_1(32688) <= 15800968;
srom_1(32689) <= 15514793;
srom_1(32690) <= 15195200;
srom_1(32691) <= 14843689;
srom_1(32692) <= 14461908;
srom_1(32693) <= 14051647;
srom_1(32694) <= 13614830;
srom_1(32695) <= 13153506;
srom_1(32696) <= 12669837;
srom_1(32697) <= 12166092;
srom_1(32698) <= 11644634;
srom_1(32699) <= 11107906;
srom_1(32700) <= 10558427;
srom_1(32701) <= 9998773;
srom_1(32702) <= 9431568;
srom_1(32703) <= 8859473;
srom_1(32704) <= 8285169;
srom_1(32705) <= 7711350;
srom_1(32706) <= 7140708;
srom_1(32707) <= 6575917;
srom_1(32708) <= 6019626;
srom_1(32709) <= 5474445;
srom_1(32710) <= 4942929;
srom_1(32711) <= 4427570;
srom_1(32712) <= 3930787;
srom_1(32713) <= 3454908;
srom_1(32714) <= 3002164;
srom_1(32715) <= 2574680;
srom_1(32716) <= 2174459;
srom_1(32717) <= 1803378;
srom_1(32718) <= 1463178;
srom_1(32719) <= 1155453;
srom_1(32720) <= 881647;
srom_1(32721) <= 643044;
srom_1(32722) <= 440762;
srom_1(32723) <= 275751;
srom_1(32724) <= 148783;
srom_1(32725) <= 60455;
srom_1(32726) <= 11181;
srom_1(32727) <= 1191;
srom_1(32728) <= 30533;
srom_1(32729) <= 99068;
srom_1(32730) <= 206476;
srom_1(32731) <= 352253;
srom_1(32732) <= 535715;
srom_1(32733) <= 756002;
srom_1(32734) <= 1012080;
srom_1(32735) <= 1302750;
srom_1(32736) <= 1626648;
srom_1(32737) <= 1982255;
srom_1(32738) <= 2367904;
srom_1(32739) <= 2781786;
srom_1(32740) <= 3221960;
srom_1(32741) <= 3686362;
srom_1(32742) <= 4172815;
srom_1(32743) <= 4679037;
srom_1(32744) <= 5202654;
srom_1(32745) <= 5741212;
srom_1(32746) <= 6292184;
srom_1(32747) <= 6852986;
srom_1(32748) <= 7420990;
srom_1(32749) <= 7993532;
srom_1(32750) <= 8567926;
srom_1(32751) <= 9141479;
srom_1(32752) <= 9711502;
srom_1(32753) <= 10275321;
srom_1(32754) <= 10830292;
srom_1(32755) <= 11373814;
srom_1(32756) <= 11903337;
srom_1(32757) <= 12416379;
srom_1(32758) <= 12910532;
srom_1(32759) <= 13383481;
srom_1(32760) <= 13833007;
srom_1(32761) <= 14257003;
srom_1(32762) <= 14653480;
srom_1(32763) <= 15020578;
srom_1(32764) <= 15356577;
srom_1(32765) <= 15659901;
srom_1(32766) <= 15929127;
srom_1(32767) <= 16162993;
srom_1(32768) <= 16360402;
srom_1(32769) <= 16520429;
srom_1(32770) <= 16642322;
srom_1(32771) <= 16725512;
srom_1(32772) <= 16769606;
srom_1(32773) <= 16774400;
srom_1(32774) <= 16739869;
srom_1(32775) <= 16666177;
srom_1(32776) <= 16553668;
srom_1(32777) <= 16402870;
srom_1(32778) <= 16214491;
srom_1(32779) <= 15989413;
srom_1(32780) <= 15728693;
srom_1(32781) <= 15433552;
srom_1(32782) <= 15105376;
srom_1(32783) <= 14745702;
srom_1(32784) <= 14356217;
srom_1(32785) <= 13938749;
srom_1(32786) <= 13495253;
srom_1(32787) <= 13027811;
srom_1(32788) <= 12538614;
srom_1(32789) <= 12029957;
srom_1(32790) <= 11504223;
srom_1(32791) <= 10963880;
srom_1(32792) <= 10411460;
srom_1(32793) <= 9849555;
srom_1(32794) <= 9280798;
srom_1(32795) <= 8707858;
srom_1(32796) <= 8133420;
srom_1(32797) <= 7560180;
srom_1(32798) <= 6990824;
srom_1(32799) <= 6428022;
srom_1(32800) <= 5874415;
srom_1(32801) <= 5332597;
srom_1(32802) <= 4805111;
srom_1(32803) <= 4294428;
srom_1(32804) <= 3802944;
srom_1(32805) <= 3332965;
srom_1(32806) <= 2886692;
srom_1(32807) <= 2466220;
srom_1(32808) <= 2073521;
srom_1(32809) <= 1710435;
srom_1(32810) <= 1378665;
srom_1(32811) <= 1079767;
srom_1(32812) <= 815143;
srom_1(32813) <= 586033;
srom_1(32814) <= 393512;
srom_1(32815) <= 238483;
srom_1(32816) <= 121673;
srom_1(32817) <= 43630;
srom_1(32818) <= 4718;
srom_1(32819) <= 5122;
srom_1(32820) <= 44839;
srom_1(32821) <= 123682;
srom_1(32822) <= 241283;
srom_1(32823) <= 397089;
srom_1(32824) <= 590370;
srom_1(32825) <= 820220;
srom_1(32826) <= 1085560;
srom_1(32827) <= 1385147;
srom_1(32828) <= 1717576;
srom_1(32829) <= 2081288;
srom_1(32830) <= 2474576;
srom_1(32831) <= 2895598;
srom_1(32832) <= 3342378;
srom_1(32833) <= 3812821;
srom_1(32834) <= 4304722;
srom_1(32835) <= 4815774;
srom_1(32836) <= 5343580;
srom_1(32837) <= 5885665;
srom_1(32838) <= 6439488;
srom_1(32839) <= 7002450;
srom_1(32840) <= 7571913;
srom_1(32841) <= 8145205;
srom_1(32842) <= 8719639;
srom_1(32843) <= 9292520;
srom_1(32844) <= 9861163;
srom_1(32845) <= 10422900;
srom_1(32846) <= 10975098;
srom_1(32847) <= 11515167;
srom_1(32848) <= 12040574;
srom_1(32849) <= 12548856;
srom_1(32850) <= 13037630;
srom_1(32851) <= 13504602;
srom_1(32852) <= 13947584;
srom_1(32853) <= 14364497;
srom_1(32854) <= 14753388;
srom_1(32855) <= 15112432;
srom_1(32856) <= 15439946;
srom_1(32857) <= 15734393;
srom_1(32858) <= 15994394;
srom_1(32859) <= 16218729;
srom_1(32860) <= 16406345;
srom_1(32861) <= 16556363;
srom_1(32862) <= 16668080;
srom_1(32863) <= 16740972;
srom_1(32864) <= 16774697;
srom_1(32865) <= 16769096;
srom_1(32866) <= 16724197;
srom_1(32867) <= 16640208;
srom_1(32868) <= 16517526;
srom_1(32869) <= 16356724;
srom_1(32870) <= 16158557;
srom_1(32871) <= 15923953;
srom_1(32872) <= 15654014;
srom_1(32873) <= 15350005;
srom_1(32874) <= 15013352;
srom_1(32875) <= 14645633;
srom_1(32876) <= 14248573;
srom_1(32877) <= 13824033;
srom_1(32878) <= 13374004;
srom_1(32879) <= 12900598;
srom_1(32880) <= 12406033;
srom_1(32881) <= 11892629;
srom_1(32882) <= 11362793;
srom_1(32883) <= 10819010;
srom_1(32884) <= 10263831;
srom_1(32885) <= 9699858;
srom_1(32886) <= 9129736;
srom_1(32887) <= 8556138;
srom_1(32888) <= 7981755;
srom_1(32889) <= 7409280;
srom_1(32890) <= 6841397;
srom_1(32891) <= 6280770;
srom_1(32892) <= 5730027;
srom_1(32893) <= 5191751;
srom_1(32894) <= 4668466;
srom_1(32895) <= 4162626;
srom_1(32896) <= 3676603;
srom_1(32897) <= 3212676;
srom_1(32898) <= 2773022;
srom_1(32899) <= 2359700;
srom_1(32900) <= 1974650;
srom_1(32901) <= 1619678;
srom_1(32902) <= 1296447;
srom_1(32903) <= 1006474;
srom_1(32904) <= 751118;
srom_1(32905) <= 531577;
srom_1(32906) <= 348880;
srom_1(32907) <= 203884;
srom_1(32908) <= 97270;
srom_1(32909) <= 29536;
srom_1(32910) <= 1001;
srom_1(32911) <= 11798;
srom_1(32912) <= 61877;
srom_1(32913) <= 151002;
srom_1(32914) <= 278757;
srom_1(32915) <= 444542;
srom_1(32916) <= 647579;
srom_1(32917) <= 886916;
srom_1(32918) <= 1161431;
srom_1(32919) <= 1469837;
srom_1(32920) <= 1810688;
srom_1(32921) <= 2182385;
srom_1(32922) <= 2583185;
srom_1(32923) <= 3011208;
srom_1(32924) <= 3464448;
srom_1(32925) <= 3940779;
srom_1(32926) <= 4437967;
srom_1(32927) <= 4953681;
srom_1(32928) <= 5485503;
srom_1(32929) <= 6030939;
srom_1(32930) <= 6587430;
srom_1(32931) <= 7152368;
srom_1(32932) <= 7723103;
srom_1(32933) <= 8296958;
srom_1(32934) <= 8871244;
srom_1(32935) <= 9443266;
srom_1(32936) <= 10010342;
srom_1(32937) <= 10569814;
srom_1(32938) <= 11119057;
srom_1(32939) <= 11655496;
srom_1(32940) <= 12176616;
srom_1(32941) <= 12679972;
srom_1(32942) <= 13163205;
srom_1(32943) <= 13624048;
srom_1(32944) <= 14060340;
srom_1(32945) <= 14470035;
srom_1(32946) <= 14851213;
srom_1(32947) <= 15202085;
srom_1(32948) <= 15521006;
srom_1(32949) <= 15806481;
srom_1(32950) <= 16057171;
srom_1(32951) <= 16271901;
srom_1(32952) <= 16449663;
srom_1(32953) <= 16589624;
srom_1(32954) <= 16691128;
srom_1(32955) <= 16753698;
srom_1(32956) <= 16777042;
srom_1(32957) <= 16761049;
srom_1(32958) <= 16705795;
srom_1(32959) <= 16611539;
srom_1(32960) <= 16478722;
srom_1(32961) <= 16307969;
srom_1(32962) <= 16100079;
srom_1(32963) <= 15856027;
srom_1(32964) <= 15576957;
srom_1(32965) <= 15264179;
srom_1(32966) <= 14919159;
srom_1(32967) <= 14543516;
srom_1(32968) <= 14139009;
srom_1(32969) <= 13707537;
srom_1(32970) <= 13251123;
srom_1(32971) <= 12771907;
srom_1(32972) <= 12272136;
srom_1(32973) <= 11754153;
srom_1(32974) <= 11220389;
srom_1(32975) <= 10673345;
srom_1(32976) <= 10115588;
srom_1(32977) <= 9549732;
srom_1(32978) <= 8978431;
srom_1(32979) <= 8404364;
srom_1(32980) <= 7830223;
srom_1(32981) <= 7258701;
srom_1(32982) <= 6692477;
srom_1(32983) <= 6134207;
srom_1(32984) <= 5586509;
srom_1(32985) <= 5051951;
srom_1(32986) <= 4533039;
srom_1(32987) <= 4032207;
srom_1(32988) <= 3551804;
srom_1(32989) <= 3094083;
srom_1(32990) <= 2661189;
srom_1(32991) <= 2255154;
srom_1(32992) <= 1877880;
srom_1(32993) <= 1531137;
srom_1(32994) <= 1216551;
srom_1(32995) <= 935597;
srom_1(32996) <= 689593;
srom_1(32997) <= 479693;
srom_1(32998) <= 306880;
srom_1(32999) <= 171965;
srom_1(33000) <= 75580;
srom_1(33001) <= 18179;
srom_1(33002) <= 29;
srom_1(33003) <= 21216;
srom_1(33004) <= 81640;
srom_1(33005) <= 181019;
srom_1(33006) <= 318886;
srom_1(33007) <= 494595;
srom_1(33008) <= 707321;
srom_1(33009) <= 956068;
srom_1(33010) <= 1239668;
srom_1(33011) <= 1556793;
srom_1(33012) <= 1905954;
srom_1(33013) <= 2285514;
srom_1(33014) <= 2693694;
srom_1(33015) <= 3128579;
srom_1(33016) <= 3588130;
srom_1(33017) <= 4070192;
srom_1(33018) <= 4572505;
srom_1(33019) <= 5092713;
srom_1(33020) <= 5628377;
srom_1(33021) <= 6176984;
srom_1(33022) <= 6735962;
srom_1(33023) <= 7302690;
srom_1(33024) <= 7874510;
srom_1(33025) <= 8448741;
srom_1(33026) <= 9022690;
srom_1(33027) <= 9593666;
srom_1(33028) <= 10158991;
srom_1(33029) <= 10716013;
srom_1(33030) <= 11262122;
srom_1(33031) <= 11794756;
srom_1(33032) <= 12311417;
srom_1(33033) <= 12809683;
srom_1(33034) <= 13287217;
srom_1(33035) <= 13741779;
srom_1(33036) <= 14171239;
srom_1(33037) <= 14573582;
srom_1(33038) <= 14946921;
srom_1(33039) <= 15289507;
srom_1(33040) <= 15599731;
srom_1(33041) <= 15876140;
srom_1(33042) <= 16117438;
srom_1(33043) <= 16322492;
srom_1(33044) <= 16490342;
srom_1(33045) <= 16620200;
srom_1(33046) <= 16711457;
srom_1(33047) <= 16763685;
srom_1(33048) <= 16776640;
srom_1(33049) <= 16750261;
srom_1(33050) <= 16684670;
srom_1(33051) <= 16580177;
srom_1(33052) <= 16437270;
srom_1(33053) <= 16256621;
srom_1(33054) <= 16039076;
srom_1(33055) <= 15785655;
srom_1(33056) <= 15497547;
srom_1(33057) <= 15176102;
srom_1(33058) <= 14822829;
srom_1(33059) <= 14439383;
srom_1(33060) <= 14027563;
srom_1(33061) <= 13589301;
srom_1(33062) <= 13126650;
srom_1(33063) <= 12641781;
srom_1(33064) <= 12136967;
srom_1(33065) <= 11614576;
srom_1(33066) <= 11077058;
srom_1(33067) <= 10526932;
srom_1(33068) <= 9966779;
srom_1(33069) <= 9399225;
srom_1(33070) <= 8826933;
srom_1(33071) <= 8252584;
srom_1(33072) <= 7678874;
srom_1(33073) <= 7108492;
srom_1(33074) <= 6544113;
srom_1(33075) <= 5988383;
srom_1(33076) <= 5443908;
srom_1(33077) <= 4913243;
srom_1(33078) <= 4398874;
srom_1(33079) <= 3903215;
srom_1(33080) <= 3428589;
srom_1(33081) <= 2977223;
srom_1(33082) <= 2551232;
srom_1(33083) <= 2152615;
srom_1(33084) <= 1783241;
srom_1(33085) <= 1444841;
srom_1(33086) <= 1139003;
srom_1(33087) <= 867161;
srom_1(33088) <= 630589;
srom_1(33089) <= 430398;
srom_1(33090) <= 267525;
srom_1(33091) <= 142735;
srom_1(33092) <= 56613;
srom_1(33093) <= 9562;
srom_1(33094) <= 1803;
srom_1(33095) <= 33374;
srom_1(33096) <= 104124;
srom_1(33097) <= 213723;
srom_1(33098) <= 361658;
srom_1(33099) <= 547233;
srom_1(33100) <= 769579;
srom_1(33101) <= 1027654;
srom_1(33102) <= 1320246;
srom_1(33103) <= 1645985;
srom_1(33104) <= 2003341;
srom_1(33105) <= 2390641;
srom_1(33106) <= 2806067;
srom_1(33107) <= 3247672;
srom_1(33108) <= 3713384;
srom_1(33109) <= 4201020;
srom_1(33110) <= 4708293;
srom_1(33111) <= 5232824;
srom_1(33112) <= 5772154;
srom_1(33113) <= 6323753;
srom_1(33114) <= 6885035;
srom_1(33115) <= 7453368;
srom_1(33116) <= 8026086;
srom_1(33117) <= 8600505;
srom_1(33118) <= 9173929;
srom_1(33119) <= 9743671;
srom_1(33120) <= 10307059;
srom_1(33121) <= 10861451;
srom_1(33122) <= 11404246;
srom_1(33123) <= 11932900;
srom_1(33124) <= 12444934;
srom_1(33125) <= 12937946;
srom_1(33126) <= 13409625;
srom_1(33127) <= 13857758;
srom_1(33128) <= 14280245;
srom_1(33129) <= 14675104;
srom_1(33130) <= 15040483;
srom_1(33131) <= 15374669;
srom_1(33132) <= 15676095;
srom_1(33133) <= 15943348;
srom_1(33134) <= 16175174;
srom_1(33135) <= 16370486;
srom_1(33136) <= 16528369;
srom_1(33137) <= 16648081;
srom_1(33138) <= 16729061;
srom_1(33139) <= 16770931;
srom_1(33140) <= 16773492;
srom_1(33141) <= 16736735;
srom_1(33142) <= 16660830;
srom_1(33143) <= 16546133;
srom_1(33144) <= 16393183;
srom_1(33145) <= 16202697;
srom_1(33146) <= 15975568;
srom_1(33147) <= 15712861;
srom_1(33148) <= 15415809;
srom_1(33149) <= 15085803;
srom_1(33150) <= 14724392;
srom_1(33151) <= 14333270;
srom_1(33152) <= 13914271;
srom_1(33153) <= 13469361;
srom_1(33154) <= 13000626;
srom_1(33155) <= 12510263;
srom_1(33156) <= 12000572;
srom_1(33157) <= 11473943;
srom_1(33158) <= 10932846;
srom_1(33159) <= 10379819;
srom_1(33160) <= 9817454;
srom_1(33161) <= 9248388;
srom_1(33162) <= 8675291;
srom_1(33163) <= 8100850;
srom_1(33164) <= 7527757;
srom_1(33165) <= 6958702;
srom_1(33166) <= 6396352;
srom_1(33167) <= 5843344;
srom_1(33168) <= 5302272;
srom_1(33169) <= 4775673;
srom_1(33170) <= 4266016;
srom_1(33171) <= 3775691;
srom_1(33172) <= 3306998;
srom_1(33173) <= 2862134;
srom_1(33174) <= 2443186;
srom_1(33175) <= 2052118;
srom_1(33176) <= 1690764;
srom_1(33177) <= 1360818;
srom_1(33178) <= 1063829;
srom_1(33179) <= 801187;
srom_1(33180) <= 574126;
srom_1(33181) <= 383709;
srom_1(33182) <= 230830;
srom_1(33183) <= 116205;
srom_1(33184) <= 40373;
srom_1(33185) <= 3689;
srom_1(33186) <= 6324;
srom_1(33187) <= 48267;
srom_1(33188) <= 129320;
srom_1(33189) <= 249104;
srom_1(33190) <= 407057;
srom_1(33191) <= 602438;
srom_1(33192) <= 834331;
srom_1(33193) <= 1101649;
srom_1(33194) <= 1403138;
srom_1(33195) <= 1737384;
srom_1(33196) <= 2102820;
srom_1(33197) <= 2497732;
srom_1(33198) <= 2920268;
srom_1(33199) <= 3368448;
srom_1(33200) <= 3840169;
srom_1(33201) <= 4333218;
srom_1(33202) <= 4845285;
srom_1(33203) <= 5373968;
srom_1(33204) <= 5916788;
srom_1(33205) <= 6471198;
srom_1(33206) <= 7034600;
srom_1(33207) <= 7604352;
srom_1(33208) <= 8177781;
srom_1(33209) <= 8752199;
srom_1(33210) <= 9324911;
srom_1(33211) <= 9893233;
srom_1(33212) <= 10454500;
srom_1(33213) <= 11006079;
srom_1(33214) <= 11545383;
srom_1(33215) <= 12069884;
srom_1(33216) <= 12577123;
srom_1(33217) <= 13064720;
srom_1(33218) <= 13530389;
srom_1(33219) <= 13971947;
srom_1(33220) <= 14387322;
srom_1(33221) <= 14774567;
srom_1(33222) <= 15131867;
srom_1(33223) <= 15457545;
srom_1(33224) <= 15750074;
srom_1(33225) <= 16008083;
srom_1(33226) <= 16230361;
srom_1(33227) <= 16415867;
srom_1(33228) <= 16563730;
srom_1(33229) <= 16673257;
srom_1(33230) <= 16743935;
srom_1(33231) <= 16775432;
srom_1(33232) <= 16767600;
srom_1(33233) <= 16720476;
srom_1(33234) <= 16634281;
srom_1(33235) <= 16509419;
srom_1(33236) <= 16346476;
srom_1(33237) <= 16146215;
srom_1(33238) <= 15909577;
srom_1(33239) <= 15637670;
srom_1(33240) <= 15331770;
srom_1(33241) <= 14993311;
srom_1(33242) <= 14623880;
srom_1(33243) <= 14225210;
srom_1(33244) <= 13799170;
srom_1(33245) <= 13347758;
srom_1(33246) <= 12873091;
srom_1(33247) <= 12377395;
srom_1(33248) <= 11862994;
srom_1(33249) <= 11332300;
srom_1(33250) <= 10787802;
srom_1(33251) <= 10232054;
srom_1(33252) <= 9667661;
srom_1(33253) <= 9097270;
srom_1(33254) <= 8523556;
srom_1(33255) <= 7949209;
srom_1(33256) <= 7376922;
srom_1(33257) <= 6809380;
srom_1(33258) <= 6249243;
srom_1(33259) <= 5699139;
srom_1(33260) <= 5161646;
srom_1(33261) <= 4639286;
srom_1(33262) <= 4134507;
srom_1(33263) <= 3649678;
srom_1(33264) <= 3187071;
srom_1(33265) <= 2748855;
srom_1(33266) <= 2337087;
srom_1(33267) <= 1953696;
srom_1(33268) <= 1600480;
srom_1(33269) <= 1279097;
srom_1(33270) <= 991052;
srom_1(33271) <= 737697;
srom_1(33272) <= 520220;
srom_1(33273) <= 339640;
srom_1(33274) <= 196805;
srom_1(33275) <= 92384;
srom_1(33276) <= 26867;
srom_1(33277) <= 560;
srom_1(33278) <= 13589;
srom_1(33279) <= 65890;
srom_1(33280) <= 157220;
srom_1(33281) <= 287149;
srom_1(33282) <= 455069;
srom_1(33283) <= 660192;
srom_1(33284) <= 901556;
srom_1(33285) <= 1178030;
srom_1(33286) <= 1488316;
srom_1(33287) <= 1830961;
srom_1(33288) <= 2204356;
srom_1(33289) <= 2606751;
srom_1(33290) <= 3036260;
srom_1(33291) <= 3490867;
srom_1(33292) <= 3968442;
srom_1(33293) <= 4466745;
srom_1(33294) <= 4983438;
srom_1(33295) <= 5516099;
srom_1(33296) <= 6062231;
srom_1(33297) <= 6619271;
srom_1(33298) <= 7184609;
srom_1(33299) <= 7755593;
srom_1(33300) <= 8329545;
srom_1(33301) <= 8903774;
srom_1(33302) <= 9475587;
srom_1(33303) <= 10042303;
srom_1(33304) <= 10601264;
srom_1(33305) <= 11149849;
srom_1(33306) <= 11685486;
srom_1(33307) <= 12205663;
srom_1(33308) <= 12707940;
srom_1(33309) <= 13189963;
srom_1(33310) <= 13649470;
srom_1(33311) <= 14084307;
srom_1(33312) <= 14492435;
srom_1(33313) <= 14871940;
srom_1(33314) <= 15221043;
srom_1(33315) <= 15538106;
srom_1(33316) <= 15821642;
srom_1(33317) <= 16070323;
srom_1(33318) <= 16282981;
srom_1(33319) <= 16458620;
srom_1(33320) <= 16596415;
srom_1(33321) <= 16695722;
srom_1(33322) <= 16756073;
srom_1(33323) <= 16777187;
srom_1(33324) <= 16758964;
srom_1(33325) <= 16701489;
srom_1(33326) <= 16605032;
srom_1(33327) <= 16470046;
srom_1(33328) <= 16297163;
srom_1(33329) <= 16087194;
srom_1(33330) <= 15841123;
srom_1(33331) <= 15560106;
srom_1(33332) <= 15245458;
srom_1(33333) <= 14898657;
srom_1(33334) <= 14521327;
srom_1(33335) <= 14115240;
srom_1(33336) <= 13682298;
srom_1(33337) <= 13224532;
srom_1(33338) <= 12744089;
srom_1(33339) <= 12243221;
srom_1(33340) <= 11724278;
srom_1(33341) <= 11189693;
srom_1(33342) <= 10641972;
srom_1(33343) <= 10083685;
srom_1(33344) <= 9517449;
srom_1(33345) <= 8945919;
srom_1(33346) <= 8371776;
srom_1(33347) <= 7797712;
srom_1(33348) <= 7226419;
srom_1(33349) <= 6660575;
srom_1(33350) <= 6102835;
srom_1(33351) <= 5555814;
srom_1(33352) <= 5022077;
srom_1(33353) <= 4504126;
srom_1(33354) <= 4004391;
srom_1(33355) <= 3525216;
srom_1(33356) <= 3068846;
srom_1(33357) <= 2637423;
srom_1(33358) <= 2232968;
srom_1(33359) <= 1857380;
srom_1(33360) <= 1512419;
srom_1(33361) <= 1199703;
srom_1(33362) <= 920698;
srom_1(33363) <= 676712;
srom_1(33364) <= 468890;
srom_1(33365) <= 298207;
srom_1(33366) <= 165462;
srom_1(33367) <= 71278;
srom_1(33368) <= 16098;
srom_1(33369) <= 178;
srom_1(33370) <= 23595;
srom_1(33371) <= 86239;
srom_1(33372) <= 187815;
srom_1(33373) <= 327847;
srom_1(33374) <= 505679;
srom_1(33375) <= 720477;
srom_1(33376) <= 971233;
srom_1(33377) <= 1256772;
srom_1(33378) <= 1575754;
srom_1(33379) <= 1926685;
srom_1(33380) <= 2307917;
srom_1(33381) <= 2717664;
srom_1(33382) <= 3154004;
srom_1(33383) <= 3614891;
srom_1(33384) <= 4098163;
srom_1(33385) <= 4601555;
srom_1(33386) <= 5122705;
srom_1(33387) <= 5659171;
srom_1(33388) <= 6208435;
srom_1(33389) <= 6767924;
srom_1(33390) <= 7335012;
srom_1(33391) <= 7907041;
srom_1(33392) <= 8481328;
srom_1(33393) <= 9055180;
srom_1(33394) <= 9625907;
srom_1(33395) <= 10190831;
srom_1(33396) <= 10747304;
srom_1(33397) <= 11292716;
srom_1(33398) <= 11824510;
srom_1(33399) <= 12340192;
srom_1(33400) <= 12837344;
srom_1(33401) <= 13313634;
srom_1(33402) <= 13766828;
srom_1(33403) <= 14194803;
srom_1(33404) <= 14595550;
srom_1(33405) <= 14967191;
srom_1(33406) <= 15307982;
srom_1(33407) <= 15616326;
srom_1(33408) <= 15890777;
srom_1(33409) <= 16130048;
srom_1(33410) <= 16333016;
srom_1(33411) <= 16498730;
srom_1(33412) <= 16626413;
srom_1(33413) <= 16715466;
srom_1(33414) <= 16765472;
srom_1(33415) <= 16776196;
srom_1(33416) <= 16747587;
srom_1(33417) <= 16679780;
srom_1(33418) <= 16573094;
srom_1(33419) <= 16428027;
srom_1(33420) <= 16245260;
srom_1(33421) <= 16025651;
srom_1(33422) <= 15770230;
srom_1(33423) <= 15480193;
srom_1(33424) <= 15156902;
srom_1(33425) <= 14801871;
srom_1(33426) <= 14416767;
srom_1(33427) <= 14003394;
srom_1(33428) <= 13563692;
srom_1(33429) <= 13099722;
srom_1(33430) <= 12613660;
srom_1(33431) <= 12107786;
srom_1(33432) <= 11584470;
srom_1(33433) <= 11046169;
srom_1(33434) <= 10495405;
srom_1(33435) <= 9934761;
srom_1(33436) <= 9366867;
srom_1(33437) <= 8794386;
srom_1(33438) <= 8220002;
srom_1(33439) <= 7646409;
srom_1(33440) <= 7076296;
srom_1(33441) <= 6512336;
srom_1(33442) <= 5957176;
srom_1(33443) <= 5413417;
srom_1(33444) <= 4883610;
srom_1(33445) <= 4370238;
srom_1(33446) <= 3875711;
srom_1(33447) <= 3402346;
srom_1(33448) <= 2952363;
srom_1(33449) <= 2527873;
srom_1(33450) <= 2130865;
srom_1(33451) <= 1763203;
srom_1(33452) <= 1426609;
srom_1(33453) <= 1122662;
srom_1(33454) <= 852788;
srom_1(33455) <= 618252;
srom_1(33456) <= 420154;
srom_1(33457) <= 259422;
srom_1(33458) <= 136812;
srom_1(33459) <= 52896;
srom_1(33460) <= 8070;
srom_1(33461) <= 2543;
srom_1(33462) <= 36341;
srom_1(33463) <= 109305;
srom_1(33464) <= 221094;
srom_1(33465) <= 371184;
srom_1(33466) <= 558869;
srom_1(33467) <= 783272;
srom_1(33468) <= 1043338;
srom_1(33469) <= 1337848;
srom_1(33470) <= 1665423;
srom_1(33471) <= 2024524;
srom_1(33472) <= 2413469;
srom_1(33473) <= 2830433;
srom_1(33474) <= 3273461;
srom_1(33475) <= 3740477;
srom_1(33476) <= 4229288;
srom_1(33477) <= 4737605;
srom_1(33478) <= 5263042;
srom_1(33479) <= 5803136;
srom_1(33480) <= 6355354;
srom_1(33481) <= 6917106;
srom_1(33482) <= 7485759;
srom_1(33483) <= 8058646;
srom_1(33484) <= 8633080;
srom_1(33485) <= 9206368;
srom_1(33486) <= 9775821;
srom_1(33487) <= 10338769;
srom_1(33488) <= 10892572;
srom_1(33489) <= 11434633;
srom_1(33490) <= 11962410;
srom_1(33491) <= 12473428;
srom_1(33492) <= 12965291;
srom_1(33493) <= 13435692;
srom_1(33494) <= 13882426;
srom_1(33495) <= 14303398;
srom_1(33496) <= 14696633;
srom_1(33497) <= 15060287;
srom_1(33498) <= 15392656;
srom_1(33499) <= 15692180;
srom_1(33500) <= 15957456;
srom_1(33501) <= 16187238;
srom_1(33502) <= 16380450;
srom_1(33503) <= 16536186;
srom_1(33504) <= 16653714;
srom_1(33505) <= 16732485;
srom_1(33506) <= 16772128;
srom_1(33507) <= 16772459;
srom_1(33508) <= 16733474;
srom_1(33509) <= 16655358;
srom_1(33510) <= 16538475;
srom_1(33511) <= 16383376;
srom_1(33512) <= 16190786;
srom_1(33513) <= 15961609;
srom_1(33514) <= 15696919;
srom_1(33515) <= 15397959;
srom_1(33516) <= 15066129;
srom_1(33517) <= 14702986;
srom_1(33518) <= 14310233;
srom_1(33519) <= 13889711;
srom_1(33520) <= 13443392;
srom_1(33521) <= 12973370;
srom_1(33522) <= 12481849;
srom_1(33523) <= 11971132;
srom_1(33524) <= 11443616;
srom_1(33525) <= 10901774;
srom_1(33526) <= 10348147;
srom_1(33527) <= 9785331;
srom_1(33528) <= 9215966;
srom_1(33529) <= 8642720;
srom_1(33530) <= 8068283;
srom_1(33531) <= 7495348;
srom_1(33532) <= 6926602;
srom_1(33533) <= 6364712;
srom_1(33534) <= 5812312;
srom_1(33535) <= 5271993;
srom_1(33536) <= 4746290;
srom_1(33537) <= 4237666;
srom_1(33538) <= 3748508;
srom_1(33539) <= 3281109;
srom_1(33540) <= 2837660;
srom_1(33541) <= 2420242;
srom_1(33542) <= 2030811;
srom_1(33543) <= 1671195;
srom_1(33544) <= 1343078;
srom_1(33545) <= 1048001;
srom_1(33546) <= 787346;
srom_1(33547) <= 562336;
srom_1(33548) <= 374026;
srom_1(33549) <= 223299;
srom_1(33550) <= 110862;
srom_1(33551) <= 37243;
srom_1(33552) <= 2786;
srom_1(33553) <= 7652;
srom_1(33554) <= 51820;
srom_1(33555) <= 135082;
srom_1(33556) <= 257048;
srom_1(33557) <= 417145;
srom_1(33558) <= 614623;
srom_1(33559) <= 848556;
srom_1(33560) <= 1117847;
srom_1(33561) <= 1421234;
srom_1(33562) <= 1757292;
srom_1(33563) <= 2124447;
srom_1(33564) <= 2520977;
srom_1(33565) <= 2945022;
srom_1(33566) <= 3394594;
srom_1(33567) <= 3867584;
srom_1(33568) <= 4361776;
srom_1(33569) <= 4874850;
srom_1(33570) <= 5404402;
srom_1(33571) <= 5947947;
srom_1(33572) <= 6502938;
srom_1(33573) <= 7066771;
srom_1(33574) <= 7636803;
srom_1(33575) <= 8210360;
srom_1(33576) <= 8784753;
srom_1(33577) <= 9357288;
srom_1(33578) <= 9925281;
srom_1(33579) <= 10486068;
srom_1(33580) <= 11037020;
srom_1(33581) <= 11575551;
srom_1(33582) <= 12099139;
srom_1(33583) <= 12605326;
srom_1(33584) <= 13091740;
srom_1(33585) <= 13556099;
srom_1(33586) <= 13996225;
srom_1(33587) <= 14410056;
srom_1(33588) <= 14795650;
srom_1(33589) <= 15151200;
srom_1(33590) <= 15475037;
srom_1(33591) <= 15765643;
srom_1(33592) <= 16021656;
srom_1(33593) <= 16241875;
srom_1(33594) <= 16425268;
srom_1(33595) <= 16570974;
srom_1(33596) <= 16678309;
srom_1(33597) <= 16746772;
srom_1(33598) <= 16776040;
srom_1(33599) <= 16765977;
srom_1(33600) <= 16716629;
srom_1(33601) <= 16628228;
srom_1(33602) <= 16501189;
srom_1(33603) <= 16336107;
srom_1(33604) <= 16133757;
srom_1(33605) <= 15895087;
srom_1(33606) <= 15621217;
srom_1(33607) <= 15313430;
srom_1(33608) <= 14973170;
srom_1(33609) <= 14602033;
srom_1(33610) <= 14201760;
srom_1(33611) <= 13774226;
srom_1(33612) <= 13321437;
srom_1(33613) <= 12845517;
srom_1(33614) <= 12348697;
srom_1(33615) <= 11833306;
srom_1(33616) <= 11301762;
srom_1(33617) <= 10756558;
srom_1(33618) <= 10200249;
srom_1(33619) <= 9635444;
srom_1(33620) <= 9064793;
srom_1(33621) <= 8490971;
srom_1(33622) <= 7916669;
srom_1(33623) <= 7344580;
srom_1(33624) <= 6777387;
srom_1(33625) <= 6217749;
srom_1(33626) <= 5668292;
srom_1(33627) <= 5131591;
srom_1(33628) <= 4610163;
srom_1(33629) <= 4106453;
srom_1(33630) <= 3622824;
srom_1(33631) <= 3161543;
srom_1(33632) <= 2724774;
srom_1(33633) <= 2314565;
srom_1(33634) <= 1932838;
srom_1(33635) <= 1581386;
srom_1(33636) <= 1261854;
srom_1(33637) <= 975742;
srom_1(33638) <= 724392;
srom_1(33639) <= 508982;
srom_1(33640) <= 330522;
srom_1(33641) <= 189849;
srom_1(33642) <= 87623;
srom_1(33643) <= 24324;
srom_1(33644) <= 247;
srom_1(33645) <= 15506;
srom_1(33646) <= 70029;
srom_1(33647) <= 163562;
srom_1(33648) <= 295664;
srom_1(33649) <= 465717;
srom_1(33650) <= 672922;
srom_1(33651) <= 916310;
srom_1(33652) <= 1194737;
srom_1(33653) <= 1506900;
srom_1(33654) <= 1851332;
srom_1(33655) <= 2226421;
srom_1(33656) <= 2630406;
srom_1(33657) <= 3061393;
srom_1(33658) <= 3517361;
srom_1(33659) <= 3996172;
srom_1(33660) <= 4495581;
srom_1(33661) <= 5013246;
srom_1(33662) <= 5546738;
srom_1(33663) <= 6093558;
srom_1(33664) <= 6651139;
srom_1(33665) <= 7216868;
srom_1(33666) <= 7788092;
srom_1(33667) <= 8362132;
srom_1(33668) <= 8936296;
srom_1(33669) <= 9507892;
srom_1(33670) <= 10074239;
srom_1(33671) <= 10632681;
srom_1(33672) <= 11180600;
srom_1(33673) <= 11715427;
srom_1(33674) <= 12234653;
srom_1(33675) <= 12735844;
srom_1(33676) <= 13216648;
srom_1(33677) <= 13674813;
srom_1(33678) <= 14108189;
srom_1(33679) <= 14514743;
srom_1(33680) <= 14892570;
srom_1(33681) <= 15239898;
srom_1(33682) <= 15555098;
srom_1(33683) <= 15836691;
srom_1(33684) <= 16083358;
srom_1(33685) <= 16293942;
srom_1(33686) <= 16467454;
srom_1(33687) <= 16603083;
srom_1(33688) <= 16700190;
srom_1(33689) <= 16758322;
srom_1(33690) <= 16777206;
srom_1(33691) <= 16756752;
srom_1(33692) <= 16697057;
srom_1(33693) <= 16598401;
srom_1(33694) <= 16461247;
srom_1(33695) <= 16286237;
srom_1(33696) <= 16074192;
srom_1(33697) <= 15826108;
srom_1(33698) <= 15543146;
srom_1(33699) <= 15226634;
srom_1(33700) <= 14878056;
srom_1(33701) <= 14499047;
srom_1(33702) <= 14091384;
srom_1(33703) <= 13656978;
srom_1(33704) <= 13197868;
srom_1(33705) <= 12716205;
srom_1(33706) <= 12214248;
srom_1(33707) <= 11694352;
srom_1(33708) <= 11158954;
srom_1(33709) <= 10610565;
srom_1(33710) <= 10051757;
srom_1(33711) <= 9485149;
srom_1(33712) <= 8913399;
srom_1(33713) <= 8339189;
srom_1(33714) <= 7765210;
srom_1(33715) <= 7194154;
srom_1(33716) <= 6628700;
srom_1(33717) <= 6071498;
srom_1(33718) <= 5525162;
srom_1(33719) <= 4992254;
srom_1(33720) <= 4475272;
srom_1(33721) <= 3976642;
srom_1(33722) <= 3498700;
srom_1(33723) <= 3043689;
srom_1(33724) <= 2613743;
srom_1(33725) <= 2210876;
srom_1(33726) <= 1836979;
srom_1(33727) <= 1493805;
srom_1(33728) <= 1182963;
srom_1(33729) <= 905911;
srom_1(33730) <= 663948;
srom_1(33731) <= 458208;
srom_1(33732) <= 289656;
srom_1(33733) <= 159084;
srom_1(33734) <= 67102;
srom_1(33735) <= 14143;
srom_1(33736) <= 454;
srom_1(33737) <= 26101;
srom_1(33738) <= 90962;
srom_1(33739) <= 194734;
srom_1(33740) <= 336929;
srom_1(33741) <= 516882;
srom_1(33742) <= 733748;
srom_1(33743) <= 986510;
srom_1(33744) <= 1273983;
srom_1(33745) <= 1594819;
srom_1(33746) <= 1947513;
srom_1(33747) <= 2330412;
srom_1(33748) <= 2741720;
srom_1(33749) <= 3179508;
srom_1(33750) <= 3641723;
srom_1(33751) <= 4126198;
srom_1(33752) <= 4630661;
srom_1(33753) <= 5152746;
srom_1(33754) <= 5690006;
srom_1(33755) <= 6239920;
srom_1(33756) <= 6799910;
srom_1(33757) <= 7367349;
srom_1(33758) <= 7939578;
srom_1(33759) <= 8513913;
srom_1(33760) <= 9087660;
srom_1(33761) <= 9658128;
srom_1(33762) <= 10222644;
srom_1(33763) <= 10778559;
srom_1(33764) <= 11323267;
srom_1(33765) <= 11854213;
srom_1(33766) <= 12368908;
srom_1(33767) <= 12864938;
srom_1(33768) <= 13339977;
srom_1(33769) <= 13791797;
srom_1(33770) <= 14218279;
srom_1(33771) <= 14617425;
srom_1(33772) <= 14987361;
srom_1(33773) <= 15326353;
srom_1(33774) <= 15632812;
srom_1(33775) <= 15905301;
srom_1(33776) <= 16142541;
srom_1(33777) <= 16343420;
srom_1(33778) <= 16506996;
srom_1(33779) <= 16632502;
srom_1(33780) <= 16719350;
srom_1(33781) <= 16767133;
srom_1(33782) <= 16775625;
srom_1(33783) <= 16744788;
srom_1(33784) <= 16674765;
srom_1(33785) <= 16565887;
srom_1(33786) <= 16418662;
srom_1(33787) <= 16233781;
srom_1(33788) <= 16012112;
srom_1(33789) <= 15754693;
srom_1(33790) <= 15462732;
srom_1(33791) <= 15137599;
srom_1(33792) <= 14780817;
srom_1(33793) <= 14394059;
srom_1(33794) <= 13979141;
srom_1(33795) <= 13538006;
srom_1(33796) <= 13072723;
srom_1(33797) <= 12585476;
srom_1(33798) <= 12078548;
srom_1(33799) <= 11554316;
srom_1(33800) <= 11015239;
srom_1(33801) <= 10463846;
srom_1(33802) <= 9902720;
srom_1(33803) <= 9334495;
srom_1(33804) <= 8761834;
srom_1(33805) <= 8187422;
srom_1(33806) <= 7613954;
srom_1(33807) <= 7044119;
srom_1(33808) <= 6480588;
srom_1(33809) <= 5926005;
srom_1(33810) <= 5382970;
srom_1(33811) <= 4854029;
srom_1(33812) <= 4341663;
srom_1(33813) <= 3848275;
srom_1(33814) <= 3376178;
srom_1(33815) <= 2927585;
srom_1(33816) <= 2504602;
srom_1(33817) <= 2109210;
srom_1(33818) <= 1743265;
srom_1(33819) <= 1408482;
srom_1(33820) <= 1106431;
srom_1(33821) <= 838529;
srom_1(33822) <= 606032;
srom_1(33823) <= 410030;
srom_1(33824) <= 251442;
srom_1(33825) <= 131012;
srom_1(33826) <= 49305;
srom_1(33827) <= 6704;
srom_1(33828) <= 3408;
srom_1(33829) <= 39434;
srom_1(33830) <= 114611;
srom_1(33831) <= 228588;
srom_1(33832) <= 380831;
srom_1(33833) <= 570624;
srom_1(33834) <= 797079;
srom_1(33835) <= 1059133;
srom_1(33836) <= 1355557;
srom_1(33837) <= 1684962;
srom_1(33838) <= 2045803;
srom_1(33839) <= 2436387;
srom_1(33840) <= 2854883;
srom_1(33841) <= 3299328;
srom_1(33842) <= 3767639;
srom_1(33843) <= 4257620;
srom_1(33844) <= 4766972;
srom_1(33845) <= 5293307;
srom_1(33846) <= 5834156;
srom_1(33847) <= 6386985;
srom_1(33848) <= 6949200;
srom_1(33849) <= 7518165;
srom_1(33850) <= 8091211;
srom_1(33851) <= 8665652;
srom_1(33852) <= 9238794;
srom_1(33853) <= 9807950;
srom_1(33854) <= 10370449;
srom_1(33855) <= 10923655;
srom_1(33856) <= 11464973;
srom_1(33857) <= 11991865;
srom_1(33858) <= 12501860;
srom_1(33859) <= 12992567;
srom_1(33860) <= 13461684;
srom_1(33861) <= 13907011;
srom_1(33862) <= 14326461;
srom_1(33863) <= 14718067;
srom_1(33864) <= 15079991;
srom_1(33865) <= 15410537;
srom_1(33866) <= 15708155;
srom_1(33867) <= 15971449;
srom_1(33868) <= 16199184;
srom_1(33869) <= 16390293;
srom_1(33870) <= 16543880;
srom_1(33871) <= 16659223;
srom_1(33872) <= 16735783;
srom_1(33873) <= 16773200;
srom_1(33874) <= 16771298;
srom_1(33875) <= 16730088;
srom_1(33876) <= 16649761;
srom_1(33877) <= 16530695;
srom_1(33878) <= 16373448;
srom_1(33879) <= 16178757;
srom_1(33880) <= 15947535;
srom_1(33881) <= 15680867;
srom_1(33882) <= 15380003;
srom_1(33883) <= 15046354;
srom_1(33884) <= 14681485;
srom_1(33885) <= 14287106;
srom_1(33886) <= 13865067;
srom_1(33887) <= 13417347;
srom_1(33888) <= 12946046;
srom_1(33889) <= 12453373;
srom_1(33890) <= 11941639;
srom_1(33891) <= 11413244;
srom_1(33892) <= 10870665;
srom_1(33893) <= 10316447;
srom_1(33894) <= 9753188;
srom_1(33895) <= 9183531;
srom_1(33896) <= 8610146;
srom_1(33897) <= 8035722;
srom_1(33898) <= 7462952;
srom_1(33899) <= 6894524;
srom_1(33900) <= 6333102;
srom_1(33901) <= 5781319;
srom_1(33902) <= 5241762;
srom_1(33903) <= 4716962;
srom_1(33904) <= 4209379;
srom_1(33905) <= 3721395;
srom_1(33906) <= 3255296;
srom_1(33907) <= 2813269;
srom_1(33908) <= 2397387;
srom_1(33909) <= 2009600;
srom_1(33910) <= 1651726;
srom_1(33911) <= 1325444;
srom_1(33912) <= 1032284;
srom_1(33913) <= 773619;
srom_1(33914) <= 550664;
srom_1(33915) <= 364464;
srom_1(33916) <= 215892;
srom_1(33917) <= 105644;
srom_1(33918) <= 34238;
srom_1(33919) <= 2009;
srom_1(33920) <= 9107;
srom_1(33921) <= 55500;
srom_1(33922) <= 140969;
srom_1(33923) <= 265115;
srom_1(33924) <= 427354;
srom_1(33925) <= 626926;
srom_1(33926) <= 862896;
srom_1(33927) <= 1134156;
srom_1(33928) <= 1439434;
srom_1(33929) <= 1777300;
srom_1(33930) <= 2146169;
srom_1(33931) <= 2544310;
srom_1(33932) <= 2969857;
srom_1(33933) <= 3420815;
srom_1(33934) <= 3895068;
srom_1(33935) <= 4390393;
srom_1(33936) <= 4904468;
srom_1(33937) <= 5434880;
srom_1(33938) <= 5979143;
srom_1(33939) <= 6534706;
srom_1(33940) <= 7098962;
srom_1(33941) <= 7669265;
srom_1(33942) <= 8242942;
srom_1(33943) <= 8817301;
srom_1(33944) <= 9389651;
srom_1(33945) <= 9957306;
srom_1(33946) <= 10517605;
srom_1(33947) <= 11067921;
srom_1(33948) <= 11605672;
srom_1(33949) <= 12128337;
srom_1(33950) <= 12633465;
srom_1(33951) <= 13118688;
srom_1(33952) <= 13581730;
srom_1(33953) <= 14020420;
srom_1(33954) <= 14432700;
srom_1(33955) <= 14816637;
srom_1(33956) <= 15170431;
srom_1(33957) <= 15492422;
srom_1(33958) <= 15781102;
srom_1(33959) <= 16035115;
srom_1(33960) <= 16253271;
srom_1(33961) <= 16434547;
srom_1(33962) <= 16578093;
srom_1(33963) <= 16683236;
srom_1(33964) <= 16749482;
srom_1(33965) <= 16776522;
srom_1(33966) <= 16764227;
srom_1(33967) <= 16712657;
srom_1(33968) <= 16622052;
srom_1(33969) <= 16492837;
srom_1(33970) <= 16325619;
srom_1(33971) <= 16121182;
srom_1(33972) <= 15880484;
srom_1(33973) <= 15604654;
srom_1(33974) <= 15294985;
srom_1(33975) <= 14952930;
srom_1(33976) <= 14580093;
srom_1(33977) <= 14178222;
srom_1(33978) <= 13749201;
srom_1(33979) <= 13295042;
srom_1(33980) <= 12817876;
srom_1(33981) <= 12319939;
srom_1(33982) <= 11803567;
srom_1(33983) <= 11271181;
srom_1(33984) <= 10725277;
srom_1(33985) <= 10168416;
srom_1(33986) <= 9603209;
srom_1(33987) <= 9032306;
srom_1(33988) <= 8458385;
srom_1(33989) <= 7884137;
srom_1(33990) <= 7312254;
srom_1(33991) <= 6745418;
srom_1(33992) <= 6186288;
srom_1(33993) <= 5637486;
srom_1(33994) <= 5101584;
srom_1(33995) <= 4581096;
srom_1(33996) <= 4078463;
srom_1(33997) <= 3596042;
srom_1(33998) <= 3136095;
srom_1(33999) <= 2700779;
srom_1(34000) <= 2292134;
srom_1(34001) <= 1912079;
srom_1(34002) <= 1562393;
srom_1(34003) <= 1244719;
srom_1(34004) <= 960544;
srom_1(34005) <= 711203;
srom_1(34006) <= 497863;
srom_1(34007) <= 321525;
srom_1(34008) <= 183017;
srom_1(34009) <= 82988;
srom_1(34010) <= 21907;
srom_1(34011) <= 60;
srom_1(34012) <= 17550;
srom_1(34013) <= 74294;
srom_1(34014) <= 170027;
srom_1(34015) <= 304300;
srom_1(34016) <= 476483;
srom_1(34017) <= 685769;
srom_1(34018) <= 931176;
srom_1(34019) <= 1211554;
srom_1(34020) <= 1525587;
srom_1(34021) <= 1871803;
srom_1(34022) <= 2248578;
srom_1(34023) <= 2654147;
srom_1(34024) <= 3086606;
srom_1(34025) <= 3543928;
srom_1(34026) <= 4023969;
srom_1(34027) <= 4524476;
srom_1(34028) <= 5043104;
srom_1(34029) <= 5577421;
srom_1(34030) <= 6124919;
srom_1(34031) <= 6683033;
srom_1(34032) <= 7249145;
srom_1(34033) <= 7820601;
srom_1(34034) <= 8394720;
srom_1(34035) <= 8968810;
srom_1(34036) <= 9540180;
srom_1(34037) <= 10106149;
srom_1(34038) <= 10664064;
srom_1(34039) <= 11211309;
srom_1(34040) <= 11745317;
srom_1(34041) <= 12263585;
srom_1(34042) <= 12763681;
srom_1(34043) <= 13243261;
srom_1(34044) <= 13700076;
srom_1(34045) <= 14131984;
srom_1(34046) <= 14536959;
srom_1(34047) <= 14913102;
srom_1(34048) <= 15258650;
srom_1(34049) <= 15571981;
srom_1(34050) <= 15851628;
srom_1(34051) <= 16096277;
srom_1(34052) <= 16304783;
srom_1(34053) <= 16476167;
srom_1(34054) <= 16609626;
srom_1(34055) <= 16704534;
srom_1(34056) <= 16760445;
srom_1(34057) <= 16777098;
srom_1(34058) <= 16754414;
srom_1(34059) <= 16692500;
srom_1(34060) <= 16591647;
srom_1(34061) <= 16452326;
srom_1(34062) <= 16275192;
srom_1(34063) <= 16061075;
srom_1(34064) <= 15810980;
srom_1(34065) <= 15526078;
srom_1(34066) <= 15207706;
srom_1(34067) <= 14857357;
srom_1(34068) <= 14476674;
srom_1(34069) <= 14067442;
srom_1(34070) <= 13631579;
srom_1(34071) <= 13171131;
srom_1(34072) <= 12688256;
srom_1(34073) <= 12185218;
srom_1(34074) <= 11664377;
srom_1(34075) <= 11128174;
srom_1(34076) <= 10579125;
srom_1(34077) <= 10019803;
srom_1(34078) <= 9452833;
srom_1(34079) <= 8880871;
srom_1(34080) <= 8306602;
srom_1(34081) <= 7732717;
srom_1(34082) <= 7161907;
srom_1(34083) <= 6596850;
srom_1(34084) <= 6040196;
srom_1(34085) <= 5494553;
srom_1(34086) <= 4962482;
srom_1(34087) <= 4446477;
srom_1(34088) <= 3948959;
srom_1(34089) <= 3472259;
srom_1(34090) <= 3018613;
srom_1(34091) <= 2590150;
srom_1(34092) <= 2188877;
srom_1(34093) <= 1816677;
srom_1(34094) <= 1475295;
srom_1(34095) <= 1166332;
srom_1(34096) <= 891237;
srom_1(34097) <= 651299;
srom_1(34098) <= 447645;
srom_1(34099) <= 281228;
srom_1(34100) <= 152829;
srom_1(34101) <= 63051;
srom_1(34102) <= 12315;
srom_1(34103) <= 857;
srom_1(34104) <= 28733;
srom_1(34105) <= 95811;
srom_1(34106) <= 201776;
srom_1(34107) <= 346133;
srom_1(34108) <= 528203;
srom_1(34109) <= 747134;
srom_1(34110) <= 1001898;
srom_1(34111) <= 1291301;
srom_1(34112) <= 1613986;
srom_1(34113) <= 1968439;
srom_1(34114) <= 2352998;
srom_1(34115) <= 2765861;
srom_1(34116) <= 3205090;
srom_1(34117) <= 3668627;
srom_1(34118) <= 4154298;
srom_1(34119) <= 4659824;
srom_1(34120) <= 5182836;
srom_1(34121) <= 5720881;
srom_1(34122) <= 6271436;
srom_1(34123) <= 6831920;
srom_1(34124) <= 7399702;
srom_1(34125) <= 7972123;
srom_1(34126) <= 8546496;
srom_1(34127) <= 9120129;
srom_1(34128) <= 9690331;
srom_1(34129) <= 10254430;
srom_1(34130) <= 10809778;
srom_1(34131) <= 11353773;
srom_1(34132) <= 11883864;
srom_1(34133) <= 12397564;
srom_1(34134) <= 12892464;
srom_1(34135) <= 13366245;
srom_1(34136) <= 13816683;
srom_1(34137) <= 14241668;
srom_1(34138) <= 14639205;
srom_1(34139) <= 15007431;
srom_1(34140) <= 15344620;
srom_1(34141) <= 15649189;
srom_1(34142) <= 15919711;
srom_1(34143) <= 16154916;
srom_1(34144) <= 16353703;
srom_1(34145) <= 16515139;
srom_1(34146) <= 16638467;
srom_1(34147) <= 16723108;
srom_1(34148) <= 16768666;
srom_1(34149) <= 16774927;
srom_1(34150) <= 16741862;
srom_1(34151) <= 16669626;
srom_1(34152) <= 16558556;
srom_1(34153) <= 16409176;
srom_1(34154) <= 16222183;
srom_1(34155) <= 15998457;
srom_1(34156) <= 15739045;
srom_1(34157) <= 15445165;
srom_1(34158) <= 15118194;
srom_1(34159) <= 14759666;
srom_1(34160) <= 14371261;
srom_1(34161) <= 13954802;
srom_1(34162) <= 13512241;
srom_1(34163) <= 13045654;
srom_1(34164) <= 12557228;
srom_1(34165) <= 12049254;
srom_1(34166) <= 11524114;
srom_1(34167) <= 10984271;
srom_1(34168) <= 10432255;
srom_1(34169) <= 9870656;
srom_1(34170) <= 9302108;
srom_1(34171) <= 8729275;
srom_1(34172) <= 8154845;
srom_1(34173) <= 7581512;
srom_1(34174) <= 7011963;
srom_1(34175) <= 6448869;
srom_1(34176) <= 5894872;
srom_1(34177) <= 5352568;
srom_1(34178) <= 4824502;
srom_1(34179) <= 4313149;
srom_1(34180) <= 3820907;
srom_1(34181) <= 3350085;
srom_1(34182) <= 2902890;
srom_1(34183) <= 2481420;
srom_1(34184) <= 2087650;
srom_1(34185) <= 1723428;
srom_1(34186) <= 1390461;
srom_1(34187) <= 1090310;
srom_1(34188) <= 824384;
srom_1(34189) <= 593929;
srom_1(34190) <= 400026;
srom_1(34191) <= 243585;
srom_1(34192) <= 125338;
srom_1(34193) <= 45840;
srom_1(34194) <= 5465;
srom_1(34195) <= 4400;
srom_1(34196) <= 42653;
srom_1(34197) <= 120042;
srom_1(34198) <= 236206;
srom_1(34199) <= 390599;
srom_1(34200) <= 582497;
srom_1(34201) <= 811001;
srom_1(34202) <= 1075039;
srom_1(34203) <= 1373372;
srom_1(34204) <= 1704603;
srom_1(34205) <= 2067177;
srom_1(34206) <= 2459394;
srom_1(34207) <= 2879416;
srom_1(34208) <= 3325272;
srom_1(34209) <= 3794872;
srom_1(34210) <= 4286013;
srom_1(34211) <= 4796393;
srom_1(34212) <= 5323618;
srom_1(34213) <= 5865216;
srom_1(34214) <= 6418647;
srom_1(34215) <= 6981315;
srom_1(34216) <= 7550583;
srom_1(34217) <= 8123781;
srom_1(34218) <= 8698220;
srom_1(34219) <= 9271208;
srom_1(34220) <= 9840057;
srom_1(34221) <= 10402099;
srom_1(34222) <= 10954700;
srom_1(34223) <= 11495267;
srom_1(34224) <= 12021266;
srom_1(34225) <= 12530230;
srom_1(34226) <= 13019773;
srom_1(34227) <= 13487599;
srom_1(34228) <= 13931513;
srom_1(34229) <= 14349435;
srom_1(34230) <= 14739405;
srom_1(34231) <= 15099594;
srom_1(34232) <= 15428312;
srom_1(34233) <= 15724019;
srom_1(34234) <= 15985328;
srom_1(34235) <= 16211013;
srom_1(34236) <= 16400016;
srom_1(34237) <= 16551451;
srom_1(34238) <= 16664607;
srom_1(34239) <= 16738955;
srom_1(34240) <= 16774144;
srom_1(34241) <= 16770011;
srom_1(34242) <= 16726575;
srom_1(34243) <= 16644040;
srom_1(34244) <= 16522791;
srom_1(34245) <= 16363399;
srom_1(34246) <= 16166610;
srom_1(34247) <= 15933347;
srom_1(34248) <= 15664705;
srom_1(34249) <= 15361942;
srom_1(34250) <= 15026479;
srom_1(34251) <= 14659889;
srom_1(34252) <= 14263891;
srom_1(34253) <= 13840341;
srom_1(34254) <= 13391226;
srom_1(34255) <= 12918652;
srom_1(34256) <= 12424836;
srom_1(34257) <= 11912092;
srom_1(34258) <= 11382825;
srom_1(34259) <= 10839517;
srom_1(34260) <= 10284716;
srom_1(34261) <= 9721024;
srom_1(34262) <= 9151084;
srom_1(34263) <= 8577568;
srom_1(34264) <= 8003165;
srom_1(34265) <= 7430571;
srom_1(34266) <= 6862469;
srom_1(34267) <= 6301523;
srom_1(34268) <= 5750365;
srom_1(34269) <= 5211578;
srom_1(34270) <= 4687689;
srom_1(34271) <= 4181155;
srom_1(34272) <= 3694352;
srom_1(34273) <= 3229561;
srom_1(34274) <= 2788963;
srom_1(34275) <= 2374623;
srom_1(34276) <= 1988485;
srom_1(34277) <= 1632360;
srom_1(34278) <= 1307917;
srom_1(34279) <= 1016678;
srom_1(34280) <= 760008;
srom_1(34281) <= 539111;
srom_1(34282) <= 355023;
srom_1(34283) <= 208608;
srom_1(34284) <= 100551;
srom_1(34285) <= 31360;
srom_1(34286) <= 1359;
srom_1(34287) <= 10689;
srom_1(34288) <= 59305;
srom_1(34289) <= 146981;
srom_1(34290) <= 273304;
srom_1(34291) <= 437683;
srom_1(34292) <= 639346;
srom_1(34293) <= 877348;
srom_1(34294) <= 1150573;
srom_1(34295) <= 1457740;
srom_1(34296) <= 1797408;
srom_1(34297) <= 2167984;
srom_1(34298) <= 2567732;
srom_1(34299) <= 2994775;
srom_1(34300) <= 3447111;
srom_1(34301) <= 3922620;
srom_1(34302) <= 4419072;
srom_1(34303) <= 4934138;
srom_1(34304) <= 5465403;
srom_1(34305) <= 6010376;
srom_1(34306) <= 6566502;
srom_1(34307) <= 7131172;
srom_1(34308) <= 7701738;
srom_1(34309) <= 8275526;
srom_1(34310) <= 8849843;
srom_1(34311) <= 9421998;
srom_1(34312) <= 9989307;
srom_1(34313) <= 10549110;
srom_1(34314) <= 11098781;
srom_1(34315) <= 11635744;
srom_1(34316) <= 12157479;
srom_1(34317) <= 12661541;
srom_1(34318) <= 13145566;
srom_1(34319) <= 13607283;
srom_1(34320) <= 14044529;
srom_1(34321) <= 14455252;
srom_1(34322) <= 14837526;
srom_1(34323) <= 15189559;
srom_1(34324) <= 15509700;
srom_1(34325) <= 15796448;
srom_1(34326) <= 16048458;
srom_1(34327) <= 16264548;
srom_1(34328) <= 16443706;
srom_1(34329) <= 16585090;
srom_1(34330) <= 16688038;
srom_1(34331) <= 16752067;
srom_1(34332) <= 16776877;
srom_1(34333) <= 16762352;
srom_1(34334) <= 16708559;
srom_1(34335) <= 16615751;
srom_1(34336) <= 16484363;
srom_1(34337) <= 16315011;
srom_1(34338) <= 16108490;
srom_1(34339) <= 15865767;
srom_1(34340) <= 15587982;
srom_1(34341) <= 15276436;
srom_1(34342) <= 14932591;
srom_1(34343) <= 14558059;
srom_1(34344) <= 14154596;
srom_1(34345) <= 13724094;
srom_1(34346) <= 13268573;
srom_1(34347) <= 12790168;
srom_1(34348) <= 12291122;
srom_1(34349) <= 11773776;
srom_1(34350) <= 11240556;
srom_1(34351) <= 10693962;
srom_1(34352) <= 10136557;
srom_1(34353) <= 9570956;
srom_1(34354) <= 8999810;
srom_1(34355) <= 8425798;
srom_1(34356) <= 7851612;
srom_1(34357) <= 7279943;
srom_1(34358) <= 6713474;
srom_1(34359) <= 6154860;
srom_1(34360) <= 5606721;
srom_1(34361) <= 5071627;
srom_1(34362) <= 4552087;
srom_1(34363) <= 4050539;
srom_1(34364) <= 3569333;
srom_1(34365) <= 3110726;
srom_1(34366) <= 2676869;
srom_1(34367) <= 2269796;
srom_1(34368) <= 1891416;
srom_1(34369) <= 1543504;
srom_1(34370) <= 1227691;
srom_1(34371) <= 945458;
srom_1(34372) <= 698129;
srom_1(34373) <= 486863;
srom_1(34374) <= 312651;
srom_1(34375) <= 176309;
srom_1(34376) <= 78478;
srom_1(34377) <= 19616;
srom_1(34378) <= 0;
srom_1(34379) <= 19720;
srom_1(34380) <= 78684;
srom_1(34381) <= 176617;
srom_1(34382) <= 313059;
srom_1(34383) <= 487370;
srom_1(34384) <= 698732;
srom_1(34385) <= 946155;
srom_1(34386) <= 1228478;
srom_1(34387) <= 1544377;
srom_1(34388) <= 1892371;
srom_1(34389) <= 2270829;
srom_1(34390) <= 2677974;
srom_1(34391) <= 3111899;
srom_1(34392) <= 3570568;
srom_1(34393) <= 4051831;
srom_1(34394) <= 4553430;
srom_1(34395) <= 5073014;
srom_1(34396) <= 5608145;
srom_1(34397) <= 6156315;
srom_1(34398) <= 6714953;
srom_1(34399) <= 7281440;
srom_1(34400) <= 7853118;
srom_1(34401) <= 8427308;
srom_1(34402) <= 9001315;
srom_1(34403) <= 9572450;
srom_1(34404) <= 10138033;
srom_1(34405) <= 10695413;
srom_1(34406) <= 11241975;
srom_1(34407) <= 11775157;
srom_1(34408) <= 12292458;
srom_1(34409) <= 12791453;
srom_1(34410) <= 13269801;
srom_1(34411) <= 13725259;
srom_1(34412) <= 14155692;
srom_1(34413) <= 14559082;
srom_1(34414) <= 14933535;
srom_1(34415) <= 15277298;
srom_1(34416) <= 15588757;
srom_1(34417) <= 15866452;
srom_1(34418) <= 16109080;
srom_1(34419) <= 16315505;
srom_1(34420) <= 16484758;
srom_1(34421) <= 16616045;
srom_1(34422) <= 16708751;
srom_1(34423) <= 16762441;
srom_1(34424) <= 16776863;
srom_1(34425) <= 16751950;
srom_1(34426) <= 16687818;
srom_1(34427) <= 16584768;
srom_1(34428) <= 16443284;
srom_1(34429) <= 16264029;
srom_1(34430) <= 16047843;
srom_1(34431) <= 15795740;
srom_1(34432) <= 15508902;
srom_1(34433) <= 15188675;
srom_1(34434) <= 14836560;
srom_1(34435) <= 14454209;
srom_1(34436) <= 14043414;
srom_1(34437) <= 13606101;
srom_1(34438) <= 13144322;
srom_1(34439) <= 12660242;
srom_1(34440) <= 12156130;
srom_1(34441) <= 11634352;
srom_1(34442) <= 11097352;
srom_1(34443) <= 10547651;
srom_1(34444) <= 9987825;
srom_1(34445) <= 9420500;
srom_1(34446) <= 8848336;
srom_1(34447) <= 8274016;
srom_1(34448) <= 7700234;
srom_1(34449) <= 7129679;
srom_1(34450) <= 6565028;
srom_1(34451) <= 6008929;
srom_1(34452) <= 5463988;
srom_1(34453) <= 4932762;
srom_1(34454) <= 4417742;
srom_1(34455) <= 3921342;
srom_1(34456) <= 3445891;
srom_1(34457) <= 2993619;
srom_1(34458) <= 2566645;
srom_1(34459) <= 2166972;
srom_1(34460) <= 1796474;
srom_1(34461) <= 1456890;
srom_1(34462) <= 1149810;
srom_1(34463) <= 876676;
srom_1(34464) <= 638768;
srom_1(34465) <= 437201;
srom_1(34466) <= 272922;
srom_1(34467) <= 146699;
srom_1(34468) <= 59126;
srom_1(34469) <= 10613;
srom_1(34470) <= 1386;
srom_1(34471) <= 31491;
srom_1(34472) <= 100784;
srom_1(34473) <= 208943;
srom_1(34474) <= 355458;
srom_1(34475) <= 539644;
srom_1(34476) <= 760636;
srom_1(34477) <= 1017398;
srom_1(34478) <= 1308726;
srom_1(34479) <= 1633255;
srom_1(34480) <= 1989461;
srom_1(34481) <= 2375676;
srom_1(34482) <= 2790087;
srom_1(34483) <= 3230751;
srom_1(34484) <= 3695603;
srom_1(34485) <= 4182461;
srom_1(34486) <= 4689044;
srom_1(34487) <= 5212975;
srom_1(34488) <= 5751798;
srom_1(34489) <= 6302985;
srom_1(34490) <= 6863953;
srom_1(34491) <= 7432070;
srom_1(34492) <= 8004673;
srom_1(34493) <= 8579077;
srom_1(34494) <= 9152587;
srom_1(34495) <= 9722514;
srom_1(34496) <= 10286187;
srom_1(34497) <= 10840961;
srom_1(34498) <= 11384235;
srom_1(34499) <= 11913462;
srom_1(34500) <= 12426159;
srom_1(34501) <= 12919923;
srom_1(34502) <= 13392438;
srom_1(34503) <= 13841488;
srom_1(34504) <= 14264968;
srom_1(34505) <= 14660891;
srom_1(34506) <= 15027402;
srom_1(34507) <= 15362781;
srom_1(34508) <= 15665456;
srom_1(34509) <= 15934007;
srom_1(34510) <= 16167175;
srom_1(34511) <= 16363867;
srom_1(34512) <= 16523160;
srom_1(34513) <= 16644307;
srom_1(34514) <= 16726741;
srom_1(34515) <= 16770074;
srom_1(34516) <= 16774103;
srom_1(34517) <= 16738810;
srom_1(34518) <= 16664361;
srom_1(34519) <= 16551103;
srom_1(34520) <= 16399568;
srom_1(34521) <= 16210468;
srom_1(34522) <= 15984688;
srom_1(34523) <= 15723287;
srom_1(34524) <= 15427491;
srom_1(34525) <= 15098688;
srom_1(34526) <= 14738419;
srom_1(34527) <= 14348373;
srom_1(34528) <= 13930380;
srom_1(34529) <= 13486400;
srom_1(34530) <= 13018514;
srom_1(34531) <= 12528918;
srom_1(34532) <= 12019905;
srom_1(34533) <= 11493865;
srom_1(34534) <= 10953263;
srom_1(34535) <= 10400634;
srom_1(34536) <= 9838570;
srom_1(34537) <= 9269707;
srom_1(34538) <= 8696712;
srom_1(34539) <= 8122272;
srom_1(34540) <= 7549081;
srom_1(34541) <= 6979827;
srom_1(34542) <= 6417179;
srom_1(34543) <= 5863776;
srom_1(34544) <= 5322213;
srom_1(34545) <= 4795029;
srom_1(34546) <= 4284697;
srom_1(34547) <= 3793609;
srom_1(34548) <= 3324069;
srom_1(34549) <= 2878278;
srom_1(34550) <= 2458327;
srom_1(34551) <= 2066185;
srom_1(34552) <= 1703691;
srom_1(34553) <= 1372545;
srom_1(34554) <= 1074299;
srom_1(34555) <= 810353;
srom_1(34556) <= 581944;
srom_1(34557) <= 390143;
srom_1(34558) <= 235850;
srom_1(34559) <= 119788;
srom_1(34560) <= 42501;
srom_1(34561) <= 4352;
srom_1(34562) <= 5519;
srom_1(34563) <= 45998;
srom_1(34564) <= 125598;
srom_1(34565) <= 243946;
srom_1(34566) <= 400487;
srom_1(34567) <= 594487;
srom_1(34568) <= 825037;
srom_1(34569) <= 1091055;
srom_1(34570) <= 1391293;
srom_1(34571) <= 1724344;
srom_1(34572) <= 2088647;
srom_1(34573) <= 2482492;
srom_1(34574) <= 2904032;
srom_1(34575) <= 3351292;
srom_1(34576) <= 3822174;
srom_1(34577) <= 4314469;
srom_1(34578) <= 4825869;
srom_1(34579) <= 5353976;
srom_1(34580) <= 5896313;
srom_1(34581) <= 6450338;
srom_1(34582) <= 7013452;
srom_1(34583) <= 7583014;
srom_1(34584) <= 8156354;
srom_1(34585) <= 8730784;
srom_1(34586) <= 9303608;
srom_1(34587) <= 9872142;
srom_1(34588) <= 10433719;
srom_1(34589) <= 10985706;
srom_1(34590) <= 11525514;
srom_1(34591) <= 12050612;
srom_1(34592) <= 12558538;
srom_1(34593) <= 13046910;
srom_1(34594) <= 13513437;
srom_1(34595) <= 13955932;
srom_1(34596) <= 14372320;
srom_1(34597) <= 14760648;
srom_1(34598) <= 15119095;
srom_1(34599) <= 15445981;
srom_1(34600) <= 15739773;
srom_1(34601) <= 15999092;
srom_1(34602) <= 16222723;
srom_1(34603) <= 16409618;
srom_1(34604) <= 16558899;
srom_1(34605) <= 16669866;
srom_1(34606) <= 16742000;
srom_1(34607) <= 16774963;
srom_1(34608) <= 16768598;
srom_1(34609) <= 16722937;
srom_1(34610) <= 16638194;
srom_1(34611) <= 16514765;
srom_1(34612) <= 16353230;
srom_1(34613) <= 16154346;
srom_1(34614) <= 15919046;
srom_1(34615) <= 15648433;
srom_1(34616) <= 15343776;
srom_1(34617) <= 15006504;
srom_1(34618) <= 14638198;
srom_1(34619) <= 14240586;
srom_1(34620) <= 13815532;
srom_1(34621) <= 13365030;
srom_1(34622) <= 12891191;
srom_1(34623) <= 12396238;
srom_1(34624) <= 11882491;
srom_1(34625) <= 11352361;
srom_1(34626) <= 10808333;
srom_1(34627) <= 10252958;
srom_1(34628) <= 9688840;
srom_1(34629) <= 9118625;
srom_1(34630) <= 8544987;
srom_1(34631) <= 7970615;
srom_1(34632) <= 7398203;
srom_1(34633) <= 6830436;
srom_1(34634) <= 6269976;
srom_1(34635) <= 5719450;
srom_1(34636) <= 5181441;
srom_1(34637) <= 4658472;
srom_1(34638) <= 4152995;
srom_1(34639) <= 3667379;
srom_1(34640) <= 3203904;
srom_1(34641) <= 2764741;
srom_1(34642) <= 2351950;
srom_1(34643) <= 1967467;
srom_1(34644) <= 1613096;
srom_1(34645) <= 1290496;
srom_1(34646) <= 1001183;
srom_1(34647) <= 746511;
srom_1(34648) <= 527676;
srom_1(34649) <= 345704;
srom_1(34650) <= 201447;
srom_1(34651) <= 95583;
srom_1(34652) <= 28608;
srom_1(34653) <= 836;
srom_1(34654) <= 12396;
srom_1(34655) <= 63236;
srom_1(34656) <= 153116;
srom_1(34657) <= 281616;
srom_1(34658) <= 448131;
srom_1(34659) <= 651883;
srom_1(34660) <= 891914;
srom_1(34661) <= 1167100;
srom_1(34662) <= 1476150;
srom_1(34663) <= 1817616;
srom_1(34664) <= 2189894;
srom_1(34665) <= 2591241;
srom_1(34666) <= 3019773;
srom_1(34667) <= 3473482;
srom_1(34668) <= 3950239;
srom_1(34669) <= 4447810;
srom_1(34670) <= 4963860;
srom_1(34671) <= 5495970;
srom_1(34672) <= 6041645;
srom_1(34673) <= 6598325;
srom_1(34674) <= 7163401;
srom_1(34675) <= 7734222;
srom_1(34676) <= 8308111;
srom_1(34677) <= 8882378;
srom_1(34678) <= 9454330;
srom_1(34679) <= 10021284;
srom_1(34680) <= 10580582;
srom_1(34681) <= 11129601;
srom_1(34682) <= 11665766;
srom_1(34683) <= 12186564;
srom_1(34684) <= 12689552;
srom_1(34685) <= 13172371;
srom_1(34686) <= 13632758;
srom_1(34687) <= 14068553;
srom_1(34688) <= 14477712;
srom_1(34689) <= 14858318;
srom_1(34690) <= 15208585;
srom_1(34691) <= 15526871;
srom_1(34692) <= 15811683;
srom_1(34693) <= 16061686;
srom_1(34694) <= 16275707;
srom_1(34695) <= 16452742;
srom_1(34696) <= 16591962;
srom_1(34697) <= 16692714;
srom_1(34698) <= 16754525;
srom_1(34699) <= 16777106;
srom_1(34700) <= 16760349;
srom_1(34701) <= 16704335;
srom_1(34702) <= 16609326;
srom_1(34703) <= 16475766;
srom_1(34704) <= 16304284;
srom_1(34705) <= 16095682;
srom_1(34706) <= 15850938;
srom_1(34707) <= 15571202;
srom_1(34708) <= 15257783;
srom_1(34709) <= 14912153;
srom_1(34710) <= 14535932;
srom_1(34711) <= 14130883;
srom_1(34712) <= 13698908;
srom_1(34713) <= 13242030;
srom_1(34714) <= 12762393;
srom_1(34715) <= 12262246;
srom_1(34716) <= 11743934;
srom_1(34717) <= 11209887;
srom_1(34718) <= 10662611;
srom_1(34719) <= 10104671;
srom_1(34720) <= 9538684;
srom_1(34721) <= 8967304;
srom_1(34722) <= 8393210;
srom_1(34723) <= 7819095;
srom_1(34724) <= 7247650;
srom_1(34725) <= 6681555;
srom_1(34726) <= 6123466;
srom_1(34727) <= 5575998;
srom_1(34728) <= 5041720;
srom_1(34729) <= 4523137;
srom_1(34730) <= 4022679;
srom_1(34731) <= 3542696;
srom_1(34732) <= 3085436;
srom_1(34733) <= 2653045;
srom_1(34734) <= 2247550;
srom_1(34735) <= 1870852;
srom_1(34736) <= 1524719;
srom_1(34737) <= 1210772;
srom_1(34738) <= 930485;
srom_1(34739) <= 685171;
srom_1(34740) <= 475982;
srom_1(34741) <= 303898;
srom_1(34742) <= 169725;
srom_1(34743) <= 74094;
srom_1(34744) <= 17452;
srom_1(34745) <= 66;
srom_1(34746) <= 22016;
srom_1(34747) <= 83200;
srom_1(34748) <= 183331;
srom_1(34749) <= 321940;
srom_1(34750) <= 498375;
srom_1(34751) <= 711811;
srom_1(34752) <= 961246;
srom_1(34753) <= 1245510;
srom_1(34754) <= 1563271;
srom_1(34755) <= 1913038;
srom_1(34756) <= 2293171;
srom_1(34757) <= 2701888;
srom_1(34758) <= 3137272;
srom_1(34759) <= 3597281;
srom_1(34760) <= 4079758;
srom_1(34761) <= 4582441;
srom_1(34762) <= 5102973;
srom_1(34763) <= 5638912;
srom_1(34764) <= 6187745;
srom_1(34765) <= 6746899;
srom_1(34766) <= 7313751;
srom_1(34767) <= 7885643;
srom_1(34768) <= 8459895;
srom_1(34769) <= 9033812;
srom_1(34770) <= 9604703;
srom_1(34771) <= 10169891;
srom_1(34772) <= 10726727;
srom_1(34773) <= 11272598;
srom_1(34774) <= 11804946;
srom_1(34775) <= 12321272;
srom_1(34776) <= 12819158;
srom_1(34777) <= 13296267;
srom_1(34778) <= 13750362;
srom_1(34779) <= 14179314;
srom_1(34780) <= 14581111;
srom_1(34781) <= 14953870;
srom_1(34782) <= 15295842;
srom_1(34783) <= 15605423;
srom_1(34784) <= 15881163;
srom_1(34785) <= 16121767;
srom_1(34786) <= 16326108;
srom_1(34787) <= 16493227;
srom_1(34788) <= 16622340;
srom_1(34789) <= 16712843;
srom_1(34790) <= 16764311;
srom_1(34791) <= 16776502;
srom_1(34792) <= 16749360;
srom_1(34793) <= 16683011;
srom_1(34794) <= 16577766;
srom_1(34795) <= 16434120;
srom_1(34796) <= 16252746;
srom_1(34797) <= 16034494;
srom_1(34798) <= 15780388;
srom_1(34799) <= 15491619;
srom_1(34800) <= 15169542;
srom_1(34801) <= 14815667;
srom_1(34802) <= 14431653;
srom_1(34803) <= 14019301;
srom_1(34804) <= 13580544;
srom_1(34805) <= 13117441;
srom_1(34806) <= 12632163;
srom_1(34807) <= 12126986;
srom_1(34808) <= 11604278;
srom_1(34809) <= 11066490;
srom_1(34810) <= 10516145;
srom_1(34811) <= 9955823;
srom_1(34812) <= 9388152;
srom_1(34813) <= 8815794;
srom_1(34814) <= 8241432;
srom_1(34815) <= 7667761;
srom_1(34816) <= 7097470;
srom_1(34817) <= 6533234;
srom_1(34818) <= 5977698;
srom_1(34819) <= 5433467;
srom_1(34820) <= 4903094;
srom_1(34821) <= 4389066;
srom_1(34822) <= 3893794;
srom_1(34823) <= 3419599;
srom_1(34824) <= 2968705;
srom_1(34825) <= 2543227;
srom_1(34826) <= 2145160;
srom_1(34827) <= 1776371;
srom_1(34828) <= 1438589;
srom_1(34829) <= 1133398;
srom_1(34830) <= 862229;
srom_1(34831) <= 626354;
srom_1(34832) <= 426878;
srom_1(34833) <= 264738;
srom_1(34834) <= 140694;
srom_1(34835) <= 55327;
srom_1(34836) <= 9037;
srom_1(34837) <= 2042;
srom_1(34838) <= 34375;
srom_1(34839) <= 105883;
srom_1(34840) <= 216232;
srom_1(34841) <= 364904;
srom_1(34842) <= 551202;
srom_1(34843) <= 774253;
srom_1(34844) <= 1033009;
srom_1(34845) <= 1326259;
srom_1(34846) <= 1652626;
srom_1(34847) <= 2010581;
srom_1(34848) <= 2398444;
srom_1(34849) <= 2814397;
srom_1(34850) <= 3256490;
srom_1(34851) <= 3722649;
srom_1(34852) <= 4210688;
srom_1(34853) <= 4718319;
srom_1(34854) <= 5243161;
srom_1(34855) <= 5782753;
srom_1(34856) <= 6334565;
srom_1(34857) <= 6896009;
srom_1(34858) <= 7464453;
srom_1(34859) <= 8037230;
srom_1(34860) <= 8611655;
srom_1(34861) <= 9185033;
srom_1(34862) <= 9754678;
srom_1(34863) <= 10317916;
srom_1(34864) <= 10872107;
srom_1(34865) <= 11414652;
srom_1(34866) <= 11943006;
srom_1(34867) <= 12454693;
srom_1(34868) <= 12947313;
srom_1(34869) <= 13418555;
srom_1(34870) <= 13866211;
srom_1(34871) <= 14288179;
srom_1(34872) <= 14682483;
srom_1(34873) <= 15047273;
srom_1(34874) <= 15380837;
srom_1(34875) <= 15681613;
srom_1(34876) <= 15948190;
srom_1(34877) <= 16179317;
srom_1(34878) <= 16373910;
srom_1(34879) <= 16531058;
srom_1(34880) <= 16650023;
srom_1(34881) <= 16730247;
srom_1(34882) <= 16771355;
srom_1(34883) <= 16773153;
srom_1(34884) <= 16735633;
srom_1(34885) <= 16658971;
srom_1(34886) <= 16543526;
srom_1(34887) <= 16389840;
srom_1(34888) <= 16198634;
srom_1(34889) <= 15970803;
srom_1(34890) <= 15707417;
srom_1(34891) <= 15409711;
srom_1(34892) <= 15079081;
srom_1(34893) <= 14717076;
srom_1(34894) <= 14325395;
srom_1(34895) <= 13905874;
srom_1(34896) <= 13460481;
srom_1(34897) <= 12991305;
srom_1(34898) <= 12500544;
srom_1(34899) <= 11990502;
srom_1(34900) <= 11463569;
srom_1(34901) <= 10922216;
srom_1(34902) <= 10368982;
srom_1(34903) <= 9806462;
srom_1(34904) <= 9237293;
srom_1(34905) <= 8664144;
srom_1(34906) <= 8089703;
srom_1(34907) <= 7516663;
srom_1(34908) <= 6947713;
srom_1(34909) <= 6385519;
srom_1(34910) <= 5832719;
srom_1(34911) <= 5291903;
srom_1(34912) <= 4765610;
srom_1(34913) <= 4256306;
srom_1(34914) <= 3766379;
srom_1(34915) <= 3298128;
srom_1(34916) <= 2853748;
srom_1(34917) <= 2435323;
srom_1(34918) <= 2044815;
srom_1(34919) <= 1684055;
srom_1(34920) <= 1354735;
srom_1(34921) <= 1058399;
srom_1(34922) <= 796437;
srom_1(34923) <= 570077;
srom_1(34924) <= 380381;
srom_1(34925) <= 228238;
srom_1(34926) <= 114363;
srom_1(34927) <= 39288;
srom_1(34928) <= 3365;
srom_1(34929) <= 6764;
srom_1(34930) <= 49469;
srom_1(34931) <= 131278;
srom_1(34932) <= 251809;
srom_1(34933) <= 410496;
srom_1(34934) <= 606595;
srom_1(34935) <= 839187;
srom_1(34936) <= 1107181;
srom_1(34937) <= 1409319;
srom_1(34938) <= 1744186;
srom_1(34939) <= 2110211;
srom_1(34940) <= 2505678;
srom_1(34941) <= 2928731;
srom_1(34942) <= 3377388;
srom_1(34943) <= 3849544;
srom_1(34944) <= 4342986;
srom_1(34945) <= 4855398;
srom_1(34946) <= 5384379;
srom_1(34947) <= 5927448;
srom_1(34948) <= 6482058;
srom_1(34949) <= 7045609;
srom_1(34950) <= 7615457;
srom_1(34951) <= 8188931;
srom_1(34952) <= 8763342;
srom_1(34953) <= 9335995;
srom_1(34954) <= 9904205;
srom_1(34955) <= 10465308;
srom_1(34956) <= 11016673;
srom_1(34957) <= 11555714;
srom_1(34958) <= 12079903;
srom_1(34959) <= 12586783;
srom_1(34960) <= 13073976;
srom_1(34961) <= 13539197;
srom_1(34962) <= 13980266;
srom_1(34963) <= 14395113;
srom_1(34964) <= 14781794;
srom_1(34965) <= 15138495;
srom_1(34966) <= 15463544;
srom_1(34967) <= 15755415;
srom_1(34968) <= 16012742;
srom_1(34969) <= 16234315;
srom_1(34970) <= 16419098;
srom_1(34971) <= 16566223;
srom_1(34972) <= 16675001;
srom_1(34973) <= 16744920;
srom_1(34974) <= 16775654;
srom_1(34975) <= 16767058;
srom_1(34976) <= 16719173;
srom_1(34977) <= 16632223;
srom_1(34978) <= 16506616;
srom_1(34979) <= 16342940;
srom_1(34980) <= 16141964;
srom_1(34981) <= 15904630;
srom_1(34982) <= 15632051;
srom_1(34983) <= 15325505;
srom_1(34984) <= 14986429;
srom_1(34985) <= 14616413;
srom_1(34986) <= 14217194;
srom_1(34987) <= 13790642;
srom_1(34988) <= 13338758;
srom_1(34989) <= 12863661;
srom_1(34990) <= 12367579;
srom_1(34991) <= 11852839;
srom_1(34992) <= 11321853;
srom_1(34993) <= 10777112;
srom_1(34994) <= 10221171;
srom_1(34995) <= 9656636;
srom_1(34996) <= 9086155;
srom_1(34997) <= 8512403;
srom_1(34998) <= 7938071;
srom_1(34999) <= 7365851;
srom_1(35000) <= 6798427;
srom_1(35001) <= 6238460;
srom_1(35002) <= 5688576;
srom_1(35003) <= 5151354;
srom_1(35004) <= 4629312;
srom_1(35005) <= 4124898;
srom_1(35006) <= 3640479;
srom_1(35007) <= 3178325;
srom_1(35008) <= 2740604;
srom_1(35009) <= 2329368;
srom_1(35010) <= 1946546;
srom_1(35011) <= 1593933;
srom_1(35012) <= 1273183;
srom_1(35013) <= 985800;
srom_1(35014) <= 733130;
srom_1(35015) <= 516360;
srom_1(35016) <= 336506;
srom_1(35017) <= 194410;
srom_1(35018) <= 90740;
srom_1(35019) <= 25982;
srom_1(35020) <= 439;
srom_1(35021) <= 14231;
srom_1(35022) <= 67293;
srom_1(35023) <= 159376;
srom_1(35024) <= 290050;
srom_1(35025) <= 458700;
srom_1(35026) <= 664536;
srom_1(35027) <= 906593;
srom_1(35028) <= 1183736;
srom_1(35029) <= 1494665;
srom_1(35030) <= 1837922;
srom_1(35031) <= 2211898;
srom_1(35032) <= 2614838;
srom_1(35033) <= 3044853;
srom_1(35034) <= 3499927;
srom_1(35035) <= 3977926;
srom_1(35036) <= 4476608;
srom_1(35037) <= 4993634;
srom_1(35038) <= 5526581;
srom_1(35039) <= 6072949;
srom_1(35040) <= 6630176;
srom_1(35041) <= 7195648;
srom_1(35042) <= 7766715;
srom_1(35043) <= 8340698;
srom_1(35044) <= 8914906;
srom_1(35045) <= 9486646;
srom_1(35046) <= 10053236;
srom_1(35047) <= 10612021;
srom_1(35048) <= 11160379;
srom_1(35049) <= 11695740;
srom_1(35050) <= 12215592;
srom_1(35051) <= 12717498;
srom_1(35052) <= 13199105;
srom_1(35053) <= 13658153;
srom_1(35054) <= 14092491;
srom_1(35055) <= 14500081;
srom_1(35056) <= 14879012;
srom_1(35057) <= 15227508;
srom_1(35058) <= 15543934;
srom_1(35059) <= 15826806;
srom_1(35060) <= 16074797;
srom_1(35061) <= 16286746;
srom_1(35062) <= 16461657;
srom_1(35063) <= 16598711;
srom_1(35064) <= 16697265;
srom_1(35065) <= 16756857;
srom_1(35066) <= 16777208;
srom_1(35067) <= 16758221;
srom_1(35068) <= 16699986;
srom_1(35069) <= 16602777;
srom_1(35070) <= 16467048;
srom_1(35071) <= 16293437;
srom_1(35072) <= 16082757;
srom_1(35073) <= 15835997;
srom_1(35074) <= 15554313;
srom_1(35075) <= 15239027;
srom_1(35076) <= 14891617;
srom_1(35077) <= 14513712;
srom_1(35078) <= 14107084;
srom_1(35079) <= 13673641;
srom_1(35080) <= 13215414;
srom_1(35081) <= 12734552;
srom_1(35082) <= 12233311;
srom_1(35083) <= 11714041;
srom_1(35084) <= 11179177;
srom_1(35085) <= 10631227;
srom_1(35086) <= 10072760;
srom_1(35087) <= 9506396;
srom_1(35088) <= 8934790;
srom_1(35089) <= 8360622;
srom_1(35090) <= 7786586;
srom_1(35091) <= 7215374;
srom_1(35092) <= 6649662;
srom_1(35093) <= 6092106;
srom_1(35094) <= 5545318;
srom_1(35095) <= 5011864;
srom_1(35096) <= 4494244;
srom_1(35097) <= 3994886;
srom_1(35098) <= 3516132;
srom_1(35099) <= 3060227;
srom_1(35100) <= 2629308;
srom_1(35101) <= 2225397;
srom_1(35102) <= 1850387;
srom_1(35103) <= 1506036;
srom_1(35104) <= 1193961;
srom_1(35105) <= 915624;
srom_1(35106) <= 672330;
srom_1(35107) <= 465221;
srom_1(35108) <= 295267;
srom_1(35109) <= 163265;
srom_1(35110) <= 69835;
srom_1(35111) <= 15414;
srom_1(35112) <= 259;
srom_1(35113) <= 24439;
srom_1(35114) <= 87841;
srom_1(35115) <= 190169;
srom_1(35116) <= 330942;
srom_1(35117) <= 509500;
srom_1(35118) <= 725006;
srom_1(35119) <= 976449;
srom_1(35120) <= 1262650;
srom_1(35121) <= 1582268;
srom_1(35122) <= 1933803;
srom_1(35123) <= 2315606;
srom_1(35124) <= 2725888;
srom_1(35125) <= 3162724;
srom_1(35126) <= 3624066;
srom_1(35127) <= 4107751;
srom_1(35128) <= 4611510;
srom_1(35129) <= 5132982;
srom_1(35130) <= 5669720;
srom_1(35131) <= 6219208;
srom_1(35132) <= 6778869;
srom_1(35133) <= 7346078;
srom_1(35134) <= 7918176;
srom_1(35135) <= 8492481;
srom_1(35136) <= 9066298;
srom_1(35137) <= 9636937;
srom_1(35138) <= 10201723;
srom_1(35139) <= 10758006;
srom_1(35140) <= 11303178;
srom_1(35141) <= 11834683;
srom_1(35142) <= 12350027;
srom_1(35143) <= 12846796;
srom_1(35144) <= 13322658;
srom_1(35145) <= 13775383;
srom_1(35146) <= 14202848;
srom_1(35147) <= 14603048;
srom_1(35148) <= 14974105;
srom_1(35149) <= 15314282;
srom_1(35150) <= 15621981;
srom_1(35151) <= 15895761;
srom_1(35152) <= 16134337;
srom_1(35153) <= 16336590;
srom_1(35154) <= 16501573;
srom_1(35155) <= 16628511;
srom_1(35156) <= 16716810;
srom_1(35157) <= 16766055;
srom_1(35158) <= 16776015;
srom_1(35159) <= 16746643;
srom_1(35160) <= 16678078;
srom_1(35161) <= 16570641;
srom_1(35162) <= 16424835;
srom_1(35163) <= 16241345;
srom_1(35164) <= 16021030;
srom_1(35165) <= 15764925;
srom_1(35166) <= 15474229;
srom_1(35167) <= 15150306;
srom_1(35168) <= 14794676;
srom_1(35169) <= 14409005;
srom_1(35170) <= 13995103;
srom_1(35171) <= 13554909;
srom_1(35172) <= 13090489;
srom_1(35173) <= 12604021;
srom_1(35174) <= 12097785;
srom_1(35175) <= 11574155;
srom_1(35176) <= 11035587;
srom_1(35177) <= 10484607;
srom_1(35178) <= 9923797;
srom_1(35179) <= 9355789;
srom_1(35180) <= 8783245;
srom_1(35181) <= 8208851;
srom_1(35182) <= 7635299;
srom_1(35183) <= 7065280;
srom_1(35184) <= 6501467;
srom_1(35185) <= 5946503;
srom_1(35186) <= 5402991;
srom_1(35187) <= 4873479;
srom_1(35188) <= 4360451;
srom_1(35189) <= 3866313;
srom_1(35190) <= 3393381;
srom_1(35191) <= 2943873;
srom_1(35192) <= 2519898;
srom_1(35193) <= 2123443;
srom_1(35194) <= 1756368;
srom_1(35195) <= 1420393;
srom_1(35196) <= 1117095;
srom_1(35197) <= 847895;
srom_1(35198) <= 614056;
srom_1(35199) <= 416675;
srom_1(35200) <= 256677;
srom_1(35201) <= 134813;
srom_1(35202) <= 51653;
srom_1(35203) <= 7588;
srom_1(35204) <= 2825;
srom_1(35205) <= 37385;
srom_1(35206) <= 111107;
srom_1(35207) <= 223645;
srom_1(35208) <= 374472;
srom_1(35209) <= 562879;
srom_1(35210) <= 787984;
srom_1(35211) <= 1048731;
srom_1(35212) <= 1343898;
srom_1(35213) <= 1672099;
srom_1(35214) <= 2031796;
srom_1(35215) <= 2421303;
srom_1(35216) <= 2838792;
srom_1(35217) <= 3282306;
srom_1(35218) <= 3749766;
srom_1(35219) <= 4238978;
srom_1(35220) <= 4747650;
srom_1(35221) <= 5273395;
srom_1(35222) <= 5813749;
srom_1(35223) <= 6366177;
srom_1(35224) <= 6928088;
srom_1(35225) <= 7496849;
srom_1(35226) <= 8069792;
srom_1(35227) <= 8644229;
srom_1(35228) <= 9217468;
srom_1(35229) <= 9786820;
srom_1(35230) <= 10349615;
srom_1(35231) <= 10903215;
srom_1(35232) <= 11445022;
srom_1(35233) <= 11972497;
srom_1(35234) <= 12483166;
srom_1(35235) <= 12974634;
srom_1(35236) <= 13444597;
srom_1(35237) <= 13890850;
srom_1(35238) <= 14311302;
srom_1(35239) <= 14703980;
srom_1(35240) <= 15067043;
srom_1(35241) <= 15398788;
srom_1(35242) <= 15697660;
srom_1(35243) <= 15962258;
srom_1(35244) <= 16191340;
srom_1(35245) <= 16383833;
srom_1(35246) <= 16538833;
srom_1(35247) <= 16655614;
srom_1(35248) <= 16733628;
srom_1(35249) <= 16772509;
srom_1(35250) <= 16772076;
srom_1(35251) <= 16732329;
srom_1(35252) <= 16653456;
srom_1(35253) <= 16535826;
srom_1(35254) <= 16379991;
srom_1(35255) <= 16186682;
srom_1(35256) <= 15956805;
srom_1(35257) <= 15691438;
srom_1(35258) <= 15391825;
srom_1(35259) <= 15059372;
srom_1(35260) <= 14695638;
srom_1(35261) <= 14302327;
srom_1(35262) <= 13881285;
srom_1(35263) <= 13434486;
srom_1(35264) <= 12964026;
srom_1(35265) <= 12472109;
srom_1(35266) <= 11961044;
srom_1(35267) <= 11433226;
srom_1(35268) <= 10891131;
srom_1(35269) <= 10337301;
srom_1(35270) <= 9774332;
srom_1(35271) <= 9204866;
srom_1(35272) <= 8631571;
srom_1(35273) <= 8057138;
srom_1(35274) <= 7484259;
srom_1(35275) <= 6915620;
srom_1(35276) <= 6353889;
srom_1(35277) <= 5801700;
srom_1(35278) <= 5261641;
srom_1(35279) <= 4736246;
srom_1(35280) <= 4227977;
srom_1(35281) <= 3739220;
srom_1(35282) <= 3272265;
srom_1(35283) <= 2829302;
srom_1(35284) <= 2412409;
srom_1(35285) <= 2023541;
srom_1(35286) <= 1664520;
srom_1(35287) <= 1337031;
srom_1(35288) <= 1042609;
srom_1(35289) <= 782635;
srom_1(35290) <= 558328;
srom_1(35291) <= 370740;
srom_1(35292) <= 220750;
srom_1(35293) <= 109062;
srom_1(35294) <= 36200;
srom_1(35295) <= 2506;
srom_1(35296) <= 8136;
srom_1(35297) <= 53066;
srom_1(35298) <= 137083;
srom_1(35299) <= 259795;
srom_1(35300) <= 420626;
srom_1(35301) <= 618821;
srom_1(35302) <= 853451;
srom_1(35303) <= 1123417;
srom_1(35304) <= 1427451;
srom_1(35305) <= 1764129;
srom_1(35306) <= 2131871;
srom_1(35307) <= 2528953;
srom_1(35308) <= 2953513;
srom_1(35309) <= 3403560;
srom_1(35310) <= 3876984;
srom_1(35311) <= 4371564;
srom_1(35312) <= 4884981;
srom_1(35313) <= 5414828;
srom_1(35314) <= 5958620;
srom_1(35315) <= 6513808;
srom_1(35316) <= 7077787;
srom_1(35317) <= 7647912;
srom_1(35318) <= 8221511;
srom_1(35319) <= 8795894;
srom_1(35320) <= 9368367;
srom_1(35321) <= 9936245;
srom_1(35322) <= 10496866;
srom_1(35323) <= 11047600;
srom_1(35324) <= 11585866;
srom_1(35325) <= 12109139;
srom_1(35326) <= 12614964;
srom_1(35327) <= 13100971;
srom_1(35328) <= 13564880;
srom_1(35329) <= 14004516;
srom_1(35330) <= 14417816;
srom_1(35331) <= 14802844;
srom_1(35332) <= 15157793;
srom_1(35333) <= 15480999;
srom_1(35334) <= 15770947;
srom_1(35335) <= 16026276;
srom_1(35336) <= 16245789;
srom_1(35337) <= 16428458;
srom_1(35338) <= 16573424;
srom_1(35339) <= 16680010;
srom_1(35340) <= 16747714;
srom_1(35341) <= 16776219;
srom_1(35342) <= 16765392;
srom_1(35343) <= 16715284;
srom_1(35344) <= 16626128;
srom_1(35345) <= 16498344;
srom_1(35346) <= 16332531;
srom_1(35347) <= 16129466;
srom_1(35348) <= 15890102;
srom_1(35349) <= 15615560;
srom_1(35350) <= 15307129;
srom_1(35351) <= 14966254;
srom_1(35352) <= 14594534;
srom_1(35353) <= 14193713;
srom_1(35354) <= 13765670;
srom_1(35355) <= 13312412;
srom_1(35356) <= 12836064;
srom_1(35357) <= 12338861;
srom_1(35358) <= 11823133;
srom_1(35359) <= 11291300;
srom_1(35360) <= 10745855;
srom_1(35361) <= 10189357;
srom_1(35362) <= 9624413;
srom_1(35363) <= 9053675;
srom_1(35364) <= 8479818;
srom_1(35365) <= 7905534;
srom_1(35366) <= 7333514;
srom_1(35367) <= 6766442;
srom_1(35368) <= 6206978;
srom_1(35369) <= 5657743;
srom_1(35370) <= 5121315;
srom_1(35371) <= 4600208;
srom_1(35372) <= 4096866;
srom_1(35373) <= 3613649;
srom_1(35374) <= 3152824;
srom_1(35375) <= 2716552;
srom_1(35376) <= 2306877;
srom_1(35377) <= 1925722;
srom_1(35378) <= 1574874;
srom_1(35379) <= 1255977;
srom_1(35380) <= 970528;
srom_1(35381) <= 719865;
srom_1(35382) <= 505163;
srom_1(35383) <= 327429;
srom_1(35384) <= 187497;
srom_1(35385) <= 86023;
srom_1(35386) <= 23482;
srom_1(35387) <= 169;
srom_1(35388) <= 16191;
srom_1(35389) <= 71475;
srom_1(35390) <= 165761;
srom_1(35391) <= 298606;
srom_1(35392) <= 469388;
srom_1(35393) <= 677306;
srom_1(35394) <= 921385;
srom_1(35395) <= 1200481;
srom_1(35396) <= 1513284;
srom_1(35397) <= 1858328;
srom_1(35398) <= 2233994;
srom_1(35399) <= 2638522;
srom_1(35400) <= 3070013;
srom_1(35401) <= 3526446;
srom_1(35402) <= 4005679;
srom_1(35403) <= 4505464;
srom_1(35404) <= 5023460;
srom_1(35405) <= 5557235;
srom_1(35406) <= 6104288;
srom_1(35407) <= 6662053;
srom_1(35408) <= 7227914;
srom_1(35409) <= 7799218;
srom_1(35410) <= 8373286;
srom_1(35411) <= 8947425;
srom_1(35412) <= 9518945;
srom_1(35413) <= 10085163;
srom_1(35414) <= 10643426;
srom_1(35415) <= 11191116;
srom_1(35416) <= 11725663;
srom_1(35417) <= 12244562;
srom_1(35418) <= 12745379;
srom_1(35419) <= 13225765;
srom_1(35420) <= 13683469;
srom_1(35421) <= 14116343;
srom_1(35422) <= 14522357;
srom_1(35423) <= 14899609;
srom_1(35424) <= 15246328;
srom_1(35425) <= 15560889;
srom_1(35426) <= 15841816;
srom_1(35427) <= 16087793;
srom_1(35428) <= 16297666;
srom_1(35429) <= 16470450;
srom_1(35430) <= 16605336;
srom_1(35431) <= 16701691;
srom_1(35432) <= 16759063;
srom_1(35433) <= 16777183;
srom_1(35434) <= 16755966;
srom_1(35435) <= 16695512;
srom_1(35436) <= 16596103;
srom_1(35437) <= 16458207;
srom_1(35438) <= 16282470;
srom_1(35439) <= 16069716;
srom_1(35440) <= 15820942;
srom_1(35441) <= 15537316;
srom_1(35442) <= 15220167;
srom_1(35443) <= 14870982;
srom_1(35444) <= 14491400;
srom_1(35445) <= 14083199;
srom_1(35446) <= 13648294;
srom_1(35447) <= 13188725;
srom_1(35448) <= 12706646;
srom_1(35449) <= 12204319;
srom_1(35450) <= 11684098;
srom_1(35451) <= 11148424;
srom_1(35452) <= 10599808;
srom_1(35453) <= 10040823;
srom_1(35454) <= 9474090;
srom_1(35455) <= 8902267;
srom_1(35456) <= 8328035;
srom_1(35457) <= 7754087;
srom_1(35458) <= 7183115;
srom_1(35459) <= 6617796;
srom_1(35460) <= 6060780;
srom_1(35461) <= 5514681;
srom_1(35462) <= 4982058;
srom_1(35463) <= 4465410;
srom_1(35464) <= 3967159;
srom_1(35465) <= 3489642;
srom_1(35466) <= 3035098;
srom_1(35467) <= 2605658;
srom_1(35468) <= 2203336;
srom_1(35469) <= 1830019;
srom_1(35470) <= 1487458;
srom_1(35471) <= 1177259;
srom_1(35472) <= 900876;
srom_1(35473) <= 659605;
srom_1(35474) <= 454579;
srom_1(35475) <= 286758;
srom_1(35476) <= 156929;
srom_1(35477) <= 65701;
srom_1(35478) <= 13503;
srom_1(35479) <= 578;
srom_1(35480) <= 26987;
srom_1(35481) <= 92607;
srom_1(35482) <= 197130;
srom_1(35483) <= 340066;
srom_1(35484) <= 520743;
srom_1(35485) <= 738316;
srom_1(35486) <= 991764;
srom_1(35487) <= 1279898;
srom_1(35488) <= 1601367;
srom_1(35489) <= 1954664;
srom_1(35490) <= 2338132;
srom_1(35491) <= 2749973;
srom_1(35492) <= 3188255;
srom_1(35493) <= 3650923;
srom_1(35494) <= 4135808;
srom_1(35495) <= 4640636;
srom_1(35496) <= 5163040;
srom_1(35497) <= 5700569;
srom_1(35498) <= 6250703;
srom_1(35499) <= 6810863;
srom_1(35500) <= 7378421;
srom_1(35501) <= 7950716;
srom_1(35502) <= 8525065;
srom_1(35503) <= 9098774;
srom_1(35504) <= 9669153;
srom_1(35505) <= 10233526;
srom_1(35506) <= 10789249;
srom_1(35507) <= 11333713;
srom_1(35508) <= 11864368;
srom_1(35509) <= 12378723;
srom_1(35510) <= 12874367;
srom_1(35511) <= 13348976;
srom_1(35512) <= 13800324;
srom_1(35513) <= 14226294;
srom_1(35514) <= 14624890;
srom_1(35515) <= 14994242;
srom_1(35516) <= 15332617;
srom_1(35517) <= 15638430;
srom_1(35518) <= 15910245;
srom_1(35519) <= 16146790;
srom_1(35520) <= 16346953;
srom_1(35521) <= 16509797;
srom_1(35522) <= 16634558;
srom_1(35523) <= 16720651;
srom_1(35524) <= 16767672;
srom_1(35525) <= 16775400;
srom_1(35526) <= 16743801;
srom_1(35527) <= 16673020;
srom_1(35528) <= 16563392;
srom_1(35529) <= 16415429;
srom_1(35530) <= 16229825;
srom_1(35531) <= 16007451;
srom_1(35532) <= 15749350;
srom_1(35533) <= 15456732;
srom_1(35534) <= 15130969;
srom_1(35535) <= 14773588;
srom_1(35536) <= 14386267;
srom_1(35537) <= 13970820;
srom_1(35538) <= 13529196;
srom_1(35539) <= 13063466;
srom_1(35540) <= 12575815;
srom_1(35541) <= 12068528;
srom_1(35542) <= 11543984;
srom_1(35543) <= 11004644;
srom_1(35544) <= 10453037;
srom_1(35545) <= 9891748;
srom_1(35546) <= 9323411;
srom_1(35547) <= 8750691;
srom_1(35548) <= 8176272;
srom_1(35549) <= 7602849;
srom_1(35550) <= 7033111;
srom_1(35551) <= 6469729;
srom_1(35552) <= 5915345;
srom_1(35553) <= 5372559;
srom_1(35554) <= 4843917;
srom_1(35555) <= 4331897;
srom_1(35556) <= 3838900;
srom_1(35557) <= 3367239;
srom_1(35558) <= 2919124;
srom_1(35559) <= 2496657;
srom_1(35560) <= 2101820;
srom_1(35561) <= 1736464;
srom_1(35562) <= 1402302;
srom_1(35563) <= 1100901;
srom_1(35564) <= 833675;
srom_1(35565) <= 601876;
srom_1(35566) <= 406592;
srom_1(35567) <= 248739;
srom_1(35568) <= 129056;
srom_1(35569) <= 48105;
srom_1(35570) <= 6265;
srom_1(35571) <= 3734;
srom_1(35572) <= 40521;
srom_1(35573) <= 116456;
srom_1(35574) <= 231182;
srom_1(35575) <= 384160;
srom_1(35576) <= 574675;
srom_1(35577) <= 801831;
srom_1(35578) <= 1064564;
srom_1(35579) <= 1361643;
srom_1(35580) <= 1691673;
srom_1(35581) <= 2053108;
srom_1(35582) <= 2444251;
srom_1(35583) <= 2863270;
srom_1(35584) <= 3308199;
srom_1(35585) <= 3776952;
srom_1(35586) <= 4267331;
srom_1(35587) <= 4777035;
srom_1(35588) <= 5303676;
srom_1(35589) <= 5844783;
srom_1(35590) <= 6397818;
srom_1(35591) <= 6960190;
srom_1(35592) <= 7529259;
srom_1(35593) <= 8102358;
srom_1(35594) <= 8676800;
srom_1(35595) <= 9249890;
srom_1(35596) <= 9818941;
srom_1(35597) <= 10381285;
srom_1(35598) <= 10934285;
srom_1(35599) <= 11475347;
srom_1(35600) <= 12001934;
srom_1(35601) <= 12511577;
srom_1(35602) <= 13001886;
srom_1(35603) <= 13470562;
srom_1(35604) <= 13915407;
srom_1(35605) <= 14334335;
srom_1(35606) <= 14725381;
srom_1(35607) <= 15086712;
srom_1(35608) <= 15416633;
srom_1(35609) <= 15713597;
srom_1(35610) <= 15976212;
srom_1(35611) <= 16203246;
srom_1(35612) <= 16393635;
srom_1(35613) <= 16546485;
srom_1(35614) <= 16661080;
srom_1(35615) <= 16736883;
srom_1(35616) <= 16773537;
srom_1(35617) <= 16770872;
srom_1(35618) <= 16728900;
srom_1(35619) <= 16647817;
srom_1(35620) <= 16528003;
srom_1(35621) <= 16370022;
srom_1(35622) <= 16174612;
srom_1(35623) <= 15942692;
srom_1(35624) <= 15675348;
srom_1(35625) <= 15373833;
srom_1(35626) <= 15039563;
srom_1(35627) <= 14674104;
srom_1(35628) <= 14279170;
srom_1(35629) <= 13856613;
srom_1(35630) <= 13408415;
srom_1(35631) <= 12936678;
srom_1(35632) <= 12443612;
srom_1(35633) <= 11931532;
srom_1(35634) <= 11402837;
srom_1(35635) <= 10860008;
srom_1(35636) <= 10305590;
srom_1(35637) <= 9742182;
srom_1(35638) <= 9172426;
srom_1(35639) <= 8598996;
srom_1(35640) <= 8024578;
srom_1(35641) <= 7451868;
srom_1(35642) <= 6883550;
srom_1(35643) <= 6322290;
srom_1(35644) <= 5770720;
srom_1(35645) <= 5231425;
srom_1(35646) <= 4706936;
srom_1(35647) <= 4199712;
srom_1(35648) <= 3712131;
srom_1(35649) <= 3246479;
srom_1(35650) <= 2804941;
srom_1(35651) <= 2389586;
srom_1(35652) <= 2002363;
srom_1(35653) <= 1645087;
srom_1(35654) <= 1319433;
srom_1(35655) <= 1026930;
srom_1(35656) <= 768948;
srom_1(35657) <= 546697;
srom_1(35658) <= 361219;
srom_1(35659) <= 213385;
srom_1(35660) <= 103887;
srom_1(35661) <= 33239;
srom_1(35662) <= 1772;
srom_1(35663) <= 9634;
srom_1(35664) <= 56788;
srom_1(35665) <= 143013;
srom_1(35666) <= 267904;
srom_1(35667) <= 430875;
srom_1(35668) <= 631164;
srom_1(35669) <= 867829;
srom_1(35670) <= 1139763;
srom_1(35671) <= 1445688;
srom_1(35672) <= 1784171;
srom_1(35673) <= 2153625;
srom_1(35674) <= 2552316;
srom_1(35675) <= 2978376;
srom_1(35676) <= 3429807;
srom_1(35677) <= 3904491;
srom_1(35678) <= 4400202;
srom_1(35679) <= 4914617;
srom_1(35680) <= 5445322;
srom_1(35681) <= 5989829;
srom_1(35682) <= 6545585;
srom_1(35683) <= 7109984;
srom_1(35684) <= 7680378;
srom_1(35685) <= 8254094;
srom_1(35686) <= 8828440;
srom_1(35687) <= 9400724;
srom_1(35688) <= 9968262;
srom_1(35689) <= 10528392;
srom_1(35690) <= 11078488;
srom_1(35691) <= 11615970;
srom_1(35692) <= 12138318;
srom_1(35693) <= 12643082;
srom_1(35694) <= 13127896;
srom_1(35695) <= 13590485;
srom_1(35696) <= 14028681;
srom_1(35697) <= 14440429;
srom_1(35698) <= 14823797;
srom_1(35699) <= 15176989;
srom_1(35700) <= 15498348;
srom_1(35701) <= 15786367;
srom_1(35702) <= 16039695;
srom_1(35703) <= 16257144;
srom_1(35704) <= 16437696;
srom_1(35705) <= 16580502;
srom_1(35706) <= 16684894;
srom_1(35707) <= 16750381;
srom_1(35708) <= 16776658;
srom_1(35709) <= 16763600;
srom_1(35710) <= 16711268;
srom_1(35711) <= 16619909;
srom_1(35712) <= 16489950;
srom_1(35713) <= 16322002;
srom_1(35714) <= 16116851;
srom_1(35715) <= 15875460;
srom_1(35716) <= 15598960;
srom_1(35717) <= 15288648;
srom_1(35718) <= 14945980;
srom_1(35719) <= 14572562;
srom_1(35720) <= 14170145;
srom_1(35721) <= 13740617;
srom_1(35722) <= 13285991;
srom_1(35723) <= 12808400;
srom_1(35724) <= 12310082;
srom_1(35725) <= 11793376;
srom_1(35726) <= 11260704;
srom_1(35727) <= 10714563;
srom_1(35728) <= 10157515;
srom_1(35729) <= 9592172;
srom_1(35730) <= 9021185;
srom_1(35731) <= 8447232;
srom_1(35732) <= 7873003;
srom_1(35733) <= 7301193;
srom_1(35734) <= 6734482;
srom_1(35735) <= 6175528;
srom_1(35736) <= 5626951;
srom_1(35737) <= 5091325;
srom_1(35738) <= 4571161;
srom_1(35739) <= 4068898;
srom_1(35740) <= 3586892;
srom_1(35741) <= 3127403;
srom_1(35742) <= 2692585;
srom_1(35743) <= 2284478;
srom_1(35744) <= 1904996;
srom_1(35745) <= 1555917;
srom_1(35746) <= 1238879;
srom_1(35747) <= 955368;
srom_1(35748) <= 706715;
srom_1(35749) <= 494084;
srom_1(35750) <= 318474;
srom_1(35751) <= 180708;
srom_1(35752) <= 81431;
srom_1(35753) <= 21109;
srom_1(35754) <= 25;
srom_1(35755) <= 18278;
srom_1(35756) <= 75783;
srom_1(35757) <= 172269;
srom_1(35758) <= 307284;
srom_1(35759) <= 480196;
srom_1(35760) <= 690193;
srom_1(35761) <= 936290;
srom_1(35762) <= 1217334;
srom_1(35763) <= 1532006;
srom_1(35764) <= 1878832;
srom_1(35765) <= 2256184;
srom_1(35766) <= 2662292;
srom_1(35767) <= 3095254;
srom_1(35768) <= 3553038;
srom_1(35769) <= 4033497;
srom_1(35770) <= 4534380;
srom_1(35771) <= 5053336;
srom_1(35772) <= 5587932;
srom_1(35773) <= 6135661;
srom_1(35774) <= 6693956;
srom_1(35775) <= 7260197;
srom_1(35776) <= 7831729;
srom_1(35777) <= 8405874;
srom_1(35778) <= 8979937;
srom_1(35779) <= 9551227;
srom_1(35780) <= 10117065;
srom_1(35781) <= 10674798;
srom_1(35782) <= 11221810;
srom_1(35783) <= 11755536;
srom_1(35784) <= 12273474;
srom_1(35785) <= 12773194;
srom_1(35786) <= 13252353;
srom_1(35787) <= 13708705;
srom_1(35788) <= 14140108;
srom_1(35789) <= 14544541;
srom_1(35790) <= 14920107;
srom_1(35791) <= 15265044;
srom_1(35792) <= 15577735;
srom_1(35793) <= 15856714;
srom_1(35794) <= 16100673;
srom_1(35795) <= 16308466;
srom_1(35796) <= 16479121;
srom_1(35797) <= 16611837;
srom_1(35798) <= 16705991;
srom_1(35799) <= 16761142;
srom_1(35800) <= 16777032;
srom_1(35801) <= 16753585;
srom_1(35802) <= 16690912;
srom_1(35803) <= 16589306;
srom_1(35804) <= 16449245;
srom_1(35805) <= 16271385;
srom_1(35806) <= 16056559;
srom_1(35807) <= 15805776;
srom_1(35808) <= 15520211;
srom_1(35809) <= 15201204;
srom_1(35810) <= 14850250;
srom_1(35811) <= 14468995;
srom_1(35812) <= 14059227;
srom_1(35813) <= 13622868;
srom_1(35814) <= 13161963;
srom_1(35815) <= 12678675;
srom_1(35816) <= 12175269;
srom_1(35817) <= 11654106;
srom_1(35818) <= 11117630;
srom_1(35819) <= 10568356;
srom_1(35820) <= 10008861;
srom_1(35821) <= 9441768;
srom_1(35822) <= 8869736;
srom_1(35823) <= 8295449;
srom_1(35824) <= 7721598;
srom_1(35825) <= 7150875;
srom_1(35826) <= 6585956;
srom_1(35827) <= 6029490;
srom_1(35828) <= 5484087;
srom_1(35829) <= 4952304;
srom_1(35830) <= 4436636;
srom_1(35831) <= 3939499;
srom_1(35832) <= 3463226;
srom_1(35833) <= 3010049;
srom_1(35834) <= 2582095;
srom_1(35835) <= 2181369;
srom_1(35836) <= 1809751;
srom_1(35837) <= 1468984;
srom_1(35838) <= 1160665;
srom_1(35839) <= 886241;
srom_1(35840) <= 646997;
srom_1(35841) <= 444057;
srom_1(35842) <= 278371;
srom_1(35843) <= 150717;
srom_1(35844) <= 61694;
srom_1(35845) <= 11718;
srom_1(35846) <= 1024;
srom_1(35847) <= 29662;
srom_1(35848) <= 97499;
srom_1(35849) <= 204215;
srom_1(35850) <= 349311;
srom_1(35851) <= 532106;
srom_1(35852) <= 751742;
srom_1(35853) <= 1007191;
srom_1(35854) <= 1297253;
srom_1(35855) <= 1620569;
srom_1(35856) <= 1975623;
srom_1(35857) <= 2360750;
srom_1(35858) <= 2774143;
srom_1(35859) <= 3213865;
srom_1(35860) <= 3677852;
srom_1(35861) <= 4163930;
srom_1(35862) <= 4669819;
srom_1(35863) <= 5193146;
srom_1(35864) <= 5731459;
srom_1(35865) <= 6282231;
srom_1(35866) <= 6842881;
srom_1(35867) <= 7410779;
srom_1(35868) <= 7983263;
srom_1(35869) <= 8557648;
srom_1(35870) <= 9131239;
srom_1(35871) <= 9701349;
srom_1(35872) <= 10265302;
srom_1(35873) <= 10820455;
srom_1(35874) <= 11364205;
srom_1(35875) <= 11894000;
srom_1(35876) <= 12407358;
srom_1(35877) <= 12901870;
srom_1(35878) <= 13375218;
srom_1(35879) <= 13825182;
srom_1(35880) <= 14249653;
srom_1(35881) <= 14646638;
srom_1(35882) <= 15014278;
srom_1(35883) <= 15350848;
srom_1(35884) <= 15654769;
srom_1(35885) <= 15924617;
srom_1(35886) <= 16159125;
srom_1(35887) <= 16357196;
srom_1(35888) <= 16517898;
srom_1(35889) <= 16640480;
srom_1(35890) <= 16724366;
srom_1(35891) <= 16769162;
srom_1(35892) <= 16774660;
srom_1(35893) <= 16740832;
srom_1(35894) <= 16667838;
srom_1(35895) <= 16556019;
srom_1(35896) <= 16405901;
srom_1(35897) <= 16218187;
srom_1(35898) <= 15993757;
srom_1(35899) <= 15733664;
srom_1(35900) <= 15439128;
srom_1(35901) <= 15111529;
srom_1(35902) <= 14752405;
srom_1(35903) <= 14363438;
srom_1(35904) <= 13946453;
srom_1(35905) <= 13503405;
srom_1(35906) <= 13036373;
srom_1(35907) <= 12547545;
srom_1(35908) <= 12039215;
srom_1(35909) <= 11513766;
srom_1(35910) <= 10973662;
srom_1(35911) <= 10421436;
srom_1(35912) <= 9859677;
srom_1(35913) <= 9291019;
srom_1(35914) <= 8718130;
srom_1(35915) <= 8143696;
srom_1(35916) <= 7570410;
srom_1(35917) <= 7000961;
srom_1(35918) <= 6438019;
srom_1(35919) <= 5884225;
srom_1(35920) <= 5342174;
srom_1(35921) <= 4814408;
srom_1(35922) <= 4303404;
srom_1(35923) <= 3811556;
srom_1(35924) <= 3341172;
srom_1(35925) <= 2894457;
srom_1(35926) <= 2473506;
srom_1(35927) <= 2080292;
srom_1(35928) <= 1716661;
srom_1(35929) <= 1384317;
srom_1(35930) <= 1084818;
srom_1(35931) <= 819569;
srom_1(35932) <= 589814;
srom_1(35933) <= 396630;
srom_1(35934) <= 240923;
srom_1(35935) <= 123424;
srom_1(35936) <= 44683;
srom_1(35937) <= 5069;
srom_1(35938) <= 4769;
srom_1(35939) <= 43783;
srom_1(35940) <= 121930;
srom_1(35941) <= 238841;
srom_1(35942) <= 393969;
srom_1(35943) <= 586588;
srom_1(35944) <= 815792;
srom_1(35945) <= 1080508;
srom_1(35946) <= 1379494;
srom_1(35947) <= 1711348;
srom_1(35948) <= 2074515;
srom_1(35949) <= 2467290;
srom_1(35950) <= 2887832;
srom_1(35951) <= 3334169;
srom_1(35952) <= 3804208;
srom_1(35953) <= 4295746;
srom_1(35954) <= 4806476;
srom_1(35955) <= 5334003;
srom_1(35956) <= 5875855;
srom_1(35957) <= 6429490;
srom_1(35958) <= 6992312;
srom_1(35959) <= 7561682;
srom_1(35960) <= 8134929;
srom_1(35961) <= 8709366;
srom_1(35962) <= 9282299;
srom_1(35963) <= 9851041;
srom_1(35964) <= 10412925;
srom_1(35965) <= 10965317;
srom_1(35966) <= 11505625;
srom_1(35967) <= 12031317;
srom_1(35968) <= 12539926;
srom_1(35969) <= 13029069;
srom_1(35970) <= 13496451;
srom_1(35971) <= 13939880;
srom_1(35972) <= 14357278;
srom_1(35973) <= 14746687;
srom_1(35974) <= 15106280;
srom_1(35975) <= 15434372;
srom_1(35976) <= 15729424;
srom_1(35977) <= 15990052;
srom_1(35978) <= 16215034;
srom_1(35979) <= 16403316;
srom_1(35980) <= 16554014;
srom_1(35981) <= 16666421;
srom_1(35982) <= 16740011;
srom_1(35983) <= 16774439;
srom_1(35984) <= 16769542;
srom_1(35985) <= 16725344;
srom_1(35986) <= 16642053;
srom_1(35987) <= 16520058;
srom_1(35988) <= 16359932;
srom_1(35989) <= 16162426;
srom_1(35990) <= 15928465;
srom_1(35991) <= 15659148;
srom_1(35992) <= 15355736;
srom_1(35993) <= 15019654;
srom_1(35994) <= 14652476;
srom_1(35995) <= 14255924;
srom_1(35996) <= 13831859;
srom_1(35997) <= 13382268;
srom_1(35998) <= 12909261;
srom_1(35999) <= 12415054;
srom_1(36000) <= 11901967;
srom_1(36001) <= 11372403;
srom_1(36002) <= 10828848;
srom_1(36003) <= 10273850;
srom_1(36004) <= 9710011;
srom_1(36005) <= 9139975;
srom_1(36006) <= 8566416;
srom_1(36007) <= 7992024;
srom_1(36008) <= 7419491;
srom_1(36009) <= 6851502;
srom_1(36010) <= 6290722;
srom_1(36011) <= 5739779;
srom_1(36012) <= 5201258;
srom_1(36013) <= 4677683;
srom_1(36014) <= 4171510;
srom_1(36015) <= 3685112;
srom_1(36016) <= 3220770;
srom_1(36017) <= 2780663;
srom_1(36018) <= 2366853;
srom_1(36019) <= 1981281;
srom_1(36020) <= 1625755;
srom_1(36021) <= 1301942;
srom_1(36022) <= 1011362;
srom_1(36023) <= 755375;
srom_1(36024) <= 535184;
srom_1(36025) <= 351820;
srom_1(36026) <= 206143;
srom_1(36027) <= 98837;
srom_1(36028) <= 30404;
srom_1(36029) <= 1166;
srom_1(36030) <= 11259;
srom_1(36031) <= 60636;
srom_1(36032) <= 149067;
srom_1(36033) <= 276135;
srom_1(36034) <= 441245;
srom_1(36035) <= 643624;
srom_1(36036) <= 882321;
srom_1(36037) <= 1156218;
srom_1(36038) <= 1464030;
srom_1(36039) <= 1804313;
srom_1(36040) <= 2175473;
srom_1(36041) <= 2575768;
srom_1(36042) <= 3003322;
srom_1(36043) <= 3456129;
srom_1(36044) <= 3932066;
srom_1(36045) <= 4428901;
srom_1(36046) <= 4944305;
srom_1(36047) <= 5475860;
srom_1(36048) <= 6021074;
srom_1(36049) <= 6577391;
srom_1(36050) <= 7142200;
srom_1(36051) <= 7712855;
srom_1(36052) <= 8286678;
srom_1(36053) <= 8860980;
srom_1(36054) <= 9433066;
srom_1(36055) <= 10000255;
srom_1(36056) <= 10559885;
srom_1(36057) <= 11109334;
srom_1(36058) <= 11646025;
srom_1(36059) <= 12167440;
srom_1(36060) <= 12671135;
srom_1(36061) <= 13154748;
srom_1(36062) <= 13616011;
srom_1(36063) <= 14052761;
srom_1(36064) <= 14462949;
srom_1(36065) <= 14844653;
srom_1(36066) <= 15196083;
srom_1(36067) <= 15515589;
srom_1(36068) <= 15801675;
srom_1(36069) <= 16052998;
srom_1(36070) <= 16268381;
srom_1(36071) <= 16446812;
srom_1(36072) <= 16587456;
srom_1(36073) <= 16689653;
srom_1(36074) <= 16752923;
srom_1(36075) <= 16776969;
srom_1(36076) <= 16761680;
srom_1(36077) <= 16707127;
srom_1(36078) <= 16613566;
srom_1(36079) <= 16481434;
srom_1(36080) <= 16311353;
srom_1(36081) <= 16104119;
srom_1(36082) <= 15860705;
srom_1(36083) <= 15582251;
srom_1(36084) <= 15270064;
srom_1(36085) <= 14925607;
srom_1(36086) <= 14550496;
srom_1(36087) <= 14146490;
srom_1(36088) <= 13715483;
srom_1(36089) <= 13259496;
srom_1(36090) <= 12780669;
srom_1(36091) <= 12281245;
srom_1(36092) <= 11763568;
srom_1(36093) <= 11230064;
srom_1(36094) <= 10683235;
srom_1(36095) <= 10125647;
srom_1(36096) <= 9559912;
srom_1(36097) <= 8988685;
srom_1(36098) <= 8414644;
srom_1(36099) <= 7840481;
srom_1(36100) <= 7268889;
srom_1(36101) <= 6702547;
srom_1(36102) <= 6144111;
srom_1(36103) <= 5596201;
srom_1(36104) <= 5061385;
srom_1(36105) <= 4542172;
srom_1(36106) <= 4040996;
srom_1(36107) <= 3560208;
srom_1(36108) <= 3102061;
srom_1(36109) <= 2668705;
srom_1(36110) <= 2262171;
srom_1(36111) <= 1884367;
srom_1(36112) <= 1537063;
srom_1(36113) <= 1221888;
srom_1(36114) <= 940321;
srom_1(36115) <= 693681;
srom_1(36116) <= 483125;
srom_1(36117) <= 309641;
srom_1(36118) <= 174042;
srom_1(36119) <= 76964;
srom_1(36120) <= 18861;
srom_1(36121) <= 8;
srom_1(36122) <= 20491;
srom_1(36123) <= 80216;
srom_1(36124) <= 178901;
srom_1(36125) <= 316085;
srom_1(36126) <= 491123;
srom_1(36127) <= 703196;
srom_1(36128) <= 951307;
srom_1(36129) <= 1234295;
srom_1(36130) <= 1550832;
srom_1(36131) <= 1899434;
srom_1(36132) <= 2278465;
srom_1(36133) <= 2686150;
srom_1(36134) <= 3120575;
srom_1(36135) <= 3579703;
srom_1(36136) <= 4061382;
srom_1(36137) <= 4563353;
srom_1(36138) <= 5083262;
srom_1(36139) <= 5618671;
srom_1(36140) <= 6167069;
srom_1(36141) <= 6725884;
srom_1(36142) <= 7292497;
srom_1(36143) <= 7864250;
srom_1(36144) <= 8438461;
srom_1(36145) <= 9012439;
srom_1(36146) <= 9583491;
srom_1(36147) <= 10148940;
srom_1(36148) <= 10706135;
srom_1(36149) <= 11252461;
srom_1(36150) <= 11785358;
srom_1(36151) <= 12302327;
srom_1(36152) <= 12800943;
srom_1(36153) <= 13278867;
srom_1(36154) <= 13733860;
srom_1(36155) <= 14163787;
srom_1(36156) <= 14566632;
srom_1(36157) <= 14940506;
srom_1(36158) <= 15283657;
srom_1(36159) <= 15594473;
srom_1(36160) <= 15871500;
srom_1(36161) <= 16113436;
srom_1(36162) <= 16319148;
srom_1(36163) <= 16487670;
srom_1(36164) <= 16618214;
srom_1(36165) <= 16710166;
srom_1(36166) <= 16763095;
srom_1(36167) <= 16776754;
srom_1(36168) <= 16751078;
srom_1(36169) <= 16686187;
srom_1(36170) <= 16582386;
srom_1(36171) <= 16440161;
srom_1(36172) <= 16260180;
srom_1(36173) <= 16043287;
srom_1(36174) <= 15790498;
srom_1(36175) <= 15502999;
srom_1(36176) <= 15182138;
srom_1(36177) <= 14829420;
srom_1(36178) <= 14446499;
srom_1(36179) <= 14035170;
srom_1(36180) <= 13597363;
srom_1(36181) <= 13135130;
srom_1(36182) <= 12650639;
srom_1(36183) <= 12146161;
srom_1(36184) <= 11624064;
srom_1(36185) <= 11086794;
srom_1(36186) <= 10536871;
srom_1(36187) <= 9976875;
srom_1(36188) <= 9409430;
srom_1(36189) <= 8837199;
srom_1(36190) <= 8262864;
srom_1(36191) <= 7689118;
srom_1(36192) <= 7118653;
srom_1(36193) <= 6554143;
srom_1(36194) <= 5998235;
srom_1(36195) <= 5453537;
srom_1(36196) <= 4922602;
srom_1(36197) <= 4407921;
srom_1(36198) <= 3911906;
srom_1(36199) <= 3436884;
srom_1(36200) <= 2985082;
srom_1(36201) <= 2558620;
srom_1(36202) <= 2159496;
srom_1(36203) <= 1789583;
srom_1(36204) <= 1450614;
srom_1(36205) <= 1144181;
srom_1(36206) <= 871719;
srom_1(36207) <= 634506;
srom_1(36208) <= 433655;
srom_1(36209) <= 270107;
srom_1(36210) <= 144630;
srom_1(36211) <= 57811;
srom_1(36212) <= 10059;
srom_1(36213) <= 1597;
srom_1(36214) <= 32464;
srom_1(36215) <= 102516;
srom_1(36216) <= 211424;
srom_1(36217) <= 358678;
srom_1(36218) <= 543587;
srom_1(36219) <= 765283;
srom_1(36220) <= 1022729;
srom_1(36221) <= 1314715;
srom_1(36222) <= 1639874;
srom_1(36223) <= 1996679;
srom_1(36224) <= 2383458;
srom_1(36225) <= 2798398;
srom_1(36226) <= 3239552;
srom_1(36227) <= 3704852;
srom_1(36228) <= 4192115;
srom_1(36229) <= 4699057;
srom_1(36230) <= 5223301;
srom_1(36231) <= 5762388;
srom_1(36232) <= 6313790;
srom_1(36233) <= 6874922;
srom_1(36234) <= 7443152;
srom_1(36235) <= 8015816;
srom_1(36236) <= 8590227;
srom_1(36237) <= 9163694;
srom_1(36238) <= 9733525;
srom_1(36239) <= 10297050;
srom_1(36240) <= 10851625;
srom_1(36241) <= 11394651;
srom_1(36242) <= 11923580;
srom_1(36243) <= 12435932;
srom_1(36244) <= 12929305;
srom_1(36245) <= 13401385;
srom_1(36246) <= 13849959;
srom_1(36247) <= 14272922;
srom_1(36248) <= 14668292;
srom_1(36249) <= 15034214;
srom_1(36250) <= 15368973;
srom_1(36251) <= 15670998;
srom_1(36252) <= 15938874;
srom_1(36253) <= 16171344;
srom_1(36254) <= 16367318;
srom_1(36255) <= 16525877;
srom_1(36256) <= 16646278;
srom_1(36257) <= 16727955;
srom_1(36258) <= 16770527;
srom_1(36259) <= 16773792;
srom_1(36260) <= 16737737;
srom_1(36261) <= 16662530;
srom_1(36262) <= 16548523;
srom_1(36263) <= 16396252;
srom_1(36264) <= 16206431;
srom_1(36265) <= 15979948;
srom_1(36266) <= 15717868;
srom_1(36267) <= 15421418;
srom_1(36268) <= 15091988;
srom_1(36269) <= 14731125;
srom_1(36270) <= 14340519;
srom_1(36271) <= 13922002;
srom_1(36272) <= 13477538;
srom_1(36273) <= 13009209;
srom_1(36274) <= 12519213;
srom_1(36275) <= 12009848;
srom_1(36276) <= 11483501;
srom_1(36277) <= 10942641;
srom_1(36278) <= 10389804;
srom_1(36279) <= 9827583;
srom_1(36280) <= 9258614;
srom_1(36281) <= 8685565;
srom_1(36282) <= 8111124;
srom_1(36283) <= 7537984;
srom_1(36284) <= 6968833;
srom_1(36285) <= 6406340;
srom_1(36286) <= 5853142;
srom_1(36287) <= 5311834;
srom_1(36288) <= 4784954;
srom_1(36289) <= 4274972;
srom_1(36290) <= 3784281;
srom_1(36291) <= 3315181;
srom_1(36292) <= 2869873;
srom_1(36293) <= 2450443;
srom_1(36294) <= 2058860;
srom_1(36295) <= 1696959;
srom_1(36296) <= 1366437;
srom_1(36297) <= 1068845;
srom_1(36298) <= 805577;
srom_1(36299) <= 577869;
srom_1(36300) <= 386788;
srom_1(36301) <= 233231;
srom_1(36302) <= 117917;
srom_1(36303) <= 41387;
srom_1(36304) <= 4000;
srom_1(36305) <= 5931;
srom_1(36306) <= 47172;
srom_1(36307) <= 127528;
srom_1(36308) <= 246623;
srom_1(36309) <= 403899;
srom_1(36310) <= 598618;
srom_1(36311) <= 829867;
srom_1(36312) <= 1096562;
srom_1(36313) <= 1397451;
srom_1(36314) <= 1731124;
srom_1(36315) <= 2096017;
srom_1(36316) <= 2490417;
srom_1(36317) <= 2912477;
srom_1(36318) <= 3360215;
srom_1(36319) <= 3831534;
srom_1(36320) <= 4324222;
srom_1(36321) <= 4835970;
srom_1(36322) <= 5364377;
srom_1(36323) <= 5906965;
srom_1(36324) <= 6461191;
srom_1(36325) <= 7024456;
srom_1(36326) <= 7594117;
srom_1(36327) <= 8167504;
srom_1(36328) <= 8741928;
srom_1(36329) <= 9314695;
srom_1(36330) <= 9883119;
srom_1(36331) <= 10444535;
srom_1(36332) <= 10996309;
srom_1(36333) <= 11535856;
srom_1(36334) <= 12060644;
srom_1(36335) <= 12568212;
srom_1(36336) <= 13056181;
srom_1(36337) <= 13522262;
srom_1(36338) <= 13964270;
srom_1(36339) <= 14380131;
srom_1(36340) <= 14767896;
srom_1(36341) <= 15125747;
srom_1(36342) <= 15452004;
srom_1(36343) <= 15745139;
srom_1(36344) <= 16003777;
srom_1(36345) <= 16226704;
srom_1(36346) <= 16412876;
srom_1(36347) <= 16561419;
srom_1(36348) <= 16671638;
srom_1(36349) <= 16743014;
srom_1(36350) <= 16775214;
srom_1(36351) <= 16768085;
srom_1(36352) <= 16721663;
srom_1(36353) <= 16636164;
srom_1(36354) <= 16511989;
srom_1(36355) <= 16349722;
srom_1(36356) <= 16150121;
srom_1(36357) <= 15914125;
srom_1(36358) <= 15642838;
srom_1(36359) <= 15337534;
srom_1(36360) <= 14999644;
srom_1(36361) <= 14630753;
srom_1(36362) <= 14232590;
srom_1(36363) <= 13807022;
srom_1(36364) <= 13356046;
srom_1(36365) <= 12881776;
srom_1(36366) <= 12386436;
srom_1(36367) <= 11872348;
srom_1(36368) <= 11341924;
srom_1(36369) <= 10797651;
srom_1(36370) <= 10242081;
srom_1(36371) <= 9677820;
srom_1(36372) <= 9107513;
srom_1(36373) <= 8533835;
srom_1(36374) <= 7959475;
srom_1(36375) <= 7387129;
srom_1(36376) <= 6819478;
srom_1(36377) <= 6259185;
srom_1(36378) <= 5708879;
srom_1(36379) <= 5171138;
srom_1(36380) <= 4648485;
srom_1(36381) <= 4143371;
srom_1(36382) <= 3658164;
srom_1(36383) <= 3195140;
srom_1(36384) <= 2756470;
srom_1(36385) <= 2344211;
srom_1(36386) <= 1960296;
srom_1(36387) <= 1606525;
srom_1(36388) <= 1284559;
srom_1(36389) <= 995905;
srom_1(36390) <= 741918;
srom_1(36391) <= 523790;
srom_1(36392) <= 342542;
srom_1(36393) <= 199025;
srom_1(36394) <= 93912;
srom_1(36395) <= 27695;
srom_1(36396) <= 686;
srom_1(36397) <= 13010;
srom_1(36398) <= 64610;
srom_1(36399) <= 155245;
srom_1(36400) <= 284489;
srom_1(36401) <= 451735;
srom_1(36402) <= 656200;
srom_1(36403) <= 896926;
srom_1(36404) <= 1172782;
srom_1(36405) <= 1482476;
srom_1(36406) <= 1824555;
srom_1(36407) <= 2197415;
srom_1(36408) <= 2599307;
srom_1(36409) <= 3028348;
srom_1(36410) <= 3482525;
srom_1(36411) <= 3959708;
srom_1(36412) <= 4457660;
srom_1(36413) <= 4974045;
srom_1(36414) <= 5506442;
srom_1(36415) <= 6052355;
srom_1(36416) <= 6609223;
srom_1(36417) <= 7174436;
srom_1(36418) <= 7745342;
srom_1(36419) <= 8319265;
srom_1(36420) <= 8893512;
srom_1(36421) <= 9465392;
srom_1(36422) <= 10032223;
srom_1(36423) <= 10591346;
srom_1(36424) <= 11140140;
srom_1(36425) <= 11676031;
srom_1(36426) <= 12196506;
srom_1(36427) <= 12699124;
srom_1(36428) <= 13181529;
srom_1(36429) <= 13641459;
srom_1(36430) <= 14076755;
srom_1(36431) <= 14485379;
srom_1(36432) <= 14865412;
srom_1(36433) <= 15215073;
srom_1(36434) <= 15532723;
srom_1(36435) <= 15816872;
srom_1(36436) <= 16066186;
srom_1(36437) <= 16279498;
srom_1(36438) <= 16455807;
srom_1(36439) <= 16594286;
srom_1(36440) <= 16694286;
srom_1(36441) <= 16755338;
srom_1(36442) <= 16777155;
srom_1(36443) <= 16759635;
srom_1(36444) <= 16702861;
srom_1(36445) <= 16607098;
srom_1(36446) <= 16472796;
srom_1(36447) <= 16300584;
srom_1(36448) <= 16091271;
srom_1(36449) <= 15845837;
srom_1(36450) <= 15565433;
srom_1(36451) <= 15251375;
srom_1(36452) <= 14905135;
srom_1(36453) <= 14528337;
srom_1(36454) <= 14122748;
srom_1(36455) <= 13690269;
srom_1(36456) <= 13232928;
srom_1(36457) <= 12752872;
srom_1(36458) <= 12252349;
srom_1(36459) <= 11733708;
srom_1(36460) <= 11199381;
srom_1(36461) <= 10651873;
srom_1(36462) <= 10093752;
srom_1(36463) <= 9527635;
srom_1(36464) <= 8956176;
srom_1(36465) <= 8382057;
srom_1(36466) <= 7807967;
srom_1(36467) <= 7236601;
srom_1(36468) <= 6670637;
srom_1(36469) <= 6112728;
srom_1(36470) <= 5565493;
srom_1(36471) <= 5031496;
srom_1(36472) <= 4513241;
srom_1(36473) <= 4013159;
srom_1(36474) <= 3533596;
srom_1(36475) <= 3076799;
srom_1(36476) <= 2644911;
srom_1(36477) <= 2239957;
srom_1(36478) <= 1863836;
srom_1(36479) <= 1518313;
srom_1(36480) <= 1205006;
srom_1(36481) <= 925386;
srom_1(36482) <= 680763;
srom_1(36483) <= 472285;
srom_1(36484) <= 300930;
srom_1(36485) <= 167500;
srom_1(36486) <= 72622;
srom_1(36487) <= 16741;
srom_1(36488) <= 118;
srom_1(36489) <= 22831;
srom_1(36490) <= 84775;
srom_1(36491) <= 185658;
srom_1(36492) <= 325007;
srom_1(36493) <= 502169;
srom_1(36494) <= 716314;
srom_1(36495) <= 966437;
srom_1(36496) <= 1251365;
srom_1(36497) <= 1569761;
srom_1(36498) <= 1920134;
srom_1(36499) <= 2300840;
srom_1(36500) <= 2710093;
srom_1(36501) <= 3145975;
srom_1(36502) <= 3606441;
srom_1(36503) <= 4089332;
srom_1(36504) <= 4592384;
srom_1(36505) <= 5113238;
srom_1(36506) <= 5649452;
srom_1(36507) <= 6198510;
srom_1(36508) <= 6757838;
srom_1(36509) <= 7324814;
srom_1(36510) <= 7896778;
srom_1(36511) <= 8471048;
srom_1(36512) <= 9044932;
srom_1(36513) <= 9615738;
srom_1(36514) <= 10180789;
srom_1(36515) <= 10737437;
srom_1(36516) <= 11283070;
srom_1(36517) <= 11815129;
srom_1(36518) <= 12331121;
srom_1(36519) <= 12828625;
srom_1(36520) <= 13305308;
srom_1(36521) <= 13758935;
srom_1(36522) <= 14187379;
srom_1(36523) <= 14588630;
srom_1(36524) <= 14960807;
srom_1(36525) <= 15302165;
srom_1(36526) <= 15611103;
srom_1(36527) <= 15886172;
srom_1(36528) <= 16126082;
srom_1(36529) <= 16329709;
srom_1(36530) <= 16496097;
srom_1(36531) <= 16624467;
srom_1(36532) <= 16714215;
srom_1(36533) <= 16764922;
srom_1(36534) <= 16776350;
srom_1(36535) <= 16748444;
srom_1(36536) <= 16681337;
srom_1(36537) <= 16575341;
srom_1(36538) <= 16430956;
srom_1(36539) <= 16248857;
srom_1(36540) <= 16029899;
srom_1(36541) <= 15775108;
srom_1(36542) <= 15485679;
srom_1(36543) <= 15162970;
srom_1(36544) <= 14808493;
srom_1(36545) <= 14423911;
srom_1(36546) <= 14011028;
srom_1(36547) <= 13571779;
srom_1(36548) <= 13108225;
srom_1(36549) <= 12622538;
srom_1(36550) <= 12116998;
srom_1(36551) <= 11593973;
srom_1(36552) <= 11055918;
srom_1(36553) <= 10505354;
srom_1(36554) <= 9944864;
srom_1(36555) <= 9377077;
srom_1(36556) <= 8804654;
srom_1(36557) <= 8230280;
srom_1(36558) <= 7656649;
srom_1(36559) <= 7086450;
srom_1(36560) <= 6522358;
srom_1(36561) <= 5967017;
srom_1(36562) <= 5423031;
srom_1(36563) <= 4892952;
srom_1(36564) <= 4379266;
srom_1(36565) <= 3884380;
srom_1(36566) <= 3410617;
srom_1(36567) <= 2960197;
srom_1(36568) <= 2535232;
srom_1(36569) <= 2137717;
srom_1(36570) <= 1769513;
srom_1(36571) <= 1432349;
srom_1(36572) <= 1127805;
srom_1(36573) <= 857310;
srom_1(36574) <= 622131;
srom_1(36575) <= 423373;
srom_1(36576) <= 261965;
srom_1(36577) <= 138667;
srom_1(36578) <= 54055;
srom_1(36579) <= 8527;
srom_1(36580) <= 2296;
srom_1(36581) <= 35391;
srom_1(36582) <= 107657;
srom_1(36583) <= 218756;
srom_1(36584) <= 368165;
srom_1(36585) <= 555186;
srom_1(36586) <= 778940;
srom_1(36587) <= 1038378;
srom_1(36588) <= 1332284;
srom_1(36589) <= 1659280;
srom_1(36590) <= 2017831;
srom_1(36591) <= 2406258;
srom_1(36592) <= 2822737;
srom_1(36593) <= 3265317;
srom_1(36594) <= 3731922;
srom_1(36595) <= 4220364;
srom_1(36596) <= 4728352;
srom_1(36597) <= 5253504;
srom_1(36598) <= 5793358;
srom_1(36599) <= 6345381;
srom_1(36600) <= 6906987;
srom_1(36601) <= 7475539;
srom_1(36602) <= 8048374;
srom_1(36603) <= 8622804;
srom_1(36604) <= 9196136;
srom_1(36605) <= 9765681;
srom_1(36606) <= 10328769;
srom_1(36607) <= 10882758;
srom_1(36608) <= 11425052;
srom_1(36609) <= 11953106;
srom_1(36610) <= 12464446;
srom_1(36611) <= 12956672;
srom_1(36612) <= 13427477;
srom_1(36613) <= 13874653;
srom_1(36614) <= 14296103;
srom_1(36615) <= 14689851;
srom_1(36616) <= 15054051;
srom_1(36617) <= 15386993;
srom_1(36618) <= 15687118;
srom_1(36619) <= 15953018;
srom_1(36620) <= 16183445;
srom_1(36621) <= 16377320;
srom_1(36622) <= 16533733;
srom_1(36623) <= 16651951;
srom_1(36624) <= 16731419;
srom_1(36625) <= 16771764;
srom_1(36626) <= 16772798;
srom_1(36627) <= 16734516;
srom_1(36628) <= 16657097;
srom_1(36629) <= 16540904;
srom_1(36630) <= 16386483;
srom_1(36631) <= 16194556;
srom_1(36632) <= 15966025;
srom_1(36633) <= 15701961;
srom_1(36634) <= 15403601;
srom_1(36635) <= 15072346;
srom_1(36636) <= 14709749;
srom_1(36637) <= 14317510;
srom_1(36638) <= 13897468;
srom_1(36639) <= 13451593;
srom_1(36640) <= 12981976;
srom_1(36641) <= 12490819;
srom_1(36642) <= 11980425;
srom_1(36643) <= 11453189;
srom_1(36644) <= 10911581;
srom_1(36645) <= 10358142;
srom_1(36646) <= 9795467;
srom_1(36647) <= 9226195;
srom_1(36648) <= 8652996;
srom_1(36649) <= 8078556;
srom_1(36650) <= 7505571;
srom_1(36651) <= 6936726;
srom_1(36652) <= 6374690;
srom_1(36653) <= 5822097;
srom_1(36654) <= 5281540;
srom_1(36655) <= 4755553;
srom_1(36656) <= 4246603;
srom_1(36657) <= 3757076;
srom_1(36658) <= 3289268;
srom_1(36659) <= 2845372;
srom_1(36660) <= 2427470;
srom_1(36661) <= 2037523;
srom_1(36662) <= 1677357;
srom_1(36663) <= 1348663;
srom_1(36664) <= 1052982;
srom_1(36665) <= 791700;
srom_1(36666) <= 566042;
srom_1(36667) <= 377068;
srom_1(36668) <= 225662;
srom_1(36669) <= 112534;
srom_1(36670) <= 38217;
srom_1(36671) <= 3057;
srom_1(36672) <= 7220;
srom_1(36673) <= 50686;
srom_1(36674) <= 133251;
srom_1(36675) <= 254529;
srom_1(36676) <= 413950;
srom_1(36677) <= 610767;
srom_1(36678) <= 844057;
srom_1(36679) <= 1112725;
srom_1(36680) <= 1415514;
srom_1(36681) <= 1751001;
srom_1(36682) <= 2117614;
srom_1(36683) <= 2513634;
srom_1(36684) <= 2937204;
srom_1(36685) <= 3386337;
srom_1(36686) <= 3858928;
srom_1(36687) <= 4352760;
srom_1(36688) <= 4865518;
srom_1(36689) <= 5394796;
srom_1(36690) <= 5938113;
srom_1(36691) <= 6492922;
srom_1(36692) <= 7056620;
srom_1(36693) <= 7626564;
srom_1(36694) <= 8200082;
srom_1(36695) <= 8774484;
srom_1(36696) <= 9347076;
srom_1(36697) <= 9915174;
srom_1(36698) <= 10476113;
srom_1(36699) <= 11027263;
srom_1(36700) <= 11566039;
srom_1(36701) <= 12089916;
srom_1(36702) <= 12596436;
srom_1(36703) <= 13083223;
srom_1(36704) <= 13547996;
srom_1(36705) <= 13988575;
srom_1(36706) <= 14402894;
srom_1(36707) <= 14789010;
srom_1(36708) <= 15145112;
srom_1(36709) <= 15469530;
srom_1(36710) <= 15760744;
srom_1(36711) <= 16017387;
srom_1(36712) <= 16238256;
srom_1(36713) <= 16422315;
srom_1(36714) <= 16568702;
srom_1(36715) <= 16676729;
srom_1(36716) <= 16745891;
srom_1(36717) <= 16775862;
srom_1(36718) <= 16766502;
srom_1(36719) <= 16717856;
srom_1(36720) <= 16630151;
srom_1(36721) <= 16503799;
srom_1(36722) <= 16339391;
srom_1(36723) <= 16137700;
srom_1(36724) <= 15899670;
srom_1(36725) <= 15626419;
srom_1(36726) <= 15319227;
srom_1(36727) <= 14979535;
srom_1(36728) <= 14608936;
srom_1(36729) <= 14209167;
srom_1(36730) <= 13782104;
srom_1(36731) <= 13329749;
srom_1(36732) <= 12854223;
srom_1(36733) <= 12357757;
srom_1(36734) <= 11842677;
srom_1(36735) <= 11311401;
srom_1(36736) <= 10766418;
srom_1(36737) <= 10210285;
srom_1(36738) <= 9645610;
srom_1(36739) <= 9075040;
srom_1(36740) <= 8501251;
srom_1(36741) <= 7926934;
srom_1(36742) <= 7354781;
srom_1(36743) <= 6787477;
srom_1(36744) <= 6227681;
srom_1(36745) <= 5678019;
srom_1(36746) <= 5141067;
srom_1(36747) <= 4619344;
srom_1(36748) <= 4115296;
srom_1(36749) <= 3631288;
srom_1(36750) <= 3169588;
srom_1(36751) <= 2732362;
srom_1(36752) <= 2321660;
srom_1(36753) <= 1939408;
srom_1(36754) <= 1587398;
srom_1(36755) <= 1267282;
srom_1(36756) <= 980560;
srom_1(36757) <= 728577;
srom_1(36758) <= 512514;
srom_1(36759) <= 333385;
srom_1(36760) <= 192030;
srom_1(36761) <= 89112;
srom_1(36762) <= 25112;
srom_1(36763) <= 332;
srom_1(36764) <= 14887;
srom_1(36765) <= 68710;
srom_1(36766) <= 161548;
srom_1(36767) <= 292965;
srom_1(36768) <= 462345;
srom_1(36769) <= 668894;
srom_1(36770) <= 911643;
srom_1(36771) <= 1189455;
srom_1(36772) <= 1501026;
srom_1(36773) <= 1844895;
srom_1(36774) <= 2219450;
srom_1(36775) <= 2622934;
srom_1(36776) <= 3053456;
srom_1(36777) <= 3508995;
srom_1(36778) <= 3987417;
srom_1(36779) <= 4486478;
srom_1(36780) <= 5003837;
srom_1(36781) <= 5537068;
srom_1(36782) <= 6083671;
srom_1(36783) <= 6641083;
srom_1(36784) <= 7206690;
srom_1(36785) <= 7777839;
srom_1(36786) <= 8351852;
srom_1(36787) <= 8926037;
srom_1(36788) <= 9497702;
srom_1(36789) <= 10064167;
srom_1(36790) <= 10622774;
srom_1(36791) <= 11170904;
srom_1(36792) <= 11705987;
srom_1(36793) <= 12225514;
srom_1(36794) <= 12727048;
srom_1(36795) <= 13208238;
srom_1(36796) <= 13666827;
srom_1(36797) <= 14100664;
srom_1(36798) <= 14507716;
srom_1(36799) <= 14886073;
srom_1(36800) <= 15233961;
srom_1(36801) <= 15549749;
srom_1(36802) <= 15831956;
srom_1(36803) <= 16079258;
srom_1(36804) <= 16290497;
srom_1(36805) <= 16464680;
srom_1(36806) <= 16600993;
srom_1(36807) <= 16698794;
srom_1(36808) <= 16757626;
srom_1(36809) <= 16777213;
srom_1(36810) <= 16757463;
srom_1(36811) <= 16698469;
srom_1(36812) <= 16600507;
srom_1(36813) <= 16464036;
srom_1(36814) <= 16289697;
srom_1(36815) <= 16078306;
srom_1(36816) <= 15830857;
srom_1(36817) <= 15548508;
srom_1(36818) <= 15232583;
srom_1(36819) <= 14884565;
srom_1(36820) <= 14506086;
srom_1(36821) <= 14098919;
srom_1(36822) <= 13664974;
srom_1(36823) <= 13206287;
srom_1(36824) <= 12725008;
srom_1(36825) <= 12223395;
srom_1(36826) <= 11703798;
srom_1(36827) <= 11168656;
srom_1(36828) <= 10620477;
srom_1(36829) <= 10061832;
srom_1(36830) <= 9495340;
srom_1(36831) <= 8923659;
srom_1(36832) <= 8349469;
srom_1(36833) <= 7775462;
srom_1(36834) <= 7204331;
srom_1(36835) <= 6638753;
srom_1(36836) <= 6081380;
srom_1(36837) <= 5534827;
srom_1(36838) <= 5001657;
srom_1(36839) <= 4484368;
srom_1(36840) <= 3985389;
srom_1(36841) <= 3507057;
srom_1(36842) <= 3051617;
srom_1(36843) <= 2621204;
srom_1(36844) <= 2217836;
srom_1(36845) <= 1843404;
srom_1(36846) <= 1499666;
srom_1(36847) <= 1188232;
srom_1(36848) <= 910563;
srom_1(36849) <= 667962;
srom_1(36850) <= 461565;
srom_1(36851) <= 292341;
srom_1(36852) <= 161082;
srom_1(36853) <= 68406;
srom_1(36854) <= 14746;
srom_1(36855) <= 354;
srom_1(36856) <= 25297;
srom_1(36857) <= 89458;
srom_1(36858) <= 192538;
srom_1(36859) <= 334051;
srom_1(36860) <= 513335;
srom_1(36861) <= 729549;
srom_1(36862) <= 981678;
srom_1(36863) <= 1268542;
srom_1(36864) <= 1588793;
srom_1(36865) <= 1940932;
srom_1(36866) <= 2323306;
srom_1(36867) <= 2734122;
srom_1(36868) <= 3171454;
srom_1(36869) <= 3633251;
srom_1(36870) <= 4117347;
srom_1(36871) <= 4621473;
srom_1(36872) <= 5143264;
srom_1(36873) <= 5680274;
srom_1(36874) <= 6229984;
srom_1(36875) <= 6789816;
srom_1(36876) <= 7357146;
srom_1(36877) <= 7929313;
srom_1(36878) <= 8503633;
srom_1(36879) <= 9077415;
srom_1(36880) <= 9647966;
srom_1(36881) <= 10212611;
srom_1(36882) <= 10768703;
srom_1(36883) <= 11313634;
srom_1(36884) <= 11844849;
srom_1(36885) <= 12359856;
srom_1(36886) <= 12856240;
srom_1(36887) <= 13331674;
srom_1(36888) <= 13783929;
srom_1(36889) <= 14210883;
srom_1(36890) <= 14610534;
srom_1(36891) <= 14981009;
srom_1(36892) <= 15320569;
srom_1(36893) <= 15627623;
srom_1(36894) <= 15900731;
srom_1(36895) <= 16138612;
srom_1(36896) <= 16340151;
srom_1(36897) <= 16504402;
srom_1(36898) <= 16630595;
srom_1(36899) <= 16718139;
srom_1(36900) <= 16766622;
srom_1(36901) <= 16775819;
srom_1(36902) <= 16745684;
srom_1(36903) <= 16676361;
srom_1(36904) <= 16568174;
srom_1(36905) <= 16421629;
srom_1(36906) <= 16237415;
srom_1(36907) <= 16016395;
srom_1(36908) <= 15759606;
srom_1(36909) <= 15468252;
srom_1(36910) <= 15143699;
srom_1(36911) <= 14787469;
srom_1(36912) <= 14401233;
srom_1(36913) <= 13986801;
srom_1(36914) <= 13546117;
srom_1(36915) <= 13081248;
srom_1(36916) <= 12594374;
srom_1(36917) <= 12087777;
srom_1(36918) <= 11563834;
srom_1(36919) <= 11025001;
srom_1(36920) <= 10473805;
srom_1(36921) <= 9912831;
srom_1(36922) <= 9344709;
srom_1(36923) <= 8772103;
srom_1(36924) <= 8197700;
srom_1(36925) <= 7624191;
srom_1(36926) <= 7054267;
srom_1(36927) <= 6490601;
srom_1(36928) <= 5935834;
srom_1(36929) <= 5392570;
srom_1(36930) <= 4863355;
srom_1(36931) <= 4350671;
srom_1(36932) <= 3856923;
srom_1(36933) <= 3384425;
srom_1(36934) <= 2935393;
srom_1(36935) <= 2511933;
srom_1(36936) <= 2116032;
srom_1(36937) <= 1749544;
srom_1(36938) <= 1414189;
srom_1(36939) <= 1111540;
srom_1(36940) <= 843015;
srom_1(36941) <= 609874;
srom_1(36942) <= 413211;
srom_1(36943) <= 253946;
srom_1(36944) <= 132828;
srom_1(36945) <= 50424;
srom_1(36946) <= 7121;
srom_1(36947) <= 3121;
srom_1(36948) <= 38444;
srom_1(36949) <= 112924;
srom_1(36950) <= 226211;
srom_1(36951) <= 377774;
srom_1(36952) <= 566903;
srom_1(36953) <= 792711;
srom_1(36954) <= 1054138;
srom_1(36955) <= 1349959;
srom_1(36956) <= 1678787;
srom_1(36957) <= 2039080;
srom_1(36958) <= 2429147;
srom_1(36959) <= 2847161;
srom_1(36960) <= 3291160;
srom_1(36961) <= 3759063;
srom_1(36962) <= 4248675;
srom_1(36963) <= 4757701;
srom_1(36964) <= 5283754;
srom_1(36965) <= 5824366;
srom_1(36966) <= 6377003;
srom_1(36967) <= 6939073;
srom_1(36968) <= 7507940;
srom_1(36969) <= 8080938;
srom_1(36970) <= 8655377;
srom_1(36971) <= 9228566;
srom_1(36972) <= 9797816;
srom_1(36973) <= 10360458;
srom_1(36974) <= 10913853;
srom_1(36975) <= 11455407;
srom_1(36976) <= 11982579;
srom_1(36977) <= 12492897;
srom_1(36978) <= 12983970;
srom_1(36979) <= 13453493;
srom_1(36980) <= 13899265;
srom_1(36981) <= 14319195;
srom_1(36982) <= 14711315;
srom_1(36983) <= 15073786;
srom_1(36984) <= 15404908;
srom_1(36985) <= 15703127;
srom_1(36986) <= 15967047;
srom_1(36987) <= 16195429;
srom_1(36988) <= 16387201;
srom_1(36989) <= 16541466;
srom_1(36990) <= 16657499;
srom_1(36991) <= 16734756;
srom_1(36992) <= 16772875;
srom_1(36993) <= 16771678;
srom_1(36994) <= 16731170;
srom_1(36995) <= 16651540;
srom_1(36996) <= 16533163;
srom_1(36997) <= 16376593;
srom_1(36998) <= 16182564;
srom_1(36999) <= 15951987;
srom_1(37000) <= 15685943;
srom_1(37001) <= 15385679;
srom_1(37002) <= 15052603;
srom_1(37003) <= 14688278;
srom_1(37004) <= 14294411;
srom_1(37005) <= 13872850;
srom_1(37006) <= 13425572;
srom_1(37007) <= 12954673;
srom_1(37008) <= 12462363;
srom_1(37009) <= 11950949;
srom_1(37010) <= 11422830;
srom_1(37011) <= 10880483;
srom_1(37012) <= 10326450;
srom_1(37013) <= 9763331;
srom_1(37014) <= 9193764;
srom_1(37015) <= 8620422;
srom_1(37016) <= 8045993;
srom_1(37017) <= 7473171;
srom_1(37018) <= 6904641;
srom_1(37019) <= 6343070;
srom_1(37020) <= 5791092;
srom_1(37021) <= 5251294;
srom_1(37022) <= 4726208;
srom_1(37023) <= 4218296;
srom_1(37024) <= 3729940;
srom_1(37025) <= 3263431;
srom_1(37026) <= 2820955;
srom_1(37027) <= 2404587;
srom_1(37028) <= 2016281;
srom_1(37029) <= 1657857;
srom_1(37030) <= 1330996;
srom_1(37031) <= 1037230;
srom_1(37032) <= 777937;
srom_1(37033) <= 554334;
srom_1(37034) <= 367468;
srom_1(37035) <= 218215;
srom_1(37036) <= 107277;
srom_1(37037) <= 35173;
srom_1(37038) <= 2240;
srom_1(37039) <= 8635;
srom_1(37040) <= 54325;
srom_1(37041) <= 139099;
srom_1(37042) <= 262557;
srom_1(37043) <= 424120;
srom_1(37044) <= 623032;
srom_1(37045) <= 858360;
srom_1(37046) <= 1128999;
srom_1(37047) <= 1433681;
srom_1(37048) <= 1770977;
srom_1(37049) <= 2139306;
srom_1(37050) <= 2536940;
srom_1(37051) <= 2962014;
srom_1(37052) <= 3412535;
srom_1(37053) <= 3886391;
srom_1(37054) <= 4381359;
srom_1(37055) <= 4895118;
srom_1(37056) <= 5425260;
srom_1(37057) <= 5969298;
srom_1(37058) <= 6524681;
srom_1(37059) <= 7088804;
srom_1(37060) <= 7659023;
srom_1(37061) <= 8232663;
srom_1(37062) <= 8807034;
srom_1(37063) <= 9379443;
srom_1(37064) <= 9947206;
srom_1(37065) <= 10507660;
srom_1(37066) <= 11058177;
srom_1(37067) <= 11596175;
srom_1(37068) <= 12119132;
srom_1(37069) <= 12624595;
srom_1(37070) <= 13110195;
srom_1(37071) <= 13573653;
srom_1(37072) <= 14012796;
srom_1(37073) <= 14425566;
srom_1(37074) <= 14810027;
srom_1(37075) <= 15164375;
srom_1(37076) <= 15486949;
srom_1(37077) <= 15776237;
srom_1(37078) <= 16030882;
srom_1(37079) <= 16249689;
srom_1(37080) <= 16431633;
srom_1(37081) <= 16575861;
srom_1(37082) <= 16681695;
srom_1(37083) <= 16748641;
srom_1(37084) <= 16776383;
srom_1(37085) <= 16764793;
srom_1(37086) <= 16713923;
srom_1(37087) <= 16624014;
srom_1(37088) <= 16495485;
srom_1(37089) <= 16328941;
srom_1(37090) <= 16125162;
srom_1(37091) <= 15885103;
srom_1(37092) <= 15609891;
srom_1(37093) <= 15300815;
srom_1(37094) <= 14959326;
srom_1(37095) <= 14587025;
srom_1(37096) <= 14185657;
srom_1(37097) <= 13757104;
srom_1(37098) <= 13303377;
srom_1(37099) <= 12826603;
srom_1(37100) <= 12329018;
srom_1(37101) <= 11812954;
srom_1(37102) <= 11280833;
srom_1(37103) <= 10735149;
srom_1(37104) <= 10178461;
srom_1(37105) <= 9613380;
srom_1(37106) <= 9042556;
srom_1(37107) <= 8468665;
srom_1(37108) <= 7894399;
srom_1(37109) <= 7322450;
srom_1(37110) <= 6755501;
srom_1(37111) <= 6196210;
srom_1(37112) <= 5647199;
srom_1(37113) <= 5111045;
srom_1(37114) <= 4590260;
srom_1(37115) <= 4087286;
srom_1(37116) <= 3604483;
srom_1(37117) <= 3144115;
srom_1(37118) <= 2708339;
srom_1(37119) <= 2299200;
srom_1(37120) <= 1918617;
srom_1(37121) <= 1568374;
srom_1(37122) <= 1250113;
srom_1(37123) <= 965327;
srom_1(37124) <= 715351;
srom_1(37125) <= 501358;
srom_1(37126) <= 324350;
srom_1(37127) <= 185159;
srom_1(37128) <= 84437;
srom_1(37129) <= 22656;
srom_1(37130) <= 105;
srom_1(37131) <= 16891;
srom_1(37132) <= 72935;
srom_1(37133) <= 167974;
srom_1(37134) <= 301563;
srom_1(37135) <= 473074;
srom_1(37136) <= 681704;
srom_1(37137) <= 926474;
srom_1(37138) <= 1206237;
srom_1(37139) <= 1519680;
srom_1(37140) <= 1865334;
srom_1(37141) <= 2241578;
srom_1(37142) <= 2646648;
srom_1(37143) <= 3078643;
srom_1(37144) <= 3535539;
srom_1(37145) <= 4015193;
srom_1(37146) <= 4515355;
srom_1(37147) <= 5033679;
srom_1(37148) <= 5567737;
srom_1(37149) <= 6115022;
srom_1(37150) <= 6672969;
srom_1(37151) <= 7238961;
srom_1(37152) <= 7810345;
srom_1(37153) <= 8384439;
srom_1(37154) <= 8958554;
srom_1(37155) <= 9529996;
srom_1(37156) <= 10096085;
srom_1(37157) <= 10654168;
srom_1(37158) <= 11201626;
srom_1(37159) <= 11735893;
srom_1(37160) <= 12254464;
srom_1(37161) <= 12754906;
srom_1(37162) <= 13234874;
srom_1(37163) <= 13692115;
srom_1(37164) <= 14124487;
srom_1(37165) <= 14529961;
srom_1(37166) <= 14906636;
srom_1(37167) <= 15252745;
srom_1(37168) <= 15566667;
srom_1(37169) <= 15846928;
srom_1(37170) <= 16092214;
srom_1(37171) <= 16301376;
srom_1(37172) <= 16473432;
srom_1(37173) <= 16607575;
srom_1(37174) <= 16703177;
srom_1(37175) <= 16759789;
srom_1(37176) <= 16777145;
srom_1(37177) <= 16755165;
srom_1(37178) <= 16693951;
srom_1(37179) <= 16593791;
srom_1(37180) <= 16455154;
srom_1(37181) <= 16278689;
srom_1(37182) <= 16065226;
srom_1(37183) <= 15815764;
srom_1(37184) <= 15531474;
srom_1(37185) <= 15213688;
srom_1(37186) <= 14863897;
srom_1(37187) <= 14483742;
srom_1(37188) <= 14075004;
srom_1(37189) <= 13639600;
srom_1(37190) <= 13179573;
srom_1(37191) <= 12697080;
srom_1(37192) <= 12194382;
srom_1(37193) <= 11673838;
srom_1(37194) <= 11137889;
srom_1(37195) <= 10589047;
srom_1(37196) <= 10029886;
srom_1(37197) <= 9463029;
srom_1(37198) <= 8891134;
srom_1(37199) <= 8316882;
srom_1(37200) <= 7742966;
srom_1(37201) <= 7172078;
srom_1(37202) <= 6606895;
srom_1(37203) <= 6050067;
srom_1(37204) <= 5504205;
srom_1(37205) <= 4971869;
srom_1(37206) <= 4455555;
srom_1(37207) <= 3957684;
srom_1(37208) <= 3480592;
srom_1(37209) <= 3026515;
srom_1(37210) <= 2597583;
srom_1(37211) <= 2195807;
srom_1(37212) <= 1823071;
srom_1(37213) <= 1481123;
srom_1(37214) <= 1171567;
srom_1(37215) <= 895854;
srom_1(37216) <= 655277;
srom_1(37217) <= 450964;
srom_1(37218) <= 283874;
srom_1(37219) <= 154789;
srom_1(37220) <= 64316;
srom_1(37221) <= 12878;
srom_1(37222) <= 716;
srom_1(37223) <= 27889;
srom_1(37224) <= 94268;
srom_1(37225) <= 199541;
srom_1(37226) <= 343216;
srom_1(37227) <= 524619;
srom_1(37228) <= 742899;
srom_1(37229) <= 997032;
srom_1(37230) <= 1285826;
srom_1(37231) <= 1607928;
srom_1(37232) <= 1961827;
srom_1(37233) <= 2345863;
srom_1(37234) <= 2758236;
srom_1(37235) <= 3197012;
srom_1(37236) <= 3660132;
srom_1(37237) <= 4145426;
srom_1(37238) <= 4650618;
srom_1(37239) <= 5173339;
srom_1(37240) <= 5711137;
srom_1(37241) <= 6261490;
srom_1(37242) <= 6821819;
srom_1(37243) <= 7389494;
srom_1(37244) <= 7961855;
srom_1(37245) <= 8536217;
srom_1(37246) <= 9109887;
srom_1(37247) <= 9680174;
srom_1(37248) <= 10244405;
srom_1(37249) <= 10799934;
srom_1(37250) <= 11344155;
srom_1(37251) <= 11874516;
srom_1(37252) <= 12388530;
srom_1(37253) <= 12883788;
srom_1(37254) <= 13357966;
srom_1(37255) <= 13808841;
srom_1(37256) <= 14234299;
srom_1(37257) <= 14632344;
srom_1(37258) <= 15001111;
srom_1(37259) <= 15338869;
srom_1(37260) <= 15644034;
srom_1(37261) <= 15915177;
srom_1(37262) <= 16151025;
srom_1(37263) <= 16350472;
srom_1(37264) <= 16512584;
srom_1(37265) <= 16636599;
srom_1(37266) <= 16721936;
srom_1(37267) <= 16768196;
srom_1(37268) <= 16775161;
srom_1(37269) <= 16742799;
srom_1(37270) <= 16671261;
srom_1(37271) <= 16560882;
srom_1(37272) <= 16412181;
srom_1(37273) <= 16225855;
srom_1(37274) <= 16002777;
srom_1(37275) <= 15743994;
srom_1(37276) <= 15450719;
srom_1(37277) <= 15124327;
srom_1(37278) <= 14766349;
srom_1(37279) <= 14378463;
srom_1(37280) <= 13962489;
srom_1(37281) <= 13520378;
srom_1(37282) <= 13054201;
srom_1(37283) <= 12566146;
srom_1(37284) <= 12058501;
srom_1(37285) <= 11533647;
srom_1(37286) <= 10994045;
srom_1(37287) <= 10442224;
srom_1(37288) <= 9880774;
srom_1(37289) <= 9312326;
srom_1(37290) <= 8739547;
srom_1(37291) <= 8165122;
srom_1(37292) <= 7591745;
srom_1(37293) <= 7022105;
srom_1(37294) <= 6458872;
srom_1(37295) <= 5904689;
srom_1(37296) <= 5362154;
srom_1(37297) <= 4833811;
srom_1(37298) <= 4322138;
srom_1(37299) <= 3829533;
srom_1(37300) <= 3358308;
srom_1(37301) <= 2910672;
srom_1(37302) <= 2488723;
srom_1(37303) <= 2094441;
srom_1(37304) <= 1729675;
srom_1(37305) <= 1396134;
srom_1(37306) <= 1095384;
srom_1(37307) <= 828834;
srom_1(37308) <= 597735;
srom_1(37309) <= 403169;
srom_1(37310) <= 246050;
srom_1(37311) <= 127114;
srom_1(37312) <= 46920;
srom_1(37313) <= 5842;
srom_1(37314) <= 4074;
srom_1(37315) <= 41624;
srom_1(37316) <= 118315;
srom_1(37317) <= 233789;
srom_1(37318) <= 387504;
srom_1(37319) <= 578739;
srom_1(37320) <= 806596;
srom_1(37321) <= 1070009;
srom_1(37322) <= 1367741;
srom_1(37323) <= 1698396;
srom_1(37324) <= 2060424;
srom_1(37325) <= 2452126;
srom_1(37326) <= 2871668;
srom_1(37327) <= 3317079;
srom_1(37328) <= 3786273;
srom_1(37329) <= 4277049;
srom_1(37330) <= 4787106;
srom_1(37331) <= 5314051;
srom_1(37332) <= 5855413;
srom_1(37333) <= 6408655;
srom_1(37334) <= 6971182;
srom_1(37335) <= 7540355;
srom_1(37336) <= 8113506;
srom_1(37337) <= 8687947;
srom_1(37338) <= 9260984;
srom_1(37339) <= 9829930;
srom_1(37340) <= 10392118;
srom_1(37341) <= 10944910;
srom_1(37342) <= 11485715;
srom_1(37343) <= 12011997;
srom_1(37344) <= 12521287;
srom_1(37345) <= 13011198;
srom_1(37346) <= 13479432;
srom_1(37347) <= 13923793;
srom_1(37348) <= 14342198;
srom_1(37349) <= 14732684;
srom_1(37350) <= 15093421;
srom_1(37351) <= 15422716;
srom_1(37352) <= 15719027;
srom_1(37353) <= 15980962;
srom_1(37354) <= 16207294;
srom_1(37355) <= 16396962;
srom_1(37356) <= 16549076;
srom_1(37357) <= 16662922;
srom_1(37358) <= 16737968;
srom_1(37359) <= 16773860;
srom_1(37360) <= 16770431;
srom_1(37361) <= 16727697;
srom_1(37362) <= 16645858;
srom_1(37363) <= 16525298;
srom_1(37364) <= 16366582;
srom_1(37365) <= 16170455;
srom_1(37366) <= 15937835;
srom_1(37367) <= 15669815;
srom_1(37368) <= 15367651;
srom_1(37369) <= 15032760;
srom_1(37370) <= 14666712;
srom_1(37371) <= 14271224;
srom_1(37372) <= 13848150;
srom_1(37373) <= 13399475;
srom_1(37374) <= 12927301;
srom_1(37375) <= 12433845;
srom_1(37376) <= 11921419;
srom_1(37377) <= 11392426;
srom_1(37378) <= 10849347;
srom_1(37379) <= 10294729;
srom_1(37380) <= 9731173;
srom_1(37381) <= 9161321;
srom_1(37382) <= 8587845;
srom_1(37383) <= 8013435;
srom_1(37384) <= 7440785;
srom_1(37385) <= 6872579;
srom_1(37386) <= 6311482;
srom_1(37387) <= 5760125;
srom_1(37388) <= 5221095;
srom_1(37389) <= 4696918;
srom_1(37390) <= 4190052;
srom_1(37391) <= 3702875;
srom_1(37392) <= 3237671;
srom_1(37393) <= 2796622;
srom_1(37394) <= 2381795;
srom_1(37395) <= 1995136;
srom_1(37396) <= 1638459;
srom_1(37397) <= 1313435;
srom_1(37398) <= 1021589;
srom_1(37399) <= 764289;
srom_1(37400) <= 542743;
srom_1(37401) <= 357989;
srom_1(37402) <= 210892;
srom_1(37403) <= 102144;
srom_1(37404) <= 32255;
srom_1(37405) <= 1550;
srom_1(37406) <= 10176;
srom_1(37407) <= 58091;
srom_1(37408) <= 145071;
srom_1(37409) <= 270707;
srom_1(37410) <= 434411;
srom_1(37411) <= 635415;
srom_1(37412) <= 872777;
srom_1(37413) <= 1145382;
srom_1(37414) <= 1451954;
srom_1(37415) <= 1791054;
srom_1(37416) <= 2161092;
srom_1(37417) <= 2560333;
srom_1(37418) <= 2986905;
srom_1(37419) <= 3438808;
srom_1(37420) <= 3913921;
srom_1(37421) <= 4410018;
srom_1(37422) <= 4924772;
srom_1(37423) <= 5455769;
srom_1(37424) <= 6000519;
srom_1(37425) <= 6556468;
srom_1(37426) <= 7121008;
srom_1(37427) <= 7691493;
srom_1(37428) <= 8265246;
srom_1(37429) <= 8839578;
srom_1(37430) <= 9411795;
srom_1(37431) <= 9979214;
srom_1(37432) <= 10539175;
srom_1(37433) <= 11089050;
srom_1(37434) <= 11626262;
srom_1(37435) <= 12148292;
srom_1(37436) <= 12652691;
srom_1(37437) <= 13137094;
srom_1(37438) <= 13599231;
srom_1(37439) <= 14036932;
srom_1(37440) <= 14448147;
srom_1(37441) <= 14830947;
srom_1(37442) <= 15183536;
srom_1(37443) <= 15504261;
srom_1(37444) <= 15791619;
srom_1(37445) <= 16044261;
srom_1(37446) <= 16261004;
srom_1(37447) <= 16440830;
srom_1(37448) <= 16582896;
srom_1(37449) <= 16686537;
srom_1(37450) <= 16751265;
srom_1(37451) <= 16776779;
srom_1(37452) <= 16762957;
srom_1(37453) <= 16709865;
srom_1(37454) <= 16617752;
srom_1(37455) <= 16487049;
srom_1(37456) <= 16318371;
srom_1(37457) <= 16112506;
srom_1(37458) <= 15870422;
srom_1(37459) <= 15593253;
srom_1(37460) <= 15282299;
srom_1(37461) <= 14939018;
srom_1(37462) <= 14565020;
srom_1(37463) <= 14162059;
srom_1(37464) <= 13732023;
srom_1(37465) <= 13276931;
srom_1(37466) <= 12798916;
srom_1(37467) <= 12300219;
srom_1(37468) <= 11783179;
srom_1(37469) <= 11250221;
srom_1(37470) <= 10703844;
srom_1(37471) <= 10146610;
srom_1(37472) <= 9581133;
srom_1(37473) <= 9010062;
srom_1(37474) <= 8436078;
srom_1(37475) <= 7861871;
srom_1(37476) <= 7290134;
srom_1(37477) <= 6723549;
srom_1(37478) <= 6164771;
srom_1(37479) <= 5616422;
srom_1(37480) <= 5081072;
srom_1(37481) <= 4561233;
srom_1(37482) <= 4059341;
srom_1(37483) <= 3577751;
srom_1(37484) <= 3118720;
srom_1(37485) <= 2684402;
srom_1(37486) <= 2276833;
srom_1(37487) <= 1897924;
srom_1(37488) <= 1549452;
srom_1(37489) <= 1233051;
srom_1(37490) <= 950205;
srom_1(37491) <= 702241;
srom_1(37492) <= 490320;
srom_1(37493) <= 315437;
srom_1(37494) <= 178412;
srom_1(37495) <= 79888;
srom_1(37496) <= 20325;
srom_1(37497) <= 5;
srom_1(37498) <= 19022;
srom_1(37499) <= 77286;
srom_1(37500) <= 174525;
srom_1(37501) <= 310283;
srom_1(37502) <= 483923;
srom_1(37503) <= 694630;
srom_1(37504) <= 941417;
srom_1(37505) <= 1223127;
srom_1(37506) <= 1538438;
srom_1(37507) <= 1885872;
srom_1(37508) <= 2263799;
srom_1(37509) <= 2670448;
srom_1(37510) <= 3103911;
srom_1(37511) <= 3562156;
srom_1(37512) <= 4043034;
srom_1(37513) <= 4544290;
srom_1(37514) <= 5063573;
srom_1(37515) <= 5598448;
srom_1(37516) <= 6146407;
srom_1(37517) <= 6704881;
srom_1(37518) <= 7271250;
srom_1(37519) <= 7842859;
srom_1(37520) <= 8417027;
srom_1(37521) <= 8991062;
srom_1(37522) <= 9562272;
srom_1(37523) <= 10127978;
srom_1(37524) <= 10685527;
srom_1(37525) <= 11232306;
srom_1(37526) <= 11765749;
srom_1(37527) <= 12283356;
srom_1(37528) <= 12782699;
srom_1(37529) <= 13261436;
srom_1(37530) <= 13717323;
srom_1(37531) <= 14148222;
srom_1(37532) <= 14552113;
srom_1(37533) <= 14927100;
srom_1(37534) <= 15271426;
srom_1(37535) <= 15583476;
srom_1(37536) <= 15861787;
srom_1(37537) <= 16105054;
srom_1(37538) <= 16312136;
srom_1(37539) <= 16482061;
srom_1(37540) <= 16614034;
srom_1(37541) <= 16707434;
srom_1(37542) <= 16761825;
srom_1(37543) <= 16776951;
srom_1(37544) <= 16752741;
srom_1(37545) <= 16689309;
srom_1(37546) <= 16586952;
srom_1(37547) <= 16446150;
srom_1(37548) <= 16267563;
srom_1(37549) <= 16052030;
srom_1(37550) <= 15800559;
srom_1(37551) <= 15514332;
srom_1(37552) <= 15194690;
srom_1(37553) <= 14843132;
srom_1(37554) <= 14461306;
srom_1(37555) <= 14051003;
srom_1(37556) <= 13614147;
srom_1(37557) <= 13152787;
srom_1(37558) <= 12669086;
srom_1(37559) <= 12165313;
srom_1(37560) <= 11643829;
srom_1(37561) <= 11107080;
srom_1(37562) <= 10557584;
srom_1(37563) <= 9997916;
srom_1(37564) <= 9430702;
srom_1(37565) <= 8858601;
srom_1(37566) <= 8284296;
srom_1(37567) <= 7710480;
srom_1(37568) <= 7139844;
srom_1(37569) <= 6575064;
srom_1(37570) <= 6018788;
srom_1(37571) <= 5473626;
srom_1(37572) <= 4942132;
srom_1(37573) <= 4426801;
srom_1(37574) <= 3930047;
srom_1(37575) <= 3454201;
srom_1(37576) <= 3001495;
srom_1(37577) <= 2574050;
srom_1(37578) <= 2173872;
srom_1(37579) <= 1802837;
srom_1(37580) <= 1462685;
srom_1(37581) <= 1155011;
srom_1(37582) <= 881257;
srom_1(37583) <= 642709;
srom_1(37584) <= 440483;
srom_1(37585) <= 275529;
srom_1(37586) <= 148620;
srom_1(37587) <= 60351;
srom_1(37588) <= 11136;
srom_1(37589) <= 1206;
srom_1(37590) <= 30607;
srom_1(37591) <= 99202;
srom_1(37592) <= 206669;
srom_1(37593) <= 352503;
srom_1(37594) <= 536022;
srom_1(37595) <= 756364;
srom_1(37596) <= 1012496;
srom_1(37597) <= 1303218;
srom_1(37598) <= 1627165;
srom_1(37599) <= 1982819;
srom_1(37600) <= 2368512;
srom_1(37601) <= 2782435;
srom_1(37602) <= 3222648;
srom_1(37603) <= 3687085;
srom_1(37604) <= 4173570;
srom_1(37605) <= 4679820;
srom_1(37606) <= 5203462;
srom_1(37607) <= 5742040;
srom_1(37608) <= 6293029;
srom_1(37609) <= 6853845;
srom_1(37610) <= 7421858;
srom_1(37611) <= 7994404;
srom_1(37612) <= 8568799;
srom_1(37613) <= 9142349;
srom_1(37614) <= 9712364;
srom_1(37615) <= 10276172;
srom_1(37616) <= 10831128;
srom_1(37617) <= 11374630;
srom_1(37618) <= 11904130;
srom_1(37619) <= 12417145;
srom_1(37620) <= 12911268;
srom_1(37621) <= 13384183;
srom_1(37622) <= 13833672;
srom_1(37623) <= 14257627;
srom_1(37624) <= 14654060;
srom_1(37625) <= 15021113;
srom_1(37626) <= 15357063;
srom_1(37627) <= 15660336;
srom_1(37628) <= 15929509;
srom_1(37629) <= 16163321;
srom_1(37630) <= 16360674;
srom_1(37631) <= 16520643;
srom_1(37632) <= 16642478;
srom_1(37633) <= 16725608;
srom_1(37634) <= 16769644;
srom_1(37635) <= 16774377;
srom_1(37636) <= 16739787;
srom_1(37637) <= 16666035;
srom_1(37638) <= 16553467;
srom_1(37639) <= 16402612;
srom_1(37640) <= 16214176;
srom_1(37641) <= 15989044;
srom_1(37642) <= 15728270;
srom_1(37643) <= 15433078;
srom_1(37644) <= 15104853;
srom_1(37645) <= 14745132;
srom_1(37646) <= 14355603;
srom_1(37647) <= 13938094;
srom_1(37648) <= 13494560;
srom_1(37649) <= 13027084;
srom_1(37650) <= 12537855;
srom_1(37651) <= 12029170;
srom_1(37652) <= 11503413;
srom_1(37653) <= 10963049;
srom_1(37654) <= 10410613;
srom_1(37655) <= 9848695;
srom_1(37656) <= 9279930;
srom_1(37657) <= 8706985;
srom_1(37658) <= 8132547;
srom_1(37659) <= 7559311;
srom_1(37660) <= 6989962;
srom_1(37661) <= 6427173;
srom_1(37662) <= 5873582;
srom_1(37663) <= 5331784;
srom_1(37664) <= 4804321;
srom_1(37665) <= 4293666;
srom_1(37666) <= 3802213;
srom_1(37667) <= 3332268;
srom_1(37668) <= 2886033;
srom_1(37669) <= 2465602;
srom_1(37670) <= 2072946;
srom_1(37671) <= 1709906;
srom_1(37672) <= 1378185;
srom_1(37673) <= 1079338;
srom_1(37674) <= 814767;
srom_1(37675) <= 585712;
srom_1(37676) <= 393248;
srom_1(37677) <= 238277;
srom_1(37678) <= 121525;
srom_1(37679) <= 43541;
srom_1(37680) <= 4689;
srom_1(37681) <= 5153;
srom_1(37682) <= 44929;
srom_1(37683) <= 123832;
srom_1(37684) <= 241491;
srom_1(37685) <= 397355;
srom_1(37686) <= 590692;
srom_1(37687) <= 820597;
srom_1(37688) <= 1085990;
srom_1(37689) <= 1385628;
srom_1(37690) <= 1718106;
srom_1(37691) <= 2081863;
srom_1(37692) <= 2475195;
srom_1(37693) <= 2896258;
srom_1(37694) <= 3343075;
srom_1(37695) <= 3813553;
srom_1(37696) <= 4305485;
srom_1(37697) <= 4816564;
srom_1(37698) <= 5344394;
srom_1(37699) <= 5886499;
srom_1(37700) <= 6440337;
srom_1(37701) <= 7003311;
srom_1(37702) <= 7572782;
srom_1(37703) <= 8146078;
srom_1(37704) <= 8720511;
srom_1(37705) <= 9293388;
srom_1(37706) <= 9862023;
srom_1(37707) <= 10423747;
srom_1(37708) <= 10975929;
srom_1(37709) <= 11515977;
srom_1(37710) <= 12041361;
srom_1(37711) <= 12549615;
srom_1(37712) <= 13038356;
srom_1(37713) <= 13505294;
srom_1(37714) <= 13948238;
srom_1(37715) <= 14365110;
srom_1(37716) <= 14753957;
srom_1(37717) <= 15112954;
srom_1(37718) <= 15440419;
srom_1(37719) <= 15734815;
srom_1(37720) <= 15994762;
srom_1(37721) <= 16219042;
srom_1(37722) <= 16406602;
srom_1(37723) <= 16556562;
srom_1(37724) <= 16668221;
srom_1(37725) <= 16741053;
srom_1(37726) <= 16774718;
srom_1(37727) <= 16769058;
srom_1(37728) <= 16724098;
srom_1(37729) <= 16640051;
srom_1(37730) <= 16517310;
srom_1(37731) <= 16356451;
srom_1(37732) <= 16158227;
srom_1(37733) <= 15923570;
srom_1(37734) <= 15653578;
srom_1(37735) <= 15349518;
srom_1(37736) <= 15012816;
srom_1(37737) <= 14645051;
srom_1(37738) <= 14247948;
srom_1(37739) <= 13823367;
srom_1(37740) <= 13373302;
srom_1(37741) <= 12899861;
srom_1(37742) <= 12405266;
srom_1(37743) <= 11891835;
srom_1(37744) <= 11361976;
srom_1(37745) <= 10818175;
srom_1(37746) <= 10262980;
srom_1(37747) <= 9698995;
srom_1(37748) <= 9128866;
srom_1(37749) <= 8555265;
srom_1(37750) <= 7980883;
srom_1(37751) <= 7408413;
srom_1(37752) <= 6840539;
srom_1(37753) <= 6279924;
srom_1(37754) <= 5729198;
srom_1(37755) <= 5190943;
srom_1(37756) <= 4667683;
srom_1(37757) <= 4161871;
srom_1(37758) <= 3675881;
srom_1(37759) <= 3211989;
srom_1(37760) <= 2772373;
srom_1(37761) <= 2359093;
srom_1(37762) <= 1974087;
srom_1(37763) <= 1619162;
srom_1(37764) <= 1295980;
srom_1(37765) <= 1006059;
srom_1(37766) <= 750757;
srom_1(37767) <= 531271;
srom_1(37768) <= 348631;
srom_1(37769) <= 203693;
srom_1(37770) <= 97137;
srom_1(37771) <= 29463;
srom_1(37772) <= 987;
srom_1(37773) <= 11844;
srom_1(37774) <= 61982;
srom_1(37775) <= 151167;
srom_1(37776) <= 278980;
srom_1(37777) <= 444822;
srom_1(37778) <= 647915;
srom_1(37779) <= 887307;
srom_1(37780) <= 1161875;
srom_1(37781) <= 1470331;
srom_1(37782) <= 1811230;
srom_1(37783) <= 2182972;
srom_1(37784) <= 2583815;
srom_1(37785) <= 3011878;
srom_1(37786) <= 3465155;
srom_1(37787) <= 3941519;
srom_1(37788) <= 4438738;
srom_1(37789) <= 4954478;
srom_1(37790) <= 5486323;
srom_1(37791) <= 6031777;
srom_1(37792) <= 6588283;
srom_1(37793) <= 7153231;
srom_1(37794) <= 7723973;
srom_1(37795) <= 8297831;
srom_1(37796) <= 8872115;
srom_1(37797) <= 9444132;
srom_1(37798) <= 10011199;
srom_1(37799) <= 10570657;
srom_1(37800) <= 11119883;
srom_1(37801) <= 11656300;
srom_1(37802) <= 12177395;
srom_1(37803) <= 12680722;
srom_1(37804) <= 13163923;
srom_1(37805) <= 13624730;
srom_1(37806) <= 14060983;
srom_1(37807) <= 14470637;
srom_1(37808) <= 14851769;
srom_1(37809) <= 15202594;
srom_1(37810) <= 15521466;
srom_1(37811) <= 15806889;
srom_1(37812) <= 16057525;
srom_1(37813) <= 16272199;
srom_1(37814) <= 16449905;
srom_1(37815) <= 16589808;
srom_1(37816) <= 16691253;
srom_1(37817) <= 16753763;
srom_1(37818) <= 16777047;
srom_1(37819) <= 16760995;
srom_1(37820) <= 16705681;
srom_1(37821) <= 16611366;
srom_1(37822) <= 16478491;
srom_1(37823) <= 16307681;
srom_1(37824) <= 16099735;
srom_1(37825) <= 15855629;
srom_1(37826) <= 15576507;
srom_1(37827) <= 15263679;
srom_1(37828) <= 14918611;
srom_1(37829) <= 14542922;
srom_1(37830) <= 14138373;
srom_1(37831) <= 13706862;
srom_1(37832) <= 13250411;
srom_1(37833) <= 12771162;
srom_1(37834) <= 12271362;
srom_1(37835) <= 11753353;
srom_1(37836) <= 11219567;
srom_1(37837) <= 10672505;
srom_1(37838) <= 10114733;
srom_1(37839) <= 9548867;
srom_1(37840) <= 8977560;
srom_1(37841) <= 8403491;
srom_1(37842) <= 7829352;
srom_1(37843) <= 7257836;
srom_1(37844) <= 6691622;
srom_1(37845) <= 6133366;
srom_1(37846) <= 5585686;
srom_1(37847) <= 5051149;
srom_1(37848) <= 4532263;
srom_1(37849) <= 4031461;
srom_1(37850) <= 3551091;
srom_1(37851) <= 3093406;
srom_1(37852) <= 2660551;
srom_1(37853) <= 2254558;
srom_1(37854) <= 1877329;
srom_1(37855) <= 1530634;
srom_1(37856) <= 1216098;
srom_1(37857) <= 935196;
srom_1(37858) <= 689247;
srom_1(37859) <= 479402;
srom_1(37860) <= 306646;
srom_1(37861) <= 171789;
srom_1(37862) <= 75464;
srom_1(37863) <= 18121;
srom_1(37864) <= 31;
srom_1(37865) <= 21278;
srom_1(37866) <= 81762;
srom_1(37867) <= 181200;
srom_1(37868) <= 319125;
srom_1(37869) <= 494891;
srom_1(37870) <= 707673;
srom_1(37871) <= 956473;
srom_1(37872) <= 1240125;
srom_1(37873) <= 1557299;
srom_1(37874) <= 1906508;
srom_1(37875) <= 2286113;
srom_1(37876) <= 2694335;
srom_1(37877) <= 3129259;
srom_1(37878) <= 3588846;
srom_1(37879) <= 4070941;
srom_1(37880) <= 4573283;
srom_1(37881) <= 5093516;
srom_1(37882) <= 5629201;
srom_1(37883) <= 6177826;
srom_1(37884) <= 6736818;
srom_1(37885) <= 7303556;
srom_1(37886) <= 7875382;
srom_1(37887) <= 8449615;
srom_1(37888) <= 9023561;
srom_1(37889) <= 9594530;
srom_1(37890) <= 10159844;
srom_1(37891) <= 10716852;
srom_1(37892) <= 11262942;
srom_1(37893) <= 11795554;
srom_1(37894) <= 12312189;
srom_1(37895) <= 12810425;
srom_1(37896) <= 13287925;
srom_1(37897) <= 13742451;
srom_1(37898) <= 14171871;
srom_1(37899) <= 14574172;
srom_1(37900) <= 14947466;
srom_1(37901) <= 15290003;
srom_1(37902) <= 15600177;
srom_1(37903) <= 15876534;
srom_1(37904) <= 16117777;
srom_1(37905) <= 16322776;
srom_1(37906) <= 16490568;
srom_1(37907) <= 16620368;
srom_1(37908) <= 16711566;
srom_1(37909) <= 16763735;
srom_1(37910) <= 16776630;
srom_1(37911) <= 16750191;
srom_1(37912) <= 16684541;
srom_1(37913) <= 16579989;
srom_1(37914) <= 16437024;
srom_1(37915) <= 16256318;
srom_1(37916) <= 16038718;
srom_1(37917) <= 15785243;
srom_1(37918) <= 15497083;
srom_1(37919) <= 15175589;
srom_1(37920) <= 14822268;
srom_1(37921) <= 14438778;
srom_1(37922) <= 14026917;
srom_1(37923) <= 13588615;
srom_1(37924) <= 13125929;
srom_1(37925) <= 12641028;
srom_1(37926) <= 12136186;
srom_1(37927) <= 11613770;
srom_1(37928) <= 11076231;
srom_1(37929) <= 10526088;
srom_1(37930) <= 9965921;
srom_1(37931) <= 9398358;
srom_1(37932) <= 8826061;
srom_1(37933) <= 8251711;
srom_1(37934) <= 7678004;
srom_1(37935) <= 7107629;
srom_1(37936) <= 6543261;
srom_1(37937) <= 5987546;
srom_1(37938) <= 5443091;
srom_1(37939) <= 4912448;
srom_1(37940) <= 4398106;
srom_1(37941) <= 3902477;
srom_1(37942) <= 3427885;
srom_1(37943) <= 2976556;
srom_1(37944) <= 2550605;
srom_1(37945) <= 2152031;
srom_1(37946) <= 1782702;
srom_1(37947) <= 1444351;
srom_1(37948) <= 1138564;
srom_1(37949) <= 866774;
srom_1(37950) <= 630257;
srom_1(37951) <= 430122;
srom_1(37952) <= 267307;
srom_1(37953) <= 142575;
srom_1(37954) <= 56512;
srom_1(37955) <= 9520;
srom_1(37956) <= 1822;
srom_1(37957) <= 33451;
srom_1(37958) <= 104261;
srom_1(37959) <= 213919;
srom_1(37960) <= 361911;
srom_1(37961) <= 547543;
srom_1(37962) <= 769945;
srom_1(37963) <= 1028072;
srom_1(37964) <= 1320716;
srom_1(37965) <= 1646504;
srom_1(37966) <= 2003908;
srom_1(37967) <= 2391252;
srom_1(37968) <= 2806719;
srom_1(37969) <= 3248362;
srom_1(37970) <= 3714109;
srom_1(37971) <= 4201777;
srom_1(37972) <= 4709078;
srom_1(37973) <= 5233633;
srom_1(37974) <= 5772984;
srom_1(37975) <= 6324599;
srom_1(37976) <= 6885894;
srom_1(37977) <= 7454236;
srom_1(37978) <= 8026959;
srom_1(37979) <= 8601378;
srom_1(37980) <= 9174799;
srom_1(37981) <= 9744533;
srom_1(37982) <= 10307909;
srom_1(37983) <= 10862285;
srom_1(37984) <= 11405061;
srom_1(37985) <= 11933692;
srom_1(37986) <= 12445698;
srom_1(37987) <= 12938680;
srom_1(37988) <= 13410324;
srom_1(37989) <= 13858420;
srom_1(37990) <= 14280866;
srom_1(37991) <= 14675682;
srom_1(37992) <= 15041015;
srom_1(37993) <= 15375153;
srom_1(37994) <= 15676528;
srom_1(37995) <= 15943728;
srom_1(37996) <= 16175499;
srom_1(37997) <= 16370755;
srom_1(37998) <= 16528580;
srom_1(37999) <= 16648233;
srom_1(38000) <= 16729155;
srom_1(38001) <= 16770964;
srom_1(38002) <= 16773466;
srom_1(38003) <= 16736649;
srom_1(38004) <= 16660685;
srom_1(38005) <= 16545930;
srom_1(38006) <= 16392922;
srom_1(38007) <= 16202380;
srom_1(38008) <= 15975196;
srom_1(38009) <= 15712436;
srom_1(38010) <= 15415332;
srom_1(38011) <= 15085277;
srom_1(38012) <= 14723819;
srom_1(38013) <= 14332654;
srom_1(38014) <= 13913614;
srom_1(38015) <= 13468666;
srom_1(38016) <= 12999896;
srom_1(38017) <= 12509502;
srom_1(38018) <= 11999783;
srom_1(38019) <= 11473131;
srom_1(38020) <= 10932014;
srom_1(38021) <= 10378970;
srom_1(38022) <= 9816593;
srom_1(38023) <= 9247520;
srom_1(38024) <= 8674418;
srom_1(38025) <= 8099977;
srom_1(38026) <= 7526889;
srom_1(38027) <= 6957841;
srom_1(38028) <= 6395504;
srom_1(38029) <= 5842512;
srom_1(38030) <= 5301460;
srom_1(38031) <= 4774885;
srom_1(38032) <= 4265255;
srom_1(38033) <= 3774962;
srom_1(38034) <= 3306303;
srom_1(38035) <= 2861477;
srom_1(38036) <= 2442570;
srom_1(38037) <= 2051546;
srom_1(38038) <= 1690238;
srom_1(38039) <= 1360342;
srom_1(38040) <= 1063403;
srom_1(38041) <= 800815;
srom_1(38042) <= 573808;
srom_1(38043) <= 383448;
srom_1(38044) <= 230626;
srom_1(38045) <= 116061;
srom_1(38046) <= 40288;
srom_1(38047) <= 3663;
srom_1(38048) <= 6358;
srom_1(38049) <= 48360;
srom_1(38050) <= 129473;
srom_1(38051) <= 249315;
srom_1(38052) <= 407326;
srom_1(38053) <= 602763;
srom_1(38054) <= 834711;
srom_1(38055) <= 1102082;
srom_1(38056) <= 1403621;
srom_1(38057) <= 1737916;
srom_1(38058) <= 2103398;
srom_1(38059) <= 2498354;
srom_1(38060) <= 2920931;
srom_1(38061) <= 3369148;
srom_1(38062) <= 3840902;
srom_1(38063) <= 4333983;
srom_1(38064) <= 4846077;
srom_1(38065) <= 5374783;
srom_1(38066) <= 5917622;
srom_1(38067) <= 6472048;
srom_1(38068) <= 7035462;
srom_1(38069) <= 7605221;
srom_1(38070) <= 8178654;
srom_1(38071) <= 8753071;
srom_1(38072) <= 9325779;
srom_1(38073) <= 9894093;
srom_1(38074) <= 10455346;
srom_1(38075) <= 11006908;
srom_1(38076) <= 11546192;
srom_1(38077) <= 12070669;
srom_1(38078) <= 12577879;
srom_1(38079) <= 13065445;
srom_1(38080) <= 13531079;
srom_1(38081) <= 13972598;
srom_1(38082) <= 14387932;
srom_1(38083) <= 14775134;
srom_1(38084) <= 15132386;
srom_1(38085) <= 15458015;
srom_1(38086) <= 15750493;
srom_1(38087) <= 16008448;
srom_1(38088) <= 16230671;
srom_1(38089) <= 16416120;
srom_1(38090) <= 16563926;
srom_1(38091) <= 16673394;
srom_1(38092) <= 16744013;
srom_1(38093) <= 16775450;
srom_1(38094) <= 16767558;
srom_1(38095) <= 16720374;
srom_1(38096) <= 16634120;
srom_1(38097) <= 16509200;
srom_1(38098) <= 16346199;
srom_1(38099) <= 16145883;
srom_1(38100) <= 15909190;
srom_1(38101) <= 15637231;
srom_1(38102) <= 15331280;
srom_1(38103) <= 14992773;
srom_1(38104) <= 14623296;
srom_1(38105) <= 14224583;
srom_1(38106) <= 13798503;
srom_1(38107) <= 13347054;
srom_1(38108) <= 12872353;
srom_1(38109) <= 12376627;
srom_1(38110) <= 11862199;
srom_1(38111) <= 11331482;
srom_1(38112) <= 10786965;
srom_1(38113) <= 10231202;
srom_1(38114) <= 9666798;
srom_1(38115) <= 9096400;
srom_1(38116) <= 8522683;
srom_1(38117) <= 7948337;
srom_1(38118) <= 7376055;
srom_1(38119) <= 6808522;
srom_1(38120) <= 6248399;
srom_1(38121) <= 5698312;
srom_1(38122) <= 5160840;
srom_1(38123) <= 4638505;
srom_1(38124) <= 4133755;
srom_1(38125) <= 3648957;
srom_1(38126) <= 3186386;
srom_1(38127) <= 2748209;
srom_1(38128) <= 2336482;
srom_1(38129) <= 1953136;
srom_1(38130) <= 1599967;
srom_1(38131) <= 1278633;
srom_1(38132) <= 990640;
srom_1(38133) <= 737339;
srom_1(38134) <= 519917;
srom_1(38135) <= 339394;
srom_1(38136) <= 196617;
srom_1(38137) <= 92255;
srom_1(38138) <= 26797;
srom_1(38139) <= 550;
srom_1(38140) <= 13638;
srom_1(38141) <= 65999;
srom_1(38142) <= 157388;
srom_1(38143) <= 287376;
srom_1(38144) <= 455353;
srom_1(38145) <= 660532;
srom_1(38146) <= 901950;
srom_1(38147) <= 1178476;
srom_1(38148) <= 1488813;
srom_1(38149) <= 1831505;
srom_1(38150) <= 2204946;
srom_1(38151) <= 2607384;
srom_1(38152) <= 3036932;
srom_1(38153) <= 3491577;
srom_1(38154) <= 3969184;
srom_1(38155) <= 4467517;
srom_1(38156) <= 4984236;
srom_1(38157) <= 5516920;
srom_1(38158) <= 6063070;
srom_1(38159) <= 6620125;
srom_1(38160) <= 7185473;
srom_1(38161) <= 7756463;
srom_1(38162) <= 8330418;
srom_1(38163) <= 8904645;
srom_1(38164) <= 9476453;
srom_1(38165) <= 10043159;
srom_1(38166) <= 10602107;
srom_1(38167) <= 11150674;
srom_1(38168) <= 11686289;
srom_1(38169) <= 12206441;
srom_1(38170) <= 12708689;
srom_1(38171) <= 13190679;
srom_1(38172) <= 13650150;
srom_1(38173) <= 14084948;
srom_1(38174) <= 14493034;
srom_1(38175) <= 14872494;
srom_1(38176) <= 15221550;
srom_1(38177) <= 15538563;
srom_1(38178) <= 15822047;
srom_1(38179) <= 16070674;
srom_1(38180) <= 16283276;
srom_1(38181) <= 16458858;
srom_1(38182) <= 16596596;
srom_1(38183) <= 16695843;
srom_1(38184) <= 16756135;
srom_1(38185) <= 16777189;
srom_1(38186) <= 16758906;
srom_1(38187) <= 16701372;
srom_1(38188) <= 16604856;
srom_1(38189) <= 16469811;
srom_1(38190) <= 16296871;
srom_1(38191) <= 16086847;
srom_1(38192) <= 15840722;
srom_1(38193) <= 15559652;
srom_1(38194) <= 15244955;
srom_1(38195) <= 14898106;
srom_1(38196) <= 14520732;
srom_1(38197) <= 14114601;
srom_1(38198) <= 13681620;
srom_1(38199) <= 13223818;
srom_1(38200) <= 12743342;
srom_1(38201) <= 12242445;
srom_1(38202) <= 11723477;
srom_1(38203) <= 11188870;
srom_1(38204) <= 10641131;
srom_1(38205) <= 10082830;
srom_1(38206) <= 9516583;
srom_1(38207) <= 8945048;
srom_1(38208) <= 8370903;
srom_1(38209) <= 7796841;
srom_1(38210) <= 7225554;
srom_1(38211) <= 6659721;
srom_1(38212) <= 6101995;
srom_1(38213) <= 5554992;
srom_1(38214) <= 5021277;
srom_1(38215) <= 4503352;
srom_1(38216) <= 4003647;
srom_1(38217) <= 3524504;
srom_1(38218) <= 3068171;
srom_1(38219) <= 2636787;
srom_1(38220) <= 2232375;
srom_1(38221) <= 1856832;
srom_1(38222) <= 1511919;
srom_1(38223) <= 1199253;
srom_1(38224) <= 920300;
srom_1(38225) <= 676369;
srom_1(38226) <= 468603;
srom_1(38227) <= 297976;
srom_1(38228) <= 165290;
srom_1(38229) <= 71165;
srom_1(38230) <= 16044;
srom_1(38231) <= 184;
srom_1(38232) <= 23661;
srom_1(38233) <= 86364;
srom_1(38234) <= 187998;
srom_1(38235) <= 328089;
srom_1(38236) <= 505978;
srom_1(38237) <= 720831;
srom_1(38238) <= 971641;
srom_1(38239) <= 1257232;
srom_1(38240) <= 1576264;
srom_1(38241) <= 1927241;
srom_1(38242) <= 2308519;
srom_1(38243) <= 2718307;
srom_1(38244) <= 3154686;
srom_1(38245) <= 3615609;
srom_1(38246) <= 4098913;
srom_1(38247) <= 4602334;
srom_1(38248) <= 5123510;
srom_1(38249) <= 5659996;
srom_1(38250) <= 6209279;
srom_1(38251) <= 6768780;
srom_1(38252) <= 7335878;
srom_1(38253) <= 7907912;
srom_1(38254) <= 8482201;
srom_1(38255) <= 9056051;
srom_1(38256) <= 9626770;
srom_1(38257) <= 10191684;
srom_1(38258) <= 10748142;
srom_1(38259) <= 11293536;
srom_1(38260) <= 11825307;
srom_1(38261) <= 12340963;
srom_1(38262) <= 12838084;
srom_1(38263) <= 13314341;
srom_1(38264) <= 13767499;
srom_1(38265) <= 14195433;
srom_1(38266) <= 14596137;
srom_1(38267) <= 14967733;
srom_1(38268) <= 15308476;
srom_1(38269) <= 15616769;
srom_1(38270) <= 15891168;
srom_1(38271) <= 16130384;
srom_1(38272) <= 16333296;
srom_1(38273) <= 16498953;
srom_1(38274) <= 16626578;
srom_1(38275) <= 16715572;
srom_1(38276) <= 16765518;
srom_1(38277) <= 16776182;
srom_1(38278) <= 16747514;
srom_1(38279) <= 16679648;
srom_1(38280) <= 16572902;
srom_1(38281) <= 16427777;
srom_1(38282) <= 16244954;
srom_1(38283) <= 16025290;
srom_1(38284) <= 15769815;
srom_1(38285) <= 15479727;
srom_1(38286) <= 15156386;
srom_1(38287) <= 14801308;
srom_1(38288) <= 14416159;
srom_1(38289) <= 14002745;
srom_1(38290) <= 13563005;
srom_1(38291) <= 13099000;
srom_1(38292) <= 12612906;
srom_1(38293) <= 12107003;
srom_1(38294) <= 11583663;
srom_1(38295) <= 11045340;
srom_1(38296) <= 10494559;
srom_1(38297) <= 9933903;
srom_1(38298) <= 9366000;
srom_1(38299) <= 8793514;
srom_1(38300) <= 8219129;
srom_1(38301) <= 7645539;
srom_1(38302) <= 7075433;
srom_1(38303) <= 6511485;
srom_1(38304) <= 5956340;
srom_1(38305) <= 5412600;
srom_1(38306) <= 4882816;
srom_1(38307) <= 4369472;
srom_1(38308) <= 3874975;
srom_1(38309) <= 3401644;
srom_1(38310) <= 2951698;
srom_1(38311) <= 2527248;
srom_1(38312) <= 2130284;
srom_1(38313) <= 1762667;
srom_1(38314) <= 1426122;
srom_1(38315) <= 1122226;
srom_1(38316) <= 852405;
srom_1(38317) <= 617923;
srom_1(38318) <= 419881;
srom_1(38319) <= 259207;
srom_1(38320) <= 136654;
srom_1(38321) <= 52798;
srom_1(38322) <= 8031;
srom_1(38323) <= 2564;
srom_1(38324) <= 36422;
srom_1(38325) <= 109446;
srom_1(38326) <= 221293;
srom_1(38327) <= 371441;
srom_1(38328) <= 559183;
srom_1(38329) <= 783640;
srom_1(38330) <= 1043760;
srom_1(38331) <= 1338322;
srom_1(38332) <= 1665945;
srom_1(38333) <= 2025093;
srom_1(38334) <= 2414082;
srom_1(38335) <= 2831087;
srom_1(38336) <= 3274154;
srom_1(38337) <= 3741204;
srom_1(38338) <= 4230047;
srom_1(38339) <= 4738391;
srom_1(38340) <= 5263852;
srom_1(38341) <= 5803966;
srom_1(38342) <= 6356201;
srom_1(38343) <= 6917966;
srom_1(38344) <= 7486628;
srom_1(38345) <= 8059519;
srom_1(38346) <= 8633953;
srom_1(38347) <= 9207237;
srom_1(38348) <= 9776682;
srom_1(38349) <= 10339618;
srom_1(38350) <= 10893405;
srom_1(38351) <= 11435446;
srom_1(38352) <= 11963200;
srom_1(38353) <= 12474191;
srom_1(38354) <= 12966023;
srom_1(38355) <= 13436390;
srom_1(38356) <= 13883086;
srom_1(38357) <= 14304017;
srom_1(38358) <= 14697208;
srom_1(38359) <= 15060817;
srom_1(38360) <= 15393137;
srom_1(38361) <= 15692610;
srom_1(38362) <= 15957832;
srom_1(38363) <= 16187560;
srom_1(38364) <= 16380716;
srom_1(38365) <= 16536393;
srom_1(38366) <= 16653864;
srom_1(38367) <= 16732575;
srom_1(38368) <= 16772159;
srom_1(38369) <= 16772429;
srom_1(38370) <= 16733385;
srom_1(38371) <= 16655209;
srom_1(38372) <= 16538269;
srom_1(38373) <= 16383111;
srom_1(38374) <= 16190465;
srom_1(38375) <= 15961233;
srom_1(38376) <= 15696491;
srom_1(38377) <= 15397479;
srom_1(38378) <= 15065600;
srom_1(38379) <= 14702411;
srom_1(38380) <= 14309614;
srom_1(38381) <= 13889051;
srom_1(38382) <= 13442695;
srom_1(38383) <= 12972639;
srom_1(38384) <= 12481086;
srom_1(38385) <= 11970343;
srom_1(38386) <= 11442803;
srom_1(38387) <= 10900941;
srom_1(38388) <= 10347298;
srom_1(38389) <= 9784470;
srom_1(38390) <= 9215097;
srom_1(38391) <= 8641847;
srom_1(38392) <= 8067410;
srom_1(38393) <= 7494480;
srom_1(38394) <= 6925742;
srom_1(38395) <= 6363864;
srom_1(38396) <= 5811481;
srom_1(38397) <= 5271183;
srom_1(38398) <= 4745503;
srom_1(38399) <= 4236907;
srom_1(38400) <= 3747780;
srom_1(38401) <= 3280416;
srom_1(38402) <= 2837005;
srom_1(38403) <= 2419628;
srom_1(38404) <= 2030242;
srom_1(38405) <= 1670672;
srom_1(38406) <= 1342604;
srom_1(38407) <= 1047578;
srom_1(38408) <= 786976;
srom_1(38409) <= 562022;
srom_1(38410) <= 373768;
srom_1(38411) <= 223099;
srom_1(38412) <= 110721;
srom_1(38413) <= 37161;
srom_1(38414) <= 2763;
srom_1(38415) <= 7690;
srom_1(38416) <= 51917;
srom_1(38417) <= 135238;
srom_1(38418) <= 257262;
srom_1(38419) <= 417417;
srom_1(38420) <= 614952;
srom_1(38421) <= 848939;
srom_1(38422) <= 1118283;
srom_1(38423) <= 1421720;
srom_1(38424) <= 1757827;
srom_1(38425) <= 2125028;
srom_1(38426) <= 2521601;
srom_1(38427) <= 2945686;
srom_1(38428) <= 3395295;
srom_1(38429) <= 3868320;
srom_1(38430) <= 4362542;
srom_1(38431) <= 4875643;
srom_1(38432) <= 5405218;
srom_1(38433) <= 5948783;
srom_1(38434) <= 6503789;
srom_1(38435) <= 7067633;
srom_1(38436) <= 7637673;
srom_1(38437) <= 8211233;
srom_1(38438) <= 8785625;
srom_1(38439) <= 9358156;
srom_1(38440) <= 9926140;
srom_1(38441) <= 10486914;
srom_1(38442) <= 11037848;
srom_1(38443) <= 11576359;
srom_1(38444) <= 12099922;
srom_1(38445) <= 12606081;
srom_1(38446) <= 13092463;
srom_1(38447) <= 13556786;
srom_1(38448) <= 13996875;
srom_1(38449) <= 14410664;
srom_1(38450) <= 14796214;
srom_1(38451) <= 15151716;
srom_1(38452) <= 15475504;
srom_1(38453) <= 15766059;
srom_1(38454) <= 16022019;
srom_1(38455) <= 16242182;
srom_1(38456) <= 16425518;
srom_1(38457) <= 16571166;
srom_1(38458) <= 16678443;
srom_1(38459) <= 16746846;
srom_1(38460) <= 16776055;
srom_1(38461) <= 16765931;
srom_1(38462) <= 16716524;
srom_1(38463) <= 16628064;
srom_1(38464) <= 16500967;
srom_1(38465) <= 16335828;
srom_1(38466) <= 16133422;
srom_1(38467) <= 15894697;
srom_1(38468) <= 15620774;
srom_1(38469) <= 15312937;
srom_1(38470) <= 14972629;
srom_1(38471) <= 14601447;
srom_1(38472) <= 14201130;
srom_1(38473) <= 13773557;
srom_1(38474) <= 13320731;
srom_1(38475) <= 12844777;
srom_1(38476) <= 12347927;
srom_1(38477) <= 11832510;
srom_1(38478) <= 11300943;
srom_1(38479) <= 10755720;
srom_1(38480) <= 10199396;
srom_1(38481) <= 9634581;
srom_1(38482) <= 9063923;
srom_1(38483) <= 8490098;
srom_1(38484) <= 7915797;
srom_1(38485) <= 7343714;
srom_1(38486) <= 6776530;
srom_1(38487) <= 6216906;
srom_1(38488) <= 5667466;
srom_1(38489) <= 5130786;
srom_1(38490) <= 4609383;
srom_1(38491) <= 4105702;
srom_1(38492) <= 3622105;
srom_1(38493) <= 3160860;
srom_1(38494) <= 2724130;
srom_1(38495) <= 2313962;
srom_1(38496) <= 1932281;
srom_1(38497) <= 1580875;
srom_1(38498) <= 1261393;
srom_1(38499) <= 975334;
srom_1(38500) <= 724037;
srom_1(38501) <= 508682;
srom_1(38502) <= 330279;
srom_1(38503) <= 189665;
srom_1(38504) <= 87498;
srom_1(38505) <= 24257;
srom_1(38506) <= 240;
srom_1(38507) <= 15559;
srom_1(38508) <= 70142;
srom_1(38509) <= 163733;
srom_1(38510) <= 295894;
srom_1(38511) <= 466004;
srom_1(38512) <= 673265;
srom_1(38513) <= 916707;
srom_1(38514) <= 1195187;
srom_1(38515) <= 1507399;
srom_1(38516) <= 1851880;
srom_1(38517) <= 2227013;
srom_1(38518) <= 2631041;
srom_1(38519) <= 3062067;
srom_1(38520) <= 3518072;
srom_1(38521) <= 3996916;
srom_1(38522) <= 4496355;
srom_1(38523) <= 5014045;
srom_1(38524) <= 5547560;
srom_1(38525) <= 6094398;
srom_1(38526) <= 6651994;
srom_1(38527) <= 7217733;
srom_1(38528) <= 7788963;
srom_1(38529) <= 8363005;
srom_1(38530) <= 8937167;
srom_1(38531) <= 9508757;
srom_1(38532) <= 10075094;
srom_1(38533) <= 10633523;
srom_1(38534) <= 11181424;
srom_1(38535) <= 11716229;
srom_1(38536) <= 12235429;
srom_1(38537) <= 12736590;
srom_1(38538) <= 13217363;
srom_1(38539) <= 13675491;
srom_1(38540) <= 14108827;
srom_1(38541) <= 14515340;
srom_1(38542) <= 14893122;
srom_1(38543) <= 15240402;
srom_1(38544) <= 15555552;
srom_1(38545) <= 15837093;
srom_1(38546) <= 16083706;
srom_1(38547) <= 16294234;
srom_1(38548) <= 16467690;
srom_1(38549) <= 16603260;
srom_1(38550) <= 16700308;
srom_1(38551) <= 16758381;
srom_1(38552) <= 16777204;
srom_1(38553) <= 16756691;
srom_1(38554) <= 16696937;
srom_1(38555) <= 16598222;
srom_1(38556) <= 16461009;
srom_1(38557) <= 16285943;
srom_1(38558) <= 16073842;
srom_1(38559) <= 15825704;
srom_1(38560) <= 15542690;
srom_1(38561) <= 15226128;
srom_1(38562) <= 14877502;
srom_1(38563) <= 14498448;
srom_1(38564) <= 14090743;
srom_1(38565) <= 13656299;
srom_1(38566) <= 13197152;
srom_1(38567) <= 12715457;
srom_1(38568) <= 12213471;
srom_1(38569) <= 11693550;
srom_1(38570) <= 11158130;
srom_1(38571) <= 10609723;
srom_1(38572) <= 10050901;
srom_1(38573) <= 9484283;
srom_1(38574) <= 8912528;
srom_1(38575) <= 8338315;
srom_1(38576) <= 7764339;
srom_1(38577) <= 7193290;
srom_1(38578) <= 6627846;
srom_1(38579) <= 6070659;
srom_1(38580) <= 5524341;
srom_1(38581) <= 4991455;
srom_1(38582) <= 4474500;
srom_1(38583) <= 3975899;
srom_1(38584) <= 3497991;
srom_1(38585) <= 3043016;
srom_1(38586) <= 2613109;
srom_1(38587) <= 2210285;
srom_1(38588) <= 1836434;
srom_1(38589) <= 1493308;
srom_1(38590) <= 1182516;
srom_1(38591) <= 905516;
srom_1(38592) <= 663607;
srom_1(38593) <= 457923;
srom_1(38594) <= 289429;
srom_1(38595) <= 158914;
srom_1(38596) <= 66992;
srom_1(38597) <= 14092;
srom_1(38598) <= 464;
srom_1(38599) <= 26170;
srom_1(38600) <= 91090;
srom_1(38601) <= 194921;
srom_1(38602) <= 337174;
srom_1(38603) <= 517184;
srom_1(38604) <= 734105;
srom_1(38605) <= 986921;
srom_1(38606) <= 1274445;
srom_1(38607) <= 1595331;
srom_1(38608) <= 1948073;
srom_1(38609) <= 2331016;
srom_1(38610) <= 2742366;
srom_1(38611) <= 3180192;
srom_1(38612) <= 3642443;
srom_1(38613) <= 4126950;
srom_1(38614) <= 4631442;
srom_1(38615) <= 5153552;
srom_1(38616) <= 5690833;
srom_1(38617) <= 6240764;
srom_1(38618) <= 6800767;
srom_1(38619) <= 7368216;
srom_1(38620) <= 7940450;
srom_1(38621) <= 8514786;
srom_1(38622) <= 9088530;
srom_1(38623) <= 9658992;
srom_1(38624) <= 10223496;
srom_1(38625) <= 10779396;
srom_1(38626) <= 11324085;
srom_1(38627) <= 11855009;
srom_1(38628) <= 12369677;
srom_1(38629) <= 12865676;
srom_1(38630) <= 13340682;
srom_1(38631) <= 13792465;
srom_1(38632) <= 14218907;
srom_1(38633) <= 14618010;
srom_1(38634) <= 14987900;
srom_1(38635) <= 15326844;
srom_1(38636) <= 15633253;
srom_1(38637) <= 15905688;
srom_1(38638) <= 16142874;
srom_1(38639) <= 16343697;
srom_1(38640) <= 16507216;
srom_1(38641) <= 16632664;
srom_1(38642) <= 16719453;
srom_1(38643) <= 16767175;
srom_1(38644) <= 16775608;
srom_1(38645) <= 16744711;
srom_1(38646) <= 16674629;
srom_1(38647) <= 16565692;
srom_1(38648) <= 16418409;
srom_1(38649) <= 16233472;
srom_1(38650) <= 16011747;
srom_1(38651) <= 15754275;
srom_1(38652) <= 15462263;
srom_1(38653) <= 15137080;
srom_1(38654) <= 14780251;
srom_1(38655) <= 14393450;
srom_1(38656) <= 13978489;
srom_1(38657) <= 13537316;
srom_1(38658) <= 13071999;
srom_1(38659) <= 12584720;
srom_1(38660) <= 12077763;
srom_1(38661) <= 11553507;
srom_1(38662) <= 11014410;
srom_1(38663) <= 10462999;
srom_1(38664) <= 9901861;
srom_1(38665) <= 9333627;
srom_1(38666) <= 8760961;
srom_1(38667) <= 8186549;
srom_1(38668) <= 7613085;
srom_1(38669) <= 7043257;
srom_1(38670) <= 6479738;
srom_1(38671) <= 5925170;
srom_1(38672) <= 5382155;
srom_1(38673) <= 4853237;
srom_1(38674) <= 4340898;
srom_1(38675) <= 3847541;
srom_1(38676) <= 3375477;
srom_1(38677) <= 2926923;
srom_1(38678) <= 2503979;
srom_1(38679) <= 2108631;
srom_1(38680) <= 1742732;
srom_1(38681) <= 1407998;
srom_1(38682) <= 1105998;
srom_1(38683) <= 838149;
srom_1(38684) <= 605706;
srom_1(38685) <= 409760;
srom_1(38686) <= 251230;
srom_1(38687) <= 130859;
srom_1(38688) <= 49211;
srom_1(38689) <= 6669;
srom_1(38690) <= 3433;
srom_1(38691) <= 39518;
srom_1(38692) <= 114755;
srom_1(38693) <= 228791;
srom_1(38694) <= 381091;
srom_1(38695) <= 570941;
srom_1(38696) <= 797450;
srom_1(38697) <= 1059558;
srom_1(38698) <= 1356033;
srom_1(38699) <= 1685487;
srom_1(38700) <= 2046374;
srom_1(38701) <= 2437002;
srom_1(38702) <= 2855539;
srom_1(38703) <= 3300023;
srom_1(38704) <= 3768368;
srom_1(38705) <= 4258380;
srom_1(38706) <= 4767759;
srom_1(38707) <= 5294118;
srom_1(38708) <= 5834988;
srom_1(38709) <= 6387833;
srom_1(38710) <= 6950060;
srom_1(38711) <= 7519033;
srom_1(38712) <= 8092084;
srom_1(38713) <= 8666525;
srom_1(38714) <= 9239663;
srom_1(38715) <= 9808810;
srom_1(38716) <= 10371298;
srom_1(38717) <= 10924487;
srom_1(38718) <= 11465785;
srom_1(38719) <= 11992654;
srom_1(38720) <= 12502621;
srom_1(38721) <= 12993297;
srom_1(38722) <= 13462379;
srom_1(38723) <= 13907669;
srom_1(38724) <= 14327078;
srom_1(38725) <= 14718640;
srom_1(38726) <= 15080518;
srom_1(38727) <= 15411015;
srom_1(38728) <= 15708582;
srom_1(38729) <= 15971822;
srom_1(38730) <= 16199503;
srom_1(38731) <= 16390556;
srom_1(38732) <= 16544084;
srom_1(38733) <= 16659369;
srom_1(38734) <= 16735869;
srom_1(38735) <= 16773227;
srom_1(38736) <= 16771265;
srom_1(38737) <= 16729995;
srom_1(38738) <= 16649609;
srom_1(38739) <= 16530485;
srom_1(38740) <= 16373180;
srom_1(38741) <= 16178433;
srom_1(38742) <= 15947156;
srom_1(38743) <= 15680435;
srom_1(38744) <= 15379521;
srom_1(38745) <= 15045823;
srom_1(38746) <= 14680907;
srom_1(38747) <= 14286485;
srom_1(38748) <= 13864406;
srom_1(38749) <= 13416648;
srom_1(38750) <= 12945312;
srom_1(38751) <= 12452609;
srom_1(38752) <= 11940848;
srom_1(38753) <= 11412429;
srom_1(38754) <= 10869830;
srom_1(38755) <= 10315597;
srom_1(38756) <= 9752326;
srom_1(38757) <= 9182661;
srom_1(38758) <= 8609273;
srom_1(38759) <= 8034849;
srom_1(38760) <= 7462084;
srom_1(38761) <= 6893665;
srom_1(38762) <= 6332255;
srom_1(38763) <= 5780489;
srom_1(38764) <= 5240952;
srom_1(38765) <= 4716176;
srom_1(38766) <= 4208622;
srom_1(38767) <= 3720669;
srom_1(38768) <= 3254605;
srom_1(38769) <= 2812617;
srom_1(38770) <= 2396776;
srom_1(38771) <= 2009033;
srom_1(38772) <= 1651206;
srom_1(38773) <= 1324973;
srom_1(38774) <= 1031864;
srom_1(38775) <= 773253;
srom_1(38776) <= 550353;
srom_1(38777) <= 364210;
srom_1(38778) <= 215695;
srom_1(38779) <= 105506;
srom_1(38780) <= 34160;
srom_1(38781) <= 1990;
srom_1(38782) <= 9148;
srom_1(38783) <= 55600;
srom_1(38784) <= 141129;
srom_1(38785) <= 265332;
srom_1(38786) <= 427629;
srom_1(38787) <= 627257;
srom_1(38788) <= 863281;
srom_1(38789) <= 1134594;
srom_1(38790) <= 1439924;
srom_1(38791) <= 1777838;
srom_1(38792) <= 2146752;
srom_1(38793) <= 2544937;
srom_1(38794) <= 2970524;
srom_1(38795) <= 3421519;
srom_1(38796) <= 3895806;
srom_1(38797) <= 4391161;
srom_1(38798) <= 4905262;
srom_1(38799) <= 5435697;
srom_1(38800) <= 5979980;
srom_1(38801) <= 6535558;
srom_1(38802) <= 7099825;
srom_1(38803) <= 7670135;
srom_1(38804) <= 8243815;
srom_1(38805) <= 8818174;
srom_1(38806) <= 9390518;
srom_1(38807) <= 9958164;
srom_1(38808) <= 10518450;
srom_1(38809) <= 11068748;
srom_1(38810) <= 11606478;
srom_1(38811) <= 12129119;
srom_1(38812) <= 12634219;
srom_1(38813) <= 13119409;
srom_1(38814) <= 13582416;
srom_1(38815) <= 14021067;
srom_1(38816) <= 14433305;
srom_1(38817) <= 14817198;
srom_1(38818) <= 15170945;
srom_1(38819) <= 15492887;
srom_1(38820) <= 15781514;
srom_1(38821) <= 16035474;
srom_1(38822) <= 16253575;
srom_1(38823) <= 16434794;
srom_1(38824) <= 16578283;
srom_1(38825) <= 16683366;
srom_1(38826) <= 16749553;
srom_1(38827) <= 16776533;
srom_1(38828) <= 16764179;
srom_1(38829) <= 16712548;
srom_1(38830) <= 16621884;
srom_1(38831) <= 16492612;
srom_1(38832) <= 16325336;
srom_1(38833) <= 16120843;
srom_1(38834) <= 15880091;
srom_1(38835) <= 15604208;
srom_1(38836) <= 15294489;
srom_1(38837) <= 14952386;
srom_1(38838) <= 14579504;
srom_1(38839) <= 14177590;
srom_1(38840) <= 13748529;
srom_1(38841) <= 13294334;
srom_1(38842) <= 12817134;
srom_1(38843) <= 12319167;
srom_1(38844) <= 11802769;
srom_1(38845) <= 11270361;
srom_1(38846) <= 10724438;
srom_1(38847) <= 10167563;
srom_1(38848) <= 9602345;
srom_1(38849) <= 9031436;
srom_1(38850) <= 8457512;
srom_1(38851) <= 7883265;
srom_1(38852) <= 7311388;
srom_1(38853) <= 6744562;
srom_1(38854) <= 6185445;
srom_1(38855) <= 5636661;
srom_1(38856) <= 5100780;
srom_1(38857) <= 4580318;
srom_1(38858) <= 4077714;
srom_1(38859) <= 3595325;
srom_1(38860) <= 3135414;
srom_1(38861) <= 2700137;
srom_1(38862) <= 2291534;
srom_1(38863) <= 1911524;
srom_1(38864) <= 1561886;
srom_1(38865) <= 1244261;
srom_1(38866) <= 960139;
srom_1(38867) <= 710851;
srom_1(38868) <= 497566;
srom_1(38869) <= 321286;
srom_1(38870) <= 182836;
srom_1(38871) <= 82866;
srom_1(38872) <= 21844;
srom_1(38873) <= 57;
srom_1(38874) <= 17606;
srom_1(38875) <= 74410;
srom_1(38876) <= 170202;
srom_1(38877) <= 304534;
srom_1(38878) <= 476774;
srom_1(38879) <= 686115;
srom_1(38880) <= 931576;
srom_1(38881) <= 1212006;
srom_1(38882) <= 1526089;
srom_1(38883) <= 1872353;
srom_1(38884) <= 2249173;
srom_1(38885) <= 2654784;
srom_1(38886) <= 3087283;
srom_1(38887) <= 3544641;
srom_1(38888) <= 4024714;
srom_1(38889) <= 4525252;
srom_1(38890) <= 5043905;
srom_1(38891) <= 5578243;
srom_1(38892) <= 6125760;
srom_1(38893) <= 6683889;
srom_1(38894) <= 7250011;
srom_1(38895) <= 7821472;
srom_1(38896) <= 8395593;
srom_1(38897) <= 8969681;
srom_1(38898) <= 9541045;
srom_1(38899) <= 10107004;
srom_1(38900) <= 10664905;
srom_1(38901) <= 11212131;
srom_1(38902) <= 11746118;
srom_1(38903) <= 12264359;
srom_1(38904) <= 12764426;
srom_1(38905) <= 13243973;
srom_1(38906) <= 13700752;
srom_1(38907) <= 14132620;
srom_1(38908) <= 14537553;
srom_1(38909) <= 14913651;
srom_1(38910) <= 15259151;
srom_1(38911) <= 15572432;
srom_1(38912) <= 15852027;
srom_1(38913) <= 16096622;
srom_1(38914) <= 16305072;
srom_1(38915) <= 16476399;
srom_1(38916) <= 16609800;
srom_1(38917) <= 16704648;
srom_1(38918) <= 16760500;
srom_1(38919) <= 16777093;
srom_1(38920) <= 16754350;
srom_1(38921) <= 16692377;
srom_1(38922) <= 16591464;
srom_1(38923) <= 16452086;
srom_1(38924) <= 16274895;
srom_1(38925) <= 16060722;
srom_1(38926) <= 15810573;
srom_1(38927) <= 15525619;
srom_1(38928) <= 15207197;
srom_1(38929) <= 14856801;
srom_1(38930) <= 14476073;
srom_1(38931) <= 14066799;
srom_1(38932) <= 13630898;
srom_1(38933) <= 13170414;
srom_1(38934) <= 12687506;
srom_1(38935) <= 12184439;
srom_1(38936) <= 11663573;
srom_1(38937) <= 11127349;
srom_1(38938) <= 10578282;
srom_1(38939) <= 10018947;
srom_1(38940) <= 9451966;
srom_1(38941) <= 8880000;
srom_1(38942) <= 8305728;
srom_1(38943) <= 7731846;
srom_1(38944) <= 7161043;
srom_1(38945) <= 6595997;
srom_1(38946) <= 6039357;
srom_1(38947) <= 5493734;
srom_1(38948) <= 4961685;
srom_1(38949) <= 4445707;
srom_1(38950) <= 3948218;
srom_1(38951) <= 3471551;
srom_1(38952) <= 3017943;
srom_1(38953) <= 2589519;
srom_1(38954) <= 2188289;
srom_1(38955) <= 1816135;
srom_1(38956) <= 1474801;
srom_1(38957) <= 1165888;
srom_1(38958) <= 890845;
srom_1(38959) <= 650962;
srom_1(38960) <= 447363;
srom_1(38961) <= 281004;
srom_1(38962) <= 152663;
srom_1(38963) <= 62944;
srom_1(38964) <= 12267;
srom_1(38965) <= 870;
srom_1(38966) <= 28805;
srom_1(38967) <= 95942;
srom_1(38968) <= 201967;
srom_1(38969) <= 346381;
srom_1(38970) <= 528508;
srom_1(38971) <= 747494;
srom_1(38972) <= 1002312;
srom_1(38973) <= 1291767;
srom_1(38974) <= 1614501;
srom_1(38975) <= 1969001;
srom_1(38976) <= 2353605;
srom_1(38977) <= 2766509;
srom_1(38978) <= 3205777;
srom_1(38979) <= 3669349;
srom_1(38980) <= 4155052;
srom_1(38981) <= 4660607;
srom_1(38982) <= 5183643;
srom_1(38983) <= 5721709;
srom_1(38984) <= 6272281;
srom_1(38985) <= 6832778;
srom_1(38986) <= 7400570;
srom_1(38987) <= 7972995;
srom_1(38988) <= 8547369;
srom_1(38989) <= 9120999;
srom_1(38990) <= 9691194;
srom_1(38991) <= 10255281;
srom_1(38992) <= 10810615;
srom_1(38993) <= 11354590;
srom_1(38994) <= 11884658;
srom_1(38995) <= 12398331;
srom_1(38996) <= 12893201;
srom_1(38997) <= 13366948;
srom_1(38998) <= 13817349;
srom_1(38999) <= 14242293;
srom_1(39000) <= 14639788;
srom_1(39001) <= 15007968;
srom_1(39002) <= 15345108;
srom_1(39003) <= 15649626;
srom_1(39004) <= 15920095;
srom_1(39005) <= 16155247;
srom_1(39006) <= 16353977;
srom_1(39007) <= 16515356;
srom_1(39008) <= 16638625;
srom_1(39009) <= 16723207;
srom_1(39010) <= 16768706;
srom_1(39011) <= 16774907;
srom_1(39012) <= 16741782;
srom_1(39013) <= 16669486;
srom_1(39014) <= 16558358;
srom_1(39015) <= 16408920;
srom_1(39016) <= 16221871;
srom_1(39017) <= 15998090;
srom_1(39018) <= 15738625;
srom_1(39019) <= 15444693;
srom_1(39020) <= 15117673;
srom_1(39021) <= 14759098;
srom_1(39022) <= 14370649;
srom_1(39023) <= 13954149;
srom_1(39024) <= 13511550;
srom_1(39025) <= 13044928;
srom_1(39026) <= 12556470;
srom_1(39027) <= 12048468;
srom_1(39028) <= 11523304;
srom_1(39029) <= 10983440;
srom_1(39030) <= 10431408;
srom_1(39031) <= 9869797;
srom_1(39032) <= 9301239;
srom_1(39033) <= 8728403;
srom_1(39034) <= 8153972;
srom_1(39035) <= 7580642;
srom_1(39036) <= 7011101;
srom_1(39037) <= 6448020;
srom_1(39038) <= 5894038;
srom_1(39039) <= 5351754;
srom_1(39040) <= 4823712;
srom_1(39041) <= 4312386;
srom_1(39042) <= 3820175;
srom_1(39043) <= 3349387;
srom_1(39044) <= 2902229;
srom_1(39045) <= 2480800;
srom_1(39046) <= 2087073;
srom_1(39047) <= 1722897;
srom_1(39048) <= 1389979;
srom_1(39049) <= 1089880;
srom_1(39050) <= 824007;
srom_1(39051) <= 593607;
srom_1(39052) <= 399760;
srom_1(39053) <= 243376;
srom_1(39054) <= 125187;
srom_1(39055) <= 45749;
srom_1(39056) <= 5433;
srom_1(39057) <= 4429;
srom_1(39058) <= 42741;
srom_1(39059) <= 120189;
srom_1(39060) <= 236411;
srom_1(39061) <= 390862;
srom_1(39062) <= 582817;
srom_1(39063) <= 811375;
srom_1(39064) <= 1075466;
srom_1(39065) <= 1373851;
srom_1(39066) <= 1705131;
srom_1(39067) <= 2067751;
srom_1(39068) <= 2460012;
srom_1(39069) <= 2880075;
srom_1(39070) <= 3325968;
srom_1(39071) <= 3795603;
srom_1(39072) <= 4286775;
srom_1(39073) <= 4797182;
srom_1(39074) <= 5324431;
srom_1(39075) <= 5866049;
srom_1(39076) <= 6419496;
srom_1(39077) <= 6982176;
srom_1(39078) <= 7551452;
srom_1(39079) <= 8124654;
srom_1(39080) <= 8699093;
srom_1(39081) <= 9272076;
srom_1(39082) <= 9840917;
srom_1(39083) <= 10402947;
srom_1(39084) <= 10955531;
srom_1(39085) <= 11496078;
srom_1(39086) <= 12022053;
srom_1(39087) <= 12530990;
srom_1(39088) <= 13020501;
srom_1(39089) <= 13488292;
srom_1(39090) <= 13932169;
srom_1(39091) <= 14350050;
srom_1(39092) <= 14739976;
srom_1(39093) <= 15100118;
srom_1(39094) <= 15428787;
srom_1(39095) <= 15724443;
srom_1(39096) <= 15985698;
srom_1(39097) <= 16211328;
srom_1(39098) <= 16400275;
srom_1(39099) <= 16551652;
srom_1(39100) <= 16664750;
srom_1(39101) <= 16739038;
srom_1(39102) <= 16774168;
srom_1(39103) <= 16769975;
srom_1(39104) <= 16726479;
srom_1(39105) <= 16643884;
srom_1(39106) <= 16522578;
srom_1(39107) <= 16363128;
srom_1(39108) <= 16166283;
srom_1(39109) <= 15932966;
srom_1(39110) <= 15664270;
srom_1(39111) <= 15361457;
srom_1(39112) <= 15025945;
srom_1(39113) <= 14659309;
srom_1(39114) <= 14263267;
srom_1(39115) <= 13839677;
srom_1(39116) <= 13390525;
srom_1(39117) <= 12917917;
srom_1(39118) <= 12424070;
srom_1(39119) <= 11911299;
srom_1(39120) <= 11382009;
srom_1(39121) <= 10838682;
srom_1(39122) <= 10283866;
srom_1(39123) <= 9720162;
srom_1(39124) <= 9150214;
srom_1(39125) <= 8576694;
srom_1(39126) <= 8002293;
srom_1(39127) <= 7429703;
srom_1(39128) <= 6861610;
srom_1(39129) <= 6300677;
srom_1(39130) <= 5749536;
srom_1(39131) <= 5210769;
srom_1(39132) <= 4686905;
srom_1(39133) <= 4180400;
srom_1(39134) <= 3693628;
srom_1(39135) <= 3228872;
srom_1(39136) <= 2788313;
srom_1(39137) <= 2374015;
srom_1(39138) <= 1987921;
srom_1(39139) <= 1631842;
srom_1(39140) <= 1307449;
srom_1(39141) <= 1016261;
srom_1(39142) <= 759645;
srom_1(39143) <= 538803;
srom_1(39144) <= 354772;
srom_1(39145) <= 208414;
srom_1(39146) <= 100417;
srom_1(39147) <= 31285;
srom_1(39148) <= 1343;
srom_1(39149) <= 10733;
srom_1(39150) <= 59409;
srom_1(39151) <= 147143;
srom_1(39152) <= 273525;
srom_1(39153) <= 437961;
srom_1(39154) <= 639680;
srom_1(39155) <= 877737;
srom_1(39156) <= 1151015;
srom_1(39157) <= 1458232;
srom_1(39158) <= 1797948;
srom_1(39159) <= 2168570;
srom_1(39160) <= 2568360;
srom_1(39161) <= 2995443;
srom_1(39162) <= 3447817;
srom_1(39163) <= 3923360;
srom_1(39164) <= 4419841;
srom_1(39165) <= 4934934;
srom_1(39166) <= 5466222;
srom_1(39167) <= 6011214;
srom_1(39168) <= 6567354;
srom_1(39169) <= 7132035;
srom_1(39170) <= 7702609;
srom_1(39171) <= 8276399;
srom_1(39172) <= 8850715;
srom_1(39173) <= 9422865;
srom_1(39174) <= 9990164;
srom_1(39175) <= 10549954;
srom_1(39176) <= 11099608;
srom_1(39177) <= 11636549;
srom_1(39178) <= 12158259;
srom_1(39179) <= 12662292;
srom_1(39180) <= 13146285;
srom_1(39181) <= 13607967;
srom_1(39182) <= 14045174;
srom_1(39183) <= 14455855;
srom_1(39184) <= 14838084;
srom_1(39185) <= 15190070;
srom_1(39186) <= 15510162;
srom_1(39187) <= 15796858;
srom_1(39188) <= 16048814;
srom_1(39189) <= 16264849;
srom_1(39190) <= 16443949;
srom_1(39191) <= 16585276;
srom_1(39192) <= 16688165;
srom_1(39193) <= 16752135;
srom_1(39194) <= 16776885;
srom_1(39195) <= 16762300;
srom_1(39196) <= 16708447;
srom_1(39197) <= 16615580;
srom_1(39198) <= 16484134;
srom_1(39199) <= 16314725;
srom_1(39200) <= 16108148;
srom_1(39201) <= 15865372;
srom_1(39202) <= 15587534;
srom_1(39203) <= 15275938;
srom_1(39204) <= 14932045;
srom_1(39205) <= 14557467;
srom_1(39206) <= 14153962;
srom_1(39207) <= 13723421;
srom_1(39208) <= 13267863;
srom_1(39209) <= 12789424;
srom_1(39210) <= 12290349;
srom_1(39211) <= 11772977;
srom_1(39212) <= 11239734;
srom_1(39213) <= 10693122;
srom_1(39214) <= 10135703;
srom_1(39215) <= 9570091;
srom_1(39216) <= 8998939;
srom_1(39217) <= 8424925;
srom_1(39218) <= 7850740;
srom_1(39219) <= 7279078;
srom_1(39220) <= 6712618;
srom_1(39221) <= 6154018;
srom_1(39222) <= 5605897;
srom_1(39223) <= 5070825;
srom_1(39224) <= 4551311;
srom_1(39225) <= 4049791;
srom_1(39226) <= 3568618;
srom_1(39227) <= 3110047;
srom_1(39228) <= 2676229;
srom_1(39229) <= 2269199;
srom_1(39230) <= 1890864;
srom_1(39231) <= 1543000;
srom_1(39232) <= 1227237;
srom_1(39233) <= 945056;
srom_1(39234) <= 697780;
srom_1(39235) <= 486570;
srom_1(39236) <= 312414;
srom_1(39237) <= 176131;
srom_1(39238) <= 78359;
srom_1(39239) <= 19557;
srom_1(39240) <= 0;
srom_1(39241) <= 19780;
srom_1(39242) <= 78804;
srom_1(39243) <= 176796;
srom_1(39244) <= 313295;
srom_1(39245) <= 487663;
srom_1(39246) <= 699081;
srom_1(39247) <= 946558;
srom_1(39248) <= 1228933;
srom_1(39249) <= 1544882;
srom_1(39250) <= 1892924;
srom_1(39251) <= 2271426;
srom_1(39252) <= 2678614;
srom_1(39253) <= 3112578;
srom_1(39254) <= 3571283;
srom_1(39255) <= 4052578;
srom_1(39256) <= 4554207;
srom_1(39257) <= 5073816;
srom_1(39258) <= 5608969;
srom_1(39259) <= 6157157;
srom_1(39260) <= 6715809;
srom_1(39261) <= 7282305;
srom_1(39262) <= 7853990;
srom_1(39263) <= 8428181;
srom_1(39264) <= 9002186;
srom_1(39265) <= 9573315;
srom_1(39266) <= 10138888;
srom_1(39267) <= 10696253;
srom_1(39268) <= 11242796;
srom_1(39269) <= 11775956;
srom_1(39270) <= 12293231;
srom_1(39271) <= 12792196;
srom_1(39272) <= 13270511;
srom_1(39273) <= 13725933;
srom_1(39274) <= 14156327;
srom_1(39275) <= 14559673;
srom_1(39276) <= 14934082;
srom_1(39277) <= 15277796;
srom_1(39278) <= 15589205;
srom_1(39279) <= 15866847;
srom_1(39280) <= 16109422;
srom_1(39281) <= 16315791;
srom_1(39282) <= 16484987;
srom_1(39283) <= 16616216;
srom_1(39284) <= 16708863;
srom_1(39285) <= 16762493;
srom_1(39286) <= 16776855;
srom_1(39287) <= 16751882;
srom_1(39288) <= 16687691;
srom_1(39289) <= 16584582;
srom_1(39290) <= 16443040;
srom_1(39291) <= 16263728;
srom_1(39292) <= 16047486;
srom_1(39293) <= 15795330;
srom_1(39294) <= 15508440;
srom_1(39295) <= 15188164;
srom_1(39296) <= 14836002;
srom_1(39297) <= 14453606;
srom_1(39298) <= 14042769;
srom_1(39299) <= 13605417;
srom_1(39300) <= 13143603;
srom_1(39301) <= 12659490;
srom_1(39302) <= 12155350;
srom_1(39303) <= 11633546;
srom_1(39304) <= 11096526;
srom_1(39305) <= 10546807;
srom_1(39306) <= 9986968;
srom_1(39307) <= 9419633;
srom_1(39308) <= 8847464;
srom_1(39309) <= 8273143;
srom_1(39310) <= 7699363;
srom_1(39311) <= 7128816;
srom_1(39312) <= 6564176;
srom_1(39313) <= 6008091;
srom_1(39314) <= 5463170;
srom_1(39315) <= 4931966;
srom_1(39316) <= 4416973;
srom_1(39317) <= 3920603;
srom_1(39318) <= 3445186;
srom_1(39319) <= 2992950;
srom_1(39320) <= 2566016;
srom_1(39321) <= 2166386;
srom_1(39322) <= 1795934;
srom_1(39323) <= 1456398;
srom_1(39324) <= 1149369;
srom_1(39325) <= 876288;
srom_1(39326) <= 638434;
srom_1(39327) <= 436923;
srom_1(39328) <= 272701;
srom_1(39329) <= 146537;
srom_1(39330) <= 59023;
srom_1(39331) <= 10569;
srom_1(39332) <= 1402;
srom_1(39333) <= 31566;
srom_1(39334) <= 100919;
srom_1(39335) <= 209136;
srom_1(39336) <= 355710;
srom_1(39337) <= 539952;
srom_1(39338) <= 760999;
srom_1(39339) <= 1017815;
srom_1(39340) <= 1309195;
srom_1(39341) <= 1633773;
srom_1(39342) <= 1990026;
srom_1(39343) <= 2376285;
srom_1(39344) <= 2790737;
srom_1(39345) <= 3231440;
srom_1(39346) <= 3696327;
srom_1(39347) <= 4183217;
srom_1(39348) <= 4689828;
srom_1(39349) <= 5213783;
srom_1(39350) <= 5752627;
srom_1(39351) <= 6303831;
srom_1(39352) <= 6864812;
srom_1(39353) <= 7432938;
srom_1(39354) <= 8005546;
srom_1(39355) <= 8579950;
srom_1(39356) <= 9153457;
srom_1(39357) <= 9723377;
srom_1(39358) <= 10287038;
srom_1(39359) <= 10841796;
srom_1(39360) <= 11385051;
srom_1(39361) <= 11914254;
srom_1(39362) <= 12426924;
srom_1(39363) <= 12920658;
srom_1(39364) <= 13393139;
srom_1(39365) <= 13842152;
srom_1(39366) <= 14265591;
srom_1(39367) <= 14661471;
srom_1(39368) <= 15027936;
srom_1(39369) <= 15363266;
srom_1(39370) <= 15665890;
srom_1(39371) <= 15934389;
srom_1(39372) <= 16167502;
srom_1(39373) <= 16364138;
srom_1(39374) <= 16523373;
srom_1(39375) <= 16644462;
srom_1(39376) <= 16726836;
srom_1(39377) <= 16770110;
srom_1(39378) <= 16774080;
srom_1(39379) <= 16738727;
srom_1(39380) <= 16664218;
srom_1(39381) <= 16550901;
srom_1(39382) <= 16399309;
srom_1(39383) <= 16210152;
srom_1(39384) <= 15984317;
srom_1(39385) <= 15722863;
srom_1(39386) <= 15427016;
srom_1(39387) <= 15098164;
srom_1(39388) <= 14737848;
srom_1(39389) <= 14347759;
srom_1(39390) <= 13929725;
srom_1(39391) <= 13485706;
srom_1(39392) <= 13017786;
srom_1(39393) <= 12528158;
srom_1(39394) <= 12019118;
srom_1(39395) <= 11493053;
srom_1(39396) <= 10952431;
srom_1(39397) <= 10399786;
srom_1(39398) <= 9837710;
srom_1(39399) <= 9268838;
srom_1(39400) <= 8695839;
srom_1(39401) <= 8121399;
srom_1(39402) <= 7548212;
srom_1(39403) <= 6978966;
srom_1(39404) <= 6416330;
srom_1(39405) <= 5862943;
srom_1(39406) <= 5321400;
srom_1(39407) <= 4794240;
srom_1(39408) <= 4283935;
srom_1(39409) <= 3792878;
srom_1(39410) <= 3323372;
srom_1(39411) <= 2877619;
srom_1(39412) <= 2457709;
srom_1(39413) <= 2065611;
srom_1(39414) <= 1703163;
srom_1(39415) <= 1372066;
srom_1(39416) <= 1073872;
srom_1(39417) <= 809979;
srom_1(39418) <= 581625;
srom_1(39419) <= 389880;
srom_1(39420) <= 235644;
srom_1(39421) <= 119641;
srom_1(39422) <= 42413;
srom_1(39423) <= 4324;
srom_1(39424) <= 5551;
srom_1(39425) <= 46089;
srom_1(39426) <= 125748;
srom_1(39427) <= 244155;
srom_1(39428) <= 400754;
srom_1(39429) <= 594810;
srom_1(39430) <= 825415;
srom_1(39431) <= 1091485;
srom_1(39432) <= 1391775;
srom_1(39433) <= 1724875;
srom_1(39434) <= 2089223;
srom_1(39435) <= 2483112;
srom_1(39436) <= 2904693;
srom_1(39437) <= 3351990;
srom_1(39438) <= 3822906;
srom_1(39439) <= 4315232;
srom_1(39440) <= 4826659;
srom_1(39441) <= 5354790;
srom_1(39442) <= 5897147;
srom_1(39443) <= 6451188;
srom_1(39444) <= 7014313;
srom_1(39445) <= 7583883;
srom_1(39446) <= 8157227;
srom_1(39447) <= 8731656;
srom_1(39448) <= 9304476;
srom_1(39449) <= 9873002;
srom_1(39450) <= 10434566;
srom_1(39451) <= 10986536;
srom_1(39452) <= 11526324;
srom_1(39453) <= 12051398;
srom_1(39454) <= 12559296;
srom_1(39455) <= 13047636;
srom_1(39456) <= 13514128;
srom_1(39457) <= 13956585;
srom_1(39458) <= 14372932;
srom_1(39459) <= 14761216;
srom_1(39460) <= 15119617;
srom_1(39461) <= 15446453;
srom_1(39462) <= 15740193;
srom_1(39463) <= 15999459;
srom_1(39464) <= 16223036;
srom_1(39465) <= 16409873;
srom_1(39466) <= 16559097;
srom_1(39467) <= 16670006;
srom_1(39468) <= 16742080;
srom_1(39469) <= 16774983;
srom_1(39470) <= 16768559;
srom_1(39471) <= 16722838;
srom_1(39472) <= 16638035;
srom_1(39473) <= 16514548;
srom_1(39474) <= 16352956;
srom_1(39475) <= 16154016;
srom_1(39476) <= 15918661;
srom_1(39477) <= 15647995;
srom_1(39478) <= 15343288;
srom_1(39479) <= 15005967;
srom_1(39480) <= 14637616;
srom_1(39481) <= 14239961;
srom_1(39482) <= 13814866;
srom_1(39483) <= 13364327;
srom_1(39484) <= 12890454;
srom_1(39485) <= 12395470;
srom_1(39486) <= 11881698;
srom_1(39487) <= 11351544;
srom_1(39488) <= 10807497;
srom_1(39489) <= 10252106;
srom_1(39490) <= 9687977;
srom_1(39491) <= 9117755;
srom_1(39492) <= 8544113;
srom_1(39493) <= 7969743;
srom_1(39494) <= 7397336;
srom_1(39495) <= 6829578;
srom_1(39496) <= 6269131;
srom_1(39497) <= 5718622;
srom_1(39498) <= 5180634;
srom_1(39499) <= 4657690;
srom_1(39500) <= 4152241;
srom_1(39501) <= 3666658;
srom_1(39502) <= 3203217;
srom_1(39503) <= 2764093;
srom_1(39504) <= 2351344;
srom_1(39505) <= 1966905;
srom_1(39506) <= 1612581;
srom_1(39507) <= 1290031;
srom_1(39508) <= 1000769;
srom_1(39509) <= 746151;
srom_1(39510) <= 527372;
srom_1(39511) <= 345456;
srom_1(39512) <= 201257;
srom_1(39513) <= 95452;
srom_1(39514) <= 28536;
srom_1(39515) <= 823;
srom_1(39516) <= 12444;
srom_1(39517) <= 63343;
srom_1(39518) <= 153283;
srom_1(39519) <= 281840;
srom_1(39520) <= 448413;
srom_1(39521) <= 652220;
srom_1(39522) <= 892306;
srom_1(39523) <= 1167545;
srom_1(39524) <= 1476645;
srom_1(39525) <= 1818158;
srom_1(39526) <= 2190483;
srom_1(39527) <= 2591872;
srom_1(39528) <= 3020444;
srom_1(39529) <= 3474190;
srom_1(39530) <= 3950981;
srom_1(39531) <= 4448581;
srom_1(39532) <= 4964657;
srom_1(39533) <= 5496790;
srom_1(39534) <= 6042483;
srom_1(39535) <= 6599178;
srom_1(39536) <= 7164265;
srom_1(39537) <= 7735092;
srom_1(39538) <= 8308985;
srom_1(39539) <= 8883250;
srom_1(39540) <= 9455196;
srom_1(39541) <= 10022141;
srom_1(39542) <= 10581425;
srom_1(39543) <= 11130426;
srom_1(39544) <= 11666570;
srom_1(39545) <= 12187343;
srom_1(39546) <= 12690302;
srom_1(39547) <= 13173089;
srom_1(39548) <= 13633439;
srom_1(39549) <= 14069195;
srom_1(39550) <= 14478313;
srom_1(39551) <= 14858874;
srom_1(39552) <= 15209093;
srom_1(39553) <= 15527330;
srom_1(39554) <= 15812090;
srom_1(39555) <= 16062038;
srom_1(39556) <= 16276004;
srom_1(39557) <= 16452983;
srom_1(39558) <= 16592145;
srom_1(39559) <= 16692838;
srom_1(39560) <= 16754589;
srom_1(39561) <= 16777110;
srom_1(39562) <= 16760294;
srom_1(39563) <= 16704220;
srom_1(39564) <= 16609152;
srom_1(39565) <= 16475534;
srom_1(39566) <= 16303994;
srom_1(39567) <= 16095337;
srom_1(39568) <= 15850539;
srom_1(39569) <= 15570750;
srom_1(39570) <= 15257282;
srom_1(39571) <= 14911604;
srom_1(39572) <= 14535338;
srom_1(39573) <= 14130247;
srom_1(39574) <= 13698232;
srom_1(39575) <= 13241318;
srom_1(39576) <= 12761648;
srom_1(39577) <= 12261471;
srom_1(39578) <= 11743133;
srom_1(39579) <= 11209065;
srom_1(39580) <= 10661771;
srom_1(39581) <= 10103816;
srom_1(39582) <= 9537819;
srom_1(39583) <= 8966433;
srom_1(39584) <= 8392337;
srom_1(39585) <= 7818223;
srom_1(39586) <= 7246785;
srom_1(39587) <= 6680700;
srom_1(39588) <= 6122625;
srom_1(39589) <= 5575176;
srom_1(39590) <= 5040919;
srom_1(39591) <= 4522361;
srom_1(39592) <= 4021934;
srom_1(39593) <= 3541983;
srom_1(39594) <= 3084760;
srom_1(39595) <= 2652408;
srom_1(39596) <= 2246955;
srom_1(39597) <= 1870303;
srom_1(39598) <= 1524217;
srom_1(39599) <= 1210320;
srom_1(39600) <= 930085;
srom_1(39601) <= 684826;
srom_1(39602) <= 475692;
srom_1(39603) <= 303665;
srom_1(39604) <= 169550;
srom_1(39605) <= 73978;
srom_1(39606) <= 17396;
srom_1(39607) <= 69;
srom_1(39608) <= 22079;
srom_1(39609) <= 83323;
srom_1(39610) <= 183513;
srom_1(39611) <= 322179;
srom_1(39612) <= 498672;
srom_1(39613) <= 712163;
srom_1(39614) <= 961652;
srom_1(39615) <= 1245968;
srom_1(39616) <= 1563779;
srom_1(39617) <= 1913593;
srom_1(39618) <= 2293771;
srom_1(39619) <= 2702530;
srom_1(39620) <= 3137953;
srom_1(39621) <= 3597998;
srom_1(39622) <= 4080508;
srom_1(39623) <= 4583220;
srom_1(39624) <= 5103776;
srom_1(39625) <= 5639737;
srom_1(39626) <= 6188588;
srom_1(39627) <= 6747755;
srom_1(39628) <= 7314617;
srom_1(39629) <= 7886515;
srom_1(39630) <= 8460768;
srom_1(39631) <= 9034682;
srom_1(39632) <= 9605567;
srom_1(39633) <= 10170745;
srom_1(39634) <= 10727566;
srom_1(39635) <= 11273418;
srom_1(39636) <= 11805743;
srom_1(39637) <= 12322044;
srom_1(39638) <= 12819899;
srom_1(39639) <= 13296975;
srom_1(39640) <= 13751033;
srom_1(39641) <= 14179946;
srom_1(39642) <= 14581700;
srom_1(39643) <= 14954414;
srom_1(39644) <= 15296337;
srom_1(39645) <= 15605869;
srom_1(39646) <= 15881555;
srom_1(39647) <= 16122105;
srom_1(39648) <= 16326390;
srom_1(39649) <= 16493452;
srom_1(39650) <= 16622507;
srom_1(39651) <= 16712951;
srom_1(39652) <= 16764360;
srom_1(39653) <= 16776491;
srom_1(39654) <= 16749289;
srom_1(39655) <= 16682880;
srom_1(39656) <= 16577577;
srom_1(39657) <= 16433873;
srom_1(39658) <= 16252442;
srom_1(39659) <= 16034135;
srom_1(39660) <= 15779975;
srom_1(39661) <= 15491155;
srom_1(39662) <= 15169028;
srom_1(39663) <= 14815105;
srom_1(39664) <= 14431047;
srom_1(39665) <= 14018653;
srom_1(39666) <= 13579858;
srom_1(39667) <= 13116720;
srom_1(39668) <= 12631410;
srom_1(39669) <= 12126204;
srom_1(39670) <= 11603471;
srom_1(39671) <= 11065662;
srom_1(39672) <= 10515300;
srom_1(39673) <= 9954965;
srom_1(39674) <= 9387285;
srom_1(39675) <= 8814922;
srom_1(39676) <= 8240559;
srom_1(39677) <= 7666891;
srom_1(39678) <= 7096607;
srom_1(39679) <= 6532382;
srom_1(39680) <= 5976861;
srom_1(39681) <= 5432650;
srom_1(39682) <= 4902300;
srom_1(39683) <= 4388299;
srom_1(39684) <= 3893056;
srom_1(39685) <= 3418895;
srom_1(39686) <= 2968038;
srom_1(39687) <= 2542601;
srom_1(39688) <= 2144577;
srom_1(39689) <= 1775834;
srom_1(39690) <= 1438100;
srom_1(39691) <= 1132959;
srom_1(39692) <= 861843;
srom_1(39693) <= 626023;
srom_1(39694) <= 426603;
srom_1(39695) <= 264521;
srom_1(39696) <= 140535;
srom_1(39697) <= 55227;
srom_1(39698) <= 8997;
srom_1(39699) <= 2062;
srom_1(39700) <= 34454;
srom_1(39701) <= 106022;
srom_1(39702) <= 216429;
srom_1(39703) <= 365159;
srom_1(39704) <= 551514;
srom_1(39705) <= 774619;
srom_1(39706) <= 1033429;
srom_1(39707) <= 1326730;
srom_1(39708) <= 1653147;
srom_1(39709) <= 2011148;
srom_1(39710) <= 2399055;
srom_1(39711) <= 2815050;
srom_1(39712) <= 3257181;
srom_1(39713) <= 3723375;
srom_1(39714) <= 4211445;
srom_1(39715) <= 4719104;
srom_1(39716) <= 5243971;
srom_1(39717) <= 5783584;
srom_1(39718) <= 6335412;
srom_1(39719) <= 6896869;
srom_1(39720) <= 7465321;
srom_1(39721) <= 8038102;
srom_1(39722) <= 8612528;
srom_1(39723) <= 9185903;
srom_1(39724) <= 9755539;
srom_1(39725) <= 10318766;
srom_1(39726) <= 10872941;
srom_1(39727) <= 11415466;
srom_1(39728) <= 11943797;
srom_1(39729) <= 12455457;
srom_1(39730) <= 12948046;
srom_1(39731) <= 13419254;
srom_1(39732) <= 13866872;
srom_1(39733) <= 14288800;
srom_1(39734) <= 14683060;
srom_1(39735) <= 15047804;
srom_1(39736) <= 15381320;
srom_1(39737) <= 15682045;
srom_1(39738) <= 15948568;
srom_1(39739) <= 16179640;
srom_1(39740) <= 16374178;
srom_1(39741) <= 16531268;
srom_1(39742) <= 16650174;
srom_1(39743) <= 16730340;
srom_1(39744) <= 16771387;
srom_1(39745) <= 16773126;
srom_1(39746) <= 16735546;
srom_1(39747) <= 16658825;
srom_1(39748) <= 16543321;
srom_1(39749) <= 16389578;
srom_1(39750) <= 16198315;
srom_1(39751) <= 15970430;
srom_1(39752) <= 15706991;
srom_1(39753) <= 15409233;
srom_1(39754) <= 15078554;
srom_1(39755) <= 14716503;
srom_1(39756) <= 14324778;
srom_1(39757) <= 13905217;
srom_1(39758) <= 13459786;
srom_1(39759) <= 12990575;
srom_1(39760) <= 12499783;
srom_1(39761) <= 11989713;
srom_1(39762) <= 11462756;
srom_1(39763) <= 10921383;
srom_1(39764) <= 10368133;
srom_1(39765) <= 9805601;
srom_1(39766) <= 9236424;
srom_1(39767) <= 8663271;
srom_1(39768) <= 8088830;
srom_1(39769) <= 7515795;
srom_1(39770) <= 6946852;
srom_1(39771) <= 6384671;
srom_1(39772) <= 5831887;
srom_1(39773) <= 5291092;
srom_1(39774) <= 4764822;
srom_1(39775) <= 4255546;
srom_1(39776) <= 3765651;
srom_1(39777) <= 3297434;
srom_1(39778) <= 2853092;
srom_1(39779) <= 2434708;
srom_1(39780) <= 2044243;
srom_1(39781) <= 1683530;
srom_1(39782) <= 1354259;
srom_1(39783) <= 1057974;
srom_1(39784) <= 796065;
srom_1(39785) <= 569761;
srom_1(39786) <= 380121;
srom_1(39787) <= 228036;
srom_1(39788) <= 114219;
srom_1(39789) <= 39203;
srom_1(39790) <= 3341;
srom_1(39791) <= 6799;
srom_1(39792) <= 49563;
srom_1(39793) <= 131432;
srom_1(39794) <= 252021;
srom_1(39795) <= 410766;
srom_1(39796) <= 606922;
srom_1(39797) <= 839568;
srom_1(39798) <= 1107614;
srom_1(39799) <= 1409804;
srom_1(39800) <= 1744720;
srom_1(39801) <= 2110791;
srom_1(39802) <= 2506300;
srom_1(39803) <= 2929394;
srom_1(39804) <= 3378089;
srom_1(39805) <= 3850279;
srom_1(39806) <= 4343751;
srom_1(39807) <= 4856190;
srom_1(39808) <= 5385195;
srom_1(39809) <= 5928283;
srom_1(39810) <= 6482909;
srom_1(39811) <= 7046471;
srom_1(39812) <= 7616327;
srom_1(39813) <= 8189804;
srom_1(39814) <= 8764214;
srom_1(39815) <= 9336862;
srom_1(39816) <= 9905064;
srom_1(39817) <= 10466154;
srom_1(39818) <= 11017502;
srom_1(39819) <= 11556523;
srom_1(39820) <= 12080688;
srom_1(39821) <= 12587539;
srom_1(39822) <= 13074700;
srom_1(39823) <= 13539887;
srom_1(39824) <= 13980917;
srom_1(39825) <= 14395723;
srom_1(39826) <= 14782360;
srom_1(39827) <= 15139014;
srom_1(39828) <= 15464013;
srom_1(39829) <= 15755833;
srom_1(39830) <= 16013106;
srom_1(39831) <= 16234625;
srom_1(39832) <= 16419351;
srom_1(39833) <= 16566418;
srom_1(39834) <= 16675136;
srom_1(39835) <= 16744997;
srom_1(39836) <= 16775671;
srom_1(39837) <= 16767015;
srom_1(39838) <= 16719071;
srom_1(39839) <= 16632061;
srom_1(39840) <= 16506396;
srom_1(39841) <= 16342663;
srom_1(39842) <= 16141631;
srom_1(39843) <= 15904242;
srom_1(39844) <= 15631610;
srom_1(39845) <= 15325013;
srom_1(39846) <= 14985889;
srom_1(39847) <= 14615828;
srom_1(39848) <= 14216566;
srom_1(39849) <= 13789974;
srom_1(39850) <= 13338053;
srom_1(39851) <= 12862922;
srom_1(39852) <= 12366810;
srom_1(39853) <= 11852043;
srom_1(39854) <= 11321035;
srom_1(39855) <= 10776275;
srom_1(39856) <= 10220319;
srom_1(39857) <= 9655773;
srom_1(39858) <= 9085285;
srom_1(39859) <= 8511530;
srom_1(39860) <= 7937199;
srom_1(39861) <= 7364984;
srom_1(39862) <= 6797570;
srom_1(39863) <= 6237616;
srom_1(39864) <= 5687750;
srom_1(39865) <= 5150548;
srom_1(39866) <= 4628531;
srom_1(39867) <= 4124146;
srom_1(39868) <= 3639759;
srom_1(39869) <= 3177640;
srom_1(39870) <= 2739958;
srom_1(39871) <= 2328764;
srom_1(39872) <= 1945987;
srom_1(39873) <= 1593421;
srom_1(39874) <= 1272721;
srom_1(39875) <= 985389;
srom_1(39876) <= 732773;
srom_1(39877) <= 516059;
srom_1(39878) <= 336261;
srom_1(39879) <= 194224;
srom_1(39880) <= 90612;
srom_1(39881) <= 25913;
srom_1(39882) <= 430;
srom_1(39883) <= 14282;
srom_1(39884) <= 67403;
srom_1(39885) <= 159546;
srom_1(39886) <= 290277;
srom_1(39887) <= 458985;
srom_1(39888) <= 664877;
srom_1(39889) <= 906988;
srom_1(39890) <= 1184184;
srom_1(39891) <= 1495163;
srom_1(39892) <= 1838468;
srom_1(39893) <= 2212489;
srom_1(39894) <= 2615471;
srom_1(39895) <= 3045526;
srom_1(39896) <= 3500637;
srom_1(39897) <= 3978669;
srom_1(39898) <= 4477380;
srom_1(39899) <= 4994433;
srom_1(39900) <= 5527402;
srom_1(39901) <= 6073788;
srom_1(39902) <= 6631030;
srom_1(39903) <= 7196513;
srom_1(39904) <= 7767586;
srom_1(39905) <= 8341571;
srom_1(39906) <= 8915777;
srom_1(39907) <= 9487511;
srom_1(39908) <= 10054092;
srom_1(39909) <= 10612863;
srom_1(39910) <= 11161203;
srom_1(39911) <= 11696542;
srom_1(39912) <= 12216369;
srom_1(39913) <= 12718246;
srom_1(39914) <= 13199820;
srom_1(39915) <= 13658832;
srom_1(39916) <= 14093131;
srom_1(39917) <= 14500679;
srom_1(39918) <= 14879566;
srom_1(39919) <= 15228014;
srom_1(39920) <= 15544390;
srom_1(39921) <= 15827209;
srom_1(39922) <= 16075147;
srom_1(39923) <= 16287040;
srom_1(39924) <= 16461894;
srom_1(39925) <= 16598890;
srom_1(39926) <= 16697386;
srom_1(39927) <= 16756918;
srom_1(39928) <= 16777209;
srom_1(39929) <= 16758162;
srom_1(39930) <= 16699868;
srom_1(39931) <= 16602599;
srom_1(39932) <= 16466813;
srom_1(39933) <= 16293144;
srom_1(39934) <= 16082409;
srom_1(39935) <= 15835595;
srom_1(39936) <= 15553859;
srom_1(39937) <= 15238523;
srom_1(39938) <= 14891065;
srom_1(39939) <= 14513115;
srom_1(39940) <= 14106445;
srom_1(39941) <= 13672962;
srom_1(39942) <= 13214700;
srom_1(39943) <= 12733805;
srom_1(39944) <= 12232535;
srom_1(39945) <= 11713239;
srom_1(39946) <= 11178353;
srom_1(39947) <= 10630385;
srom_1(39948) <= 10071904;
srom_1(39949) <= 9505530;
srom_1(39950) <= 8933918;
srom_1(39951) <= 8359749;
srom_1(39952) <= 7785715;
srom_1(39953) <= 7214509;
srom_1(39954) <= 6648808;
srom_1(39955) <= 6091266;
srom_1(39956) <= 5544497;
srom_1(39957) <= 5011064;
srom_1(39958) <= 4493470;
srom_1(39959) <= 3994142;
srom_1(39960) <= 3515421;
srom_1(39961) <= 3059552;
srom_1(39962) <= 2628673;
srom_1(39963) <= 2224804;
srom_1(39964) <= 1849839;
srom_1(39965) <= 1505537;
srom_1(39966) <= 1193512;
srom_1(39967) <= 915227;
srom_1(39968) <= 671988;
srom_1(39969) <= 464934;
srom_1(39970) <= 295037;
srom_1(39971) <= 163094;
srom_1(39972) <= 69723;
srom_1(39973) <= 15361;
srom_1(39974) <= 265;
srom_1(39975) <= 24505;
srom_1(39976) <= 87967;
srom_1(39977) <= 190354;
srom_1(39978) <= 331185;
srom_1(39979) <= 509800;
srom_1(39980) <= 725361;
srom_1(39981) <= 976858;
srom_1(39982) <= 1263111;
srom_1(39983) <= 1582778;
srom_1(39984) <= 1934360;
srom_1(39985) <= 2316208;
srom_1(39986) <= 2726532;
srom_1(39987) <= 3163407;
srom_1(39988) <= 3624785;
srom_1(39989) <= 4108502;
srom_1(39990) <= 4612290;
srom_1(39991) <= 5133787;
srom_1(39992) <= 5670546;
srom_1(39993) <= 6220051;
srom_1(39994) <= 6779726;
srom_1(39995) <= 7346945;
srom_1(39996) <= 7919048;
srom_1(39997) <= 8493354;
srom_1(39998) <= 9067168;
srom_1(39999) <= 9637801;
srom_1(40000) <= 10202575;
srom_1(40001) <= 10758843;
srom_1(40002) <= 11303997;
srom_1(40003) <= 11835479;
srom_1(40004) <= 12350797;
srom_1(40005) <= 12847536;
srom_1(40006) <= 13323365;
srom_1(40007) <= 13776053;
srom_1(40008) <= 14203477;
srom_1(40009) <= 14603634;
srom_1(40010) <= 14974646;
srom_1(40011) <= 15314774;
srom_1(40012) <= 15622423;
srom_1(40013) <= 15896150;
srom_1(40014) <= 16134672;
srom_1(40015) <= 16336870;
srom_1(40016) <= 16501795;
srom_1(40017) <= 16628675;
srom_1(40018) <= 16716914;
srom_1(40019) <= 16766100;
srom_1(40020) <= 16776000;
srom_1(40021) <= 16746569;
srom_1(40022) <= 16677944;
srom_1(40023) <= 16570448;
srom_1(40024) <= 16424585;
srom_1(40025) <= 16241038;
srom_1(40026) <= 16020668;
srom_1(40027) <= 15764509;
srom_1(40028) <= 15473761;
srom_1(40029) <= 15149789;
srom_1(40030) <= 14794112;
srom_1(40031) <= 14408397;
srom_1(40032) <= 13994453;
srom_1(40033) <= 13554221;
srom_1(40034) <= 13089766;
srom_1(40035) <= 12603266;
srom_1(40036) <= 12097001;
srom_1(40037) <= 11573347;
srom_1(40038) <= 11034758;
srom_1(40039) <= 10483761;
srom_1(40040) <= 9922939;
srom_1(40041) <= 9354921;
srom_1(40042) <= 8782373;
srom_1(40043) <= 8207978;
srom_1(40044) <= 7634429;
srom_1(40045) <= 7064418;
srom_1(40046) <= 6500616;
srom_1(40047) <= 5945667;
srom_1(40048) <= 5402175;
srom_1(40049) <= 4872686;
srom_1(40050) <= 4359685;
srom_1(40051) <= 3865577;
srom_1(40052) <= 3392679;
srom_1(40053) <= 2943209;
srom_1(40054) <= 2519274;
srom_1(40055) <= 2122862;
srom_1(40056) <= 1755833;
srom_1(40057) <= 1419907;
srom_1(40058) <= 1116659;
srom_1(40059) <= 847512;
srom_1(40060) <= 613728;
srom_1(40061) <= 416403;
srom_1(40062) <= 256463;
srom_1(40063) <= 134657;
srom_1(40064) <= 51556;
srom_1(40065) <= 7551;
srom_1(40066) <= 2847;
srom_1(40067) <= 37467;
srom_1(40068) <= 111249;
srom_1(40069) <= 223846;
srom_1(40070) <= 374730;
srom_1(40071) <= 563194;
srom_1(40072) <= 788354;
srom_1(40073) <= 1049154;
srom_1(40074) <= 1344372;
srom_1(40075) <= 1672622;
srom_1(40076) <= 2032366;
srom_1(40077) <= 2421916;
srom_1(40078) <= 2839447;
srom_1(40079) <= 3282999;
srom_1(40080) <= 3750493;
srom_1(40081) <= 4239737;
srom_1(40082) <= 4748437;
srom_1(40083) <= 5274206;
srom_1(40084) <= 5814580;
srom_1(40085) <= 6367024;
srom_1(40086) <= 6928948;
srom_1(40087) <= 7497718;
srom_1(40088) <= 8070664;
srom_1(40089) <= 8645102;
srom_1(40090) <= 9218337;
srom_1(40091) <= 9787681;
srom_1(40092) <= 10350464;
srom_1(40093) <= 10904048;
srom_1(40094) <= 11445836;
srom_1(40095) <= 11973287;
srom_1(40096) <= 12483928;
srom_1(40097) <= 12975366;
srom_1(40098) <= 13445294;
srom_1(40099) <= 13891509;
srom_1(40100) <= 14311920;
srom_1(40101) <= 14704554;
srom_1(40102) <= 15067571;
srom_1(40103) <= 15399268;
srom_1(40104) <= 15698089;
srom_1(40105) <= 15962634;
srom_1(40106) <= 16191661;
srom_1(40107) <= 16384097;
srom_1(40108) <= 16539040;
srom_1(40109) <= 16655762;
srom_1(40110) <= 16733717;
srom_1(40111) <= 16772539;
srom_1(40112) <= 16772045;
srom_1(40113) <= 16732239;
srom_1(40114) <= 16653307;
srom_1(40115) <= 16535618;
srom_1(40116) <= 16379726;
srom_1(40117) <= 16186360;
srom_1(40118) <= 15956428;
srom_1(40119) <= 15691008;
srom_1(40120) <= 15391344;
srom_1(40121) <= 15058843;
srom_1(40122) <= 14695062;
srom_1(40123) <= 14301708;
srom_1(40124) <= 13880625;
srom_1(40125) <= 13433789;
srom_1(40126) <= 12963294;
srom_1(40127) <= 12471346;
srom_1(40128) <= 11960254;
srom_1(40129) <= 11432412;
srom_1(40130) <= 10890297;
srom_1(40131) <= 10336451;
srom_1(40132) <= 9773471;
srom_1(40133) <= 9203996;
srom_1(40134) <= 8630698;
srom_1(40135) <= 8056265;
srom_1(40136) <= 7483390;
srom_1(40137) <= 6914760;
srom_1(40138) <= 6353042;
srom_1(40139) <= 5800869;
srom_1(40140) <= 5260830;
srom_1(40141) <= 4735459;
srom_1(40142) <= 4227219;
srom_1(40143) <= 3738493;
srom_1(40144) <= 3271573;
srom_1(40145) <= 2828648;
srom_1(40146) <= 2411796;
srom_1(40147) <= 2022972;
srom_1(40148) <= 1663998;
srom_1(40149) <= 1336558;
srom_1(40150) <= 1042187;
srom_1(40151) <= 782266;
srom_1(40152) <= 558015;
srom_1(40153) <= 370483;
srom_1(40154) <= 220551;
srom_1(40155) <= 108922;
srom_1(40156) <= 36119;
srom_1(40157) <= 2484;
srom_1(40158) <= 8175;
srom_1(40159) <= 53164;
srom_1(40160) <= 137240;
srom_1(40161) <= 260011;
srom_1(40162) <= 420899;
srom_1(40163) <= 619150;
srom_1(40164) <= 853835;
srom_1(40165) <= 1123853;
srom_1(40166) <= 1427939;
srom_1(40167) <= 1764665;
srom_1(40168) <= 2132453;
srom_1(40169) <= 2529578;
srom_1(40170) <= 2954178;
srom_1(40171) <= 3404262;
srom_1(40172) <= 3877720;
srom_1(40173) <= 4372330;
srom_1(40174) <= 4885775;
srom_1(40175) <= 5415645;
srom_1(40176) <= 5959456;
srom_1(40177) <= 6514659;
srom_1(40178) <= 7078649;
srom_1(40179) <= 7648782;
srom_1(40180) <= 8222384;
srom_1(40181) <= 8796766;
srom_1(40182) <= 9369234;
srom_1(40183) <= 9937103;
srom_1(40184) <= 10497711;
srom_1(40185) <= 11048429;
srom_1(40186) <= 11586673;
srom_1(40187) <= 12109921;
srom_1(40188) <= 12615719;
srom_1(40189) <= 13101694;
srom_1(40190) <= 13565567;
srom_1(40191) <= 14005164;
srom_1(40192) <= 14418424;
srom_1(40193) <= 14803407;
srom_1(40194) <= 15158309;
srom_1(40195) <= 15481466;
srom_1(40196) <= 15771361;
srom_1(40197) <= 16026637;
srom_1(40198) <= 16246095;
srom_1(40199) <= 16428707;
srom_1(40200) <= 16573616;
srom_1(40201) <= 16680142;
srom_1(40202) <= 16747787;
srom_1(40203) <= 16776233;
srom_1(40204) <= 16765346;
srom_1(40205) <= 16715178;
srom_1(40206) <= 16625963;
srom_1(40207) <= 16498121;
srom_1(40208) <= 16332251;
srom_1(40209) <= 16129130;
srom_1(40210) <= 15889711;
srom_1(40211) <= 15615116;
srom_1(40212) <= 15306635;
srom_1(40213) <= 14965712;
srom_1(40214) <= 14593947;
srom_1(40215) <= 14193083;
srom_1(40216) <= 13765000;
srom_1(40217) <= 13311705;
srom_1(40218) <= 12835323;
srom_1(40219) <= 12338090;
srom_1(40220) <= 11822336;
srom_1(40221) <= 11290481;
srom_1(40222) <= 10745017;
srom_1(40223) <= 10188504;
srom_1(40224) <= 9623550;
srom_1(40225) <= 9052805;
srom_1(40226) <= 8478945;
srom_1(40227) <= 7904662;
srom_1(40228) <= 7332648;
srom_1(40229) <= 6765586;
srom_1(40230) <= 6206134;
srom_1(40231) <= 5656917;
srom_1(40232) <= 5120510;
srom_1(40233) <= 4599429;
srom_1(40234) <= 4096115;
srom_1(40235) <= 3612931;
srom_1(40236) <= 3152142;
srom_1(40237) <= 2715908;
srom_1(40238) <= 2306276;
srom_1(40239) <= 1925165;
srom_1(40240) <= 1574364;
srom_1(40241) <= 1255517;
srom_1(40242) <= 970120;
srom_1(40243) <= 719511;
srom_1(40244) <= 504864;
srom_1(40245) <= 327188;
srom_1(40246) <= 187314;
srom_1(40247) <= 85898;
srom_1(40248) <= 23417;
srom_1(40249) <= 163;
srom_1(40250) <= 16246;
srom_1(40251) <= 71589;
srom_1(40252) <= 165933;
srom_1(40253) <= 298837;
srom_1(40254) <= 469676;
srom_1(40255) <= 677650;
srom_1(40256) <= 921783;
srom_1(40257) <= 1200931;
srom_1(40258) <= 1513784;
srom_1(40259) <= 1858876;
srom_1(40260) <= 2234588;
srom_1(40261) <= 2639158;
srom_1(40262) <= 3070689;
srom_1(40263) <= 3527157;
srom_1(40264) <= 4006423;
srom_1(40265) <= 4506238;
srom_1(40266) <= 5024260;
srom_1(40267) <= 5558057;
srom_1(40268) <= 6105128;
srom_1(40269) <= 6662907;
srom_1(40270) <= 7228779;
srom_1(40271) <= 7800089;
srom_1(40272) <= 8374159;
srom_1(40273) <= 8948297;
srom_1(40274) <= 9519810;
srom_1(40275) <= 10086019;
srom_1(40276) <= 10644268;
srom_1(40277) <= 11191939;
srom_1(40278) <= 11726464;
srom_1(40279) <= 12245337;
srom_1(40280) <= 12746125;
srom_1(40281) <= 13226479;
srom_1(40282) <= 13684146;
srom_1(40283) <= 14116981;
srom_1(40284) <= 14522953;
srom_1(40285) <= 14900159;
srom_1(40286) <= 15246831;
srom_1(40287) <= 15561341;
srom_1(40288) <= 15842217;
srom_1(40289) <= 16088140;
srom_1(40290) <= 16297957;
srom_1(40291) <= 16470684;
srom_1(40292) <= 16605512;
srom_1(40293) <= 16701808;
srom_1(40294) <= 16759120;
srom_1(40295) <= 16777181;
srom_1(40296) <= 16755904;
srom_1(40297) <= 16695390;
srom_1(40298) <= 16595923;
srom_1(40299) <= 16457969;
srom_1(40300) <= 16282175;
srom_1(40301) <= 16069365;
srom_1(40302) <= 15820537;
srom_1(40303) <= 15536859;
srom_1(40304) <= 15219660;
srom_1(40305) <= 14870428;
srom_1(40306) <= 14490800;
srom_1(40307) <= 14082557;
srom_1(40308) <= 13647614;
srom_1(40309) <= 13188009;
srom_1(40310) <= 12705897;
srom_1(40311) <= 12203541;
srom_1(40312) <= 11683295;
srom_1(40313) <= 11147599;
srom_1(40314) <= 10598966;
srom_1(40315) <= 10039967;
srom_1(40316) <= 9473224;
srom_1(40317) <= 8901395;
srom_1(40318) <= 8327162;
srom_1(40319) <= 7753216;
srom_1(40320) <= 7182251;
srom_1(40321) <= 6616942;
srom_1(40322) <= 6059941;
srom_1(40323) <= 5513860;
srom_1(40324) <= 4981260;
srom_1(40325) <= 4464638;
srom_1(40326) <= 3966417;
srom_1(40327) <= 3488933;
srom_1(40328) <= 3034425;
srom_1(40329) <= 2605025;
srom_1(40330) <= 2202746;
srom_1(40331) <= 1829475;
srom_1(40332) <= 1486962;
srom_1(40333) <= 1176813;
srom_1(40334) <= 900482;
srom_1(40335) <= 659266;
srom_1(40336) <= 454295;
srom_1(40337) <= 286531;
srom_1(40338) <= 156761;
srom_1(40339) <= 65592;
srom_1(40340) <= 13453;
srom_1(40341) <= 588;
srom_1(40342) <= 27058;
srom_1(40343) <= 92737;
srom_1(40344) <= 197318;
srom_1(40345) <= 340312;
srom_1(40346) <= 521046;
srom_1(40347) <= 738675;
srom_1(40348) <= 992176;
srom_1(40349) <= 1280362;
srom_1(40350) <= 1601881;
srom_1(40351) <= 1955225;
srom_1(40352) <= 2338737;
srom_1(40353) <= 2750620;
srom_1(40354) <= 3188940;
srom_1(40355) <= 3651644;
srom_1(40356) <= 4136561;
srom_1(40357) <= 4641418;
srom_1(40358) <= 5163846;
srom_1(40359) <= 5701396;
srom_1(40360) <= 6251548;
srom_1(40361) <= 6811721;
srom_1(40362) <= 7379288;
srom_1(40363) <= 7951589;
srom_1(40364) <= 8525938;
srom_1(40365) <= 9099644;
srom_1(40366) <= 9670016;
srom_1(40367) <= 10234378;
srom_1(40368) <= 10790085;
srom_1(40369) <= 11334531;
srom_1(40370) <= 11865162;
srom_1(40371) <= 12379491;
srom_1(40372) <= 12875105;
srom_1(40373) <= 13349680;
srom_1(40374) <= 13800991;
srom_1(40375) <= 14226921;
srom_1(40376) <= 14625474;
srom_1(40377) <= 14994780;
srom_1(40378) <= 15333107;
srom_1(40379) <= 15638869;
srom_1(40380) <= 15910632;
srom_1(40381) <= 16147122;
srom_1(40382) <= 16347229;
srom_1(40383) <= 16510016;
srom_1(40384) <= 16634718;
srom_1(40385) <= 16720752;
srom_1(40386) <= 16767713;
srom_1(40387) <= 16775382;
srom_1(40388) <= 16743723;
srom_1(40389) <= 16672883;
srom_1(40390) <= 16563196;
srom_1(40391) <= 16415175;
srom_1(40392) <= 16229515;
srom_1(40393) <= 16007086;
srom_1(40394) <= 15748931;
srom_1(40395) <= 15456261;
srom_1(40396) <= 15130449;
srom_1(40397) <= 14773022;
srom_1(40398) <= 14385656;
srom_1(40399) <= 13970168;
srom_1(40400) <= 13528506;
srom_1(40401) <= 13062741;
srom_1(40402) <= 12575058;
srom_1(40403) <= 12067743;
srom_1(40404) <= 11543175;
srom_1(40405) <= 11003815;
srom_1(40406) <= 10452190;
srom_1(40407) <= 9890889;
srom_1(40408) <= 9322543;
srom_1(40409) <= 8749818;
srom_1(40410) <= 8175399;
srom_1(40411) <= 7601979;
srom_1(40412) <= 7032249;
srom_1(40413) <= 6468879;
srom_1(40414) <= 5914511;
srom_1(40415) <= 5371745;
srom_1(40416) <= 4843126;
srom_1(40417) <= 4331133;
srom_1(40418) <= 3838166;
srom_1(40419) <= 3366539;
srom_1(40420) <= 2918462;
srom_1(40421) <= 2496036;
srom_1(40422) <= 2101242;
srom_1(40423) <= 1735932;
srom_1(40424) <= 1401819;
srom_1(40425) <= 1100469;
srom_1(40426) <= 833295;
srom_1(40427) <= 601552;
srom_1(40428) <= 406324;
srom_1(40429) <= 248528;
srom_1(40430) <= 128903;
srom_1(40431) <= 48012;
srom_1(40432) <= 6232;
srom_1(40433) <= 3760;
srom_1(40434) <= 40607;
srom_1(40435) <= 116601;
srom_1(40436) <= 231385;
srom_1(40437) <= 384422;
srom_1(40438) <= 574992;
srom_1(40439) <= 802204;
srom_1(40440) <= 1064990;
srom_1(40441) <= 1362120;
srom_1(40442) <= 1692199;
srom_1(40443) <= 2053680;
srom_1(40444) <= 2444868;
srom_1(40445) <= 2863927;
srom_1(40446) <= 3308894;
srom_1(40447) <= 3777682;
srom_1(40448) <= 4268091;
srom_1(40449) <= 4777824;
srom_1(40450) <= 5304488;
srom_1(40451) <= 5845615;
srom_1(40452) <= 6398667;
srom_1(40453) <= 6961050;
srom_1(40454) <= 7530128;
srom_1(40455) <= 8103231;
srom_1(40456) <= 8677673;
srom_1(40457) <= 9250759;
srom_1(40458) <= 9819802;
srom_1(40459) <= 10382134;
srom_1(40460) <= 10935117;
srom_1(40461) <= 11476159;
srom_1(40462) <= 12002722;
srom_1(40463) <= 12512338;
srom_1(40464) <= 13002616;
srom_1(40465) <= 13471257;
srom_1(40466) <= 13916064;
srom_1(40467) <= 14334951;
srom_1(40468) <= 14725953;
srom_1(40469) <= 15087238;
srom_1(40470) <= 15417110;
srom_1(40471) <= 15714023;
srom_1(40472) <= 15976585;
srom_1(40473) <= 16203564;
srom_1(40474) <= 16393896;
srom_1(40475) <= 16546688;
srom_1(40476) <= 16661225;
srom_1(40477) <= 16736968;
srom_1(40478) <= 16773563;
srom_1(40479) <= 16770838;
srom_1(40480) <= 16728806;
srom_1(40481) <= 16647664;
srom_1(40482) <= 16527792;
srom_1(40483) <= 16369753;
srom_1(40484) <= 16174287;
srom_1(40485) <= 15942312;
srom_1(40486) <= 15674915;
srom_1(40487) <= 15373350;
srom_1(40488) <= 15039031;
srom_1(40489) <= 14673526;
srom_1(40490) <= 14278548;
srom_1(40491) <= 13855951;
srom_1(40492) <= 13407716;
srom_1(40493) <= 12935944;
srom_1(40494) <= 12442848;
srom_1(40495) <= 11930740;
srom_1(40496) <= 11402022;
srom_1(40497) <= 10859174;
srom_1(40498) <= 10304739;
srom_1(40499) <= 9741320;
srom_1(40500) <= 9171557;
srom_1(40501) <= 8598122;
srom_1(40502) <= 8023706;
srom_1(40503) <= 7451000;
srom_1(40504) <= 6882691;
srom_1(40505) <= 6321444;
srom_1(40506) <= 5769890;
srom_1(40507) <= 5230616;
srom_1(40508) <= 4706152;
srom_1(40509) <= 4198955;
srom_1(40510) <= 3711406;
srom_1(40511) <= 3245789;
srom_1(40512) <= 2804289;
srom_1(40513) <= 2388975;
srom_1(40514) <= 2001796;
srom_1(40515) <= 1644567;
srom_1(40516) <= 1318963;
srom_1(40517) <= 1026511;
srom_1(40518) <= 768582;
srom_1(40519) <= 546387;
srom_1(40520) <= 360966;
srom_1(40521) <= 213189;
srom_1(40522) <= 103750;
srom_1(40523) <= 33161;
srom_1(40524) <= 1754;
srom_1(40525) <= 9676;
srom_1(40526) <= 56890;
srom_1(40527) <= 143173;
srom_1(40528) <= 268123;
srom_1(40529) <= 431152;
srom_1(40530) <= 631496;
srom_1(40531) <= 868216;
srom_1(40532) <= 1140202;
srom_1(40533) <= 1446178;
srom_1(40534) <= 1784710;
srom_1(40535) <= 2154209;
srom_1(40536) <= 2552944;
srom_1(40537) <= 2979044;
srom_1(40538) <= 3430511;
srom_1(40539) <= 3905229;
srom_1(40540) <= 4400971;
srom_1(40541) <= 4915412;
srom_1(40542) <= 5446140;
srom_1(40543) <= 5990666;
srom_1(40544) <= 6546437;
srom_1(40545) <= 7110847;
srom_1(40546) <= 7681249;
srom_1(40547) <= 8254967;
srom_1(40548) <= 8829312;
srom_1(40549) <= 9401591;
srom_1(40550) <= 9969119;
srom_1(40551) <= 10529236;
srom_1(40552) <= 11079315;
srom_1(40553) <= 11616776;
srom_1(40554) <= 12139099;
srom_1(40555) <= 12643835;
srom_1(40556) <= 13128616;
srom_1(40557) <= 13591170;
srom_1(40558) <= 14029327;
srom_1(40559) <= 14441033;
srom_1(40560) <= 14824358;
srom_1(40561) <= 15177502;
srom_1(40562) <= 15498811;
srom_1(40563) <= 15786778;
srom_1(40564) <= 16040053;
srom_1(40565) <= 16257447;
srom_1(40566) <= 16437942;
srom_1(40567) <= 16580690;
srom_1(40568) <= 16685023;
srom_1(40569) <= 16750451;
srom_1(40570) <= 16776668;
srom_1(40571) <= 16763550;
srom_1(40572) <= 16711159;
srom_1(40573) <= 16619741;
srom_1(40574) <= 16489724;
srom_1(40575) <= 16321718;
srom_1(40576) <= 16116511;
srom_1(40577) <= 15875066;
srom_1(40578) <= 15598513;
srom_1(40579) <= 15288152;
srom_1(40580) <= 14945435;
srom_1(40581) <= 14571972;
srom_1(40582) <= 14169512;
srom_1(40583) <= 13739944;
srom_1(40584) <= 13285282;
srom_1(40585) <= 12807657;
srom_1(40586) <= 12309310;
srom_1(40587) <= 11792578;
srom_1(40588) <= 11259883;
srom_1(40589) <= 10713724;
srom_1(40590) <= 10156661;
srom_1(40591) <= 9591308;
srom_1(40592) <= 9020314;
srom_1(40593) <= 8446358;
srom_1(40594) <= 7872132;
srom_1(40595) <= 7300327;
srom_1(40596) <= 6733626;
srom_1(40597) <= 6174685;
srom_1(40598) <= 5626127;
srom_1(40599) <= 5090522;
srom_1(40600) <= 4570383;
srom_1(40601) <= 4068150;
srom_1(40602) <= 3586176;
srom_1(40603) <= 3126723;
srom_1(40604) <= 2691944;
srom_1(40605) <= 2283879;
srom_1(40606) <= 1904441;
srom_1(40607) <= 1555410;
srom_1(40608) <= 1238422;
srom_1(40609) <= 954964;
srom_1(40610) <= 706364;
srom_1(40611) <= 493789;
srom_1(40612) <= 318236;
srom_1(40613) <= 180527;
srom_1(40614) <= 81309;
srom_1(40615) <= 21047;
srom_1(40616) <= 23;
srom_1(40617) <= 18336;
srom_1(40618) <= 75900;
srom_1(40619) <= 172445;
srom_1(40620) <= 307519;
srom_1(40621) <= 480487;
srom_1(40622) <= 690540;
srom_1(40623) <= 936691;
srom_1(40624) <= 1217787;
srom_1(40625) <= 1532509;
srom_1(40626) <= 1879382;
srom_1(40627) <= 2256779;
srom_1(40628) <= 2662931;
srom_1(40629) <= 3095932;
srom_1(40630) <= 3553752;
srom_1(40631) <= 4034244;
srom_1(40632) <= 4535155;
srom_1(40633) <= 5054137;
srom_1(40634) <= 5588755;
srom_1(40635) <= 6136503;
srom_1(40636) <= 6694811;
srom_1(40637) <= 7261062;
srom_1(40638) <= 7832601;
srom_1(40639) <= 8406747;
srom_1(40640) <= 8980808;
srom_1(40641) <= 9552092;
srom_1(40642) <= 10117919;
srom_1(40643) <= 10675638;
srom_1(40644) <= 11222632;
srom_1(40645) <= 11756336;
srom_1(40646) <= 12274248;
srom_1(40647) <= 12773938;
srom_1(40648) <= 13253065;
srom_1(40649) <= 13709380;
srom_1(40650) <= 14140744;
srom_1(40651) <= 14545134;
srom_1(40652) <= 14920655;
srom_1(40653) <= 15265544;
srom_1(40654) <= 15578185;
srom_1(40655) <= 15857112;
srom_1(40656) <= 16101016;
srom_1(40657) <= 16308754;
srom_1(40658) <= 16479352;
srom_1(40659) <= 16612010;
srom_1(40660) <= 16706105;
srom_1(40661) <= 16761196;
srom_1(40662) <= 16777026;
srom_1(40663) <= 16753519;
srom_1(40664) <= 16690787;
srom_1(40665) <= 16589123;
srom_1(40666) <= 16449003;
srom_1(40667) <= 16271086;
srom_1(40668) <= 16056205;
srom_1(40669) <= 15805368;
srom_1(40670) <= 15519751;
srom_1(40671) <= 15200694;
srom_1(40672) <= 14849693;
srom_1(40673) <= 14468393;
srom_1(40674) <= 14058584;
srom_1(40675) <= 13622185;
srom_1(40676) <= 13161245;
srom_1(40677) <= 12677924;
srom_1(40678) <= 12174489;
srom_1(40679) <= 11653301;
srom_1(40680) <= 11116804;
srom_1(40681) <= 10567513;
srom_1(40682) <= 10008004;
srom_1(40683) <= 9440902;
srom_1(40684) <= 8868865;
srom_1(40685) <= 8294575;
srom_1(40686) <= 7720727;
srom_1(40687) <= 7150011;
srom_1(40688) <= 6585103;
srom_1(40689) <= 6028652;
srom_1(40690) <= 5483268;
srom_1(40691) <= 4951508;
srom_1(40692) <= 4435865;
srom_1(40693) <= 3938759;
srom_1(40694) <= 3462519;
srom_1(40695) <= 3009379;
srom_1(40696) <= 2581465;
srom_1(40697) <= 2180782;
srom_1(40698) <= 1809210;
srom_1(40699) <= 1468490;
srom_1(40700) <= 1160222;
srom_1(40701) <= 885850;
srom_1(40702) <= 646661;
srom_1(40703) <= 443776;
srom_1(40704) <= 278148;
srom_1(40705) <= 150553;
srom_1(40706) <= 61588;
srom_1(40707) <= 11672;
srom_1(40708) <= 1038;
srom_1(40709) <= 29736;
srom_1(40710) <= 97632;
srom_1(40711) <= 204407;
srom_1(40712) <= 349560;
srom_1(40713) <= 532412;
srom_1(40714) <= 752104;
srom_1(40715) <= 1007606;
srom_1(40716) <= 1297720;
srom_1(40717) <= 1621085;
srom_1(40718) <= 1976186;
srom_1(40719) <= 2361357;
srom_1(40720) <= 2774792;
srom_1(40721) <= 3214552;
srom_1(40722) <= 3678575;
srom_1(40723) <= 4164684;
srom_1(40724) <= 4670602;
srom_1(40725) <= 5193954;
srom_1(40726) <= 5732287;
srom_1(40727) <= 6283076;
srom_1(40728) <= 6843739;
srom_1(40729) <= 7411647;
srom_1(40730) <= 7984135;
srom_1(40731) <= 8558521;
srom_1(40732) <= 9132109;
srom_1(40733) <= 9702211;
srom_1(40734) <= 10266153;
srom_1(40735) <= 10821291;
srom_1(40736) <= 11365021;
srom_1(40737) <= 11894794;
srom_1(40738) <= 12408124;
srom_1(40739) <= 12902606;
srom_1(40740) <= 13375920;
srom_1(40741) <= 13825847;
srom_1(40742) <= 14250277;
srom_1(40743) <= 14647220;
srom_1(40744) <= 15014814;
srom_1(40745) <= 15351335;
srom_1(40746) <= 15655205;
srom_1(40747) <= 15925000;
srom_1(40748) <= 16159454;
srom_1(40749) <= 16357468;
srom_1(40750) <= 16518114;
srom_1(40751) <= 16640637;
srom_1(40752) <= 16724464;
srom_1(40753) <= 16769201;
srom_1(40754) <= 16774638;
srom_1(40755) <= 16740751;
srom_1(40756) <= 16667697;
srom_1(40757) <= 16555820;
srom_1(40758) <= 16405644;
srom_1(40759) <= 16217873;
srom_1(40760) <= 15993389;
srom_1(40761) <= 15733242;
srom_1(40762) <= 15438655;
srom_1(40763) <= 15111007;
srom_1(40764) <= 14751835;
srom_1(40765) <= 14362825;
srom_1(40766) <= 13945799;
srom_1(40767) <= 13502713;
srom_1(40768) <= 13035646;
srom_1(40769) <= 12546787;
srom_1(40770) <= 12038429;
srom_1(40771) <= 11512956;
srom_1(40772) <= 10972831;
srom_1(40773) <= 10420588;
srom_1(40774) <= 9858817;
srom_1(40775) <= 9290151;
srom_1(40776) <= 8717258;
srom_1(40777) <= 8142823;
srom_1(40778) <= 7569541;
srom_1(40779) <= 7000100;
srom_1(40780) <= 6437170;
srom_1(40781) <= 5883391;
srom_1(40782) <= 5341360;
srom_1(40783) <= 4813618;
srom_1(40784) <= 4302641;
srom_1(40785) <= 3810824;
srom_1(40786) <= 3340474;
srom_1(40787) <= 2893797;
srom_1(40788) <= 2472886;
srom_1(40789) <= 2079717;
srom_1(40790) <= 1716132;
srom_1(40791) <= 1383836;
srom_1(40792) <= 1084388;
srom_1(40793) <= 819193;
srom_1(40794) <= 589492;
srom_1(40795) <= 396365;
srom_1(40796) <= 240716;
srom_1(40797) <= 123275;
srom_1(40798) <= 44593;
srom_1(40799) <= 5039;
srom_1(40800) <= 4799;
srom_1(40801) <= 43873;
srom_1(40802) <= 122078;
srom_1(40803) <= 239048;
srom_1(40804) <= 394234;
srom_1(40805) <= 586908;
srom_1(40806) <= 816168;
srom_1(40807) <= 1080937;
srom_1(40808) <= 1379974;
srom_1(40809) <= 1711877;
srom_1(40810) <= 2075090;
srom_1(40811) <= 2467908;
srom_1(40812) <= 2888491;
srom_1(40813) <= 3334866;
srom_1(40814) <= 3804940;
srom_1(40815) <= 4296508;
srom_1(40816) <= 4807265;
srom_1(40817) <= 5334817;
srom_1(40818) <= 5876688;
srom_1(40819) <= 6430339;
srom_1(40820) <= 6993173;
srom_1(40821) <= 7562551;
srom_1(40822) <= 8135802;
srom_1(40823) <= 8710239;
srom_1(40824) <= 9283167;
srom_1(40825) <= 9851901;
srom_1(40826) <= 10413773;
srom_1(40827) <= 10966148;
srom_1(40828) <= 11506436;
srom_1(40829) <= 12032103;
srom_1(40830) <= 12540685;
srom_1(40831) <= 13029796;
srom_1(40832) <= 13497144;
srom_1(40833) <= 13940535;
srom_1(40834) <= 14357892;
srom_1(40835) <= 14747256;
srom_1(40836) <= 15106803;
srom_1(40837) <= 15434846;
srom_1(40838) <= 15729846;
srom_1(40839) <= 15990421;
srom_1(40840) <= 16215349;
srom_1(40841) <= 16403574;
srom_1(40842) <= 16554214;
srom_1(40843) <= 16666563;
srom_1(40844) <= 16740093;
srom_1(40845) <= 16774461;
srom_1(40846) <= 16769505;
srom_1(40847) <= 16725247;
srom_1(40848) <= 16641896;
srom_1(40849) <= 16519843;
srom_1(40850) <= 16359660;
srom_1(40851) <= 16162097;
srom_1(40852) <= 15928082;
srom_1(40853) <= 15658712;
srom_1(40854) <= 15355250;
srom_1(40855) <= 15019119;
srom_1(40856) <= 14651895;
srom_1(40857) <= 14255300;
srom_1(40858) <= 13831194;
srom_1(40859) <= 13381567;
srom_1(40860) <= 12908525;
srom_1(40861) <= 12414288;
srom_1(40862) <= 11901173;
srom_1(40863) <= 11371587;
srom_1(40864) <= 10828013;
srom_1(40865) <= 10272999;
srom_1(40866) <= 9709148;
srom_1(40867) <= 9139106;
srom_1(40868) <= 8565543;
srom_1(40869) <= 7991151;
srom_1(40870) <= 7418623;
srom_1(40871) <= 6850644;
srom_1(40872) <= 6289876;
srom_1(40873) <= 5738950;
srom_1(40874) <= 5200450;
srom_1(40875) <= 4676900;
srom_1(40876) <= 4170755;
srom_1(40877) <= 3684389;
srom_1(40878) <= 3220083;
srom_1(40879) <= 2780013;
srom_1(40880) <= 2366245;
srom_1(40881) <= 1980717;
srom_1(40882) <= 1625238;
srom_1(40883) <= 1301475;
srom_1(40884) <= 1010946;
srom_1(40885) <= 755013;
srom_1(40886) <= 534877;
srom_1(40887) <= 351570;
srom_1(40888) <= 205951;
srom_1(40889) <= 98703;
srom_1(40890) <= 30330;
srom_1(40891) <= 1151;
srom_1(40892) <= 11304;
srom_1(40893) <= 60741;
srom_1(40894) <= 149231;
srom_1(40895) <= 276357;
srom_1(40896) <= 441525;
srom_1(40897) <= 643959;
srom_1(40898) <= 882711;
srom_1(40899) <= 1156660;
srom_1(40900) <= 1464523;
srom_1(40901) <= 1804854;
srom_1(40902) <= 2176060;
srom_1(40903) <= 2576398;
srom_1(40904) <= 3003991;
srom_1(40905) <= 3456835;
srom_1(40906) <= 3932806;
srom_1(40907) <= 4429671;
srom_1(40908) <= 4945101;
srom_1(40909) <= 5476679;
srom_1(40910) <= 6021912;
srom_1(40911) <= 6578243;
srom_1(40912) <= 7143064;
srom_1(40913) <= 7713726;
srom_1(40914) <= 8287552;
srom_1(40915) <= 8861852;
srom_1(40916) <= 9433933;
srom_1(40917) <= 10001112;
srom_1(40918) <= 10560729;
srom_1(40919) <= 11110160;
srom_1(40920) <= 11646830;
srom_1(40921) <= 12168220;
srom_1(40922) <= 12671886;
srom_1(40923) <= 13155467;
srom_1(40924) <= 13616694;
srom_1(40925) <= 14053405;
srom_1(40926) <= 14463552;
srom_1(40927) <= 14845211;
srom_1(40928) <= 15196593;
srom_1(40929) <= 15516050;
srom_1(40930) <= 15802084;
srom_1(40931) <= 16053353;
srom_1(40932) <= 16268680;
srom_1(40933) <= 16447055;
srom_1(40934) <= 16587641;
srom_1(40935) <= 16689778;
srom_1(40936) <= 16752989;
srom_1(40937) <= 16776976;
srom_1(40938) <= 16761627;
srom_1(40939) <= 16707015;
srom_1(40940) <= 16613394;
srom_1(40941) <= 16481204;
srom_1(40942) <= 16311066;
srom_1(40943) <= 16103776;
srom_1(40944) <= 15860308;
srom_1(40945) <= 15581802;
srom_1(40946) <= 15269564;
srom_1(40947) <= 14925060;
srom_1(40948) <= 14549903;
srom_1(40949) <= 14145855;
srom_1(40950) <= 13714808;
srom_1(40951) <= 13258785;
srom_1(40952) <= 12779925;
srom_1(40953) <= 12280472;
srom_1(40954) <= 11762768;
srom_1(40955) <= 11229242;
srom_1(40956) <= 10682395;
srom_1(40957) <= 10124792;
srom_1(40958) <= 9559047;
srom_1(40959) <= 8987814;
srom_1(40960) <= 8413771;
srom_1(40961) <= 7839610;
srom_1(40962) <= 7268023;
srom_1(40963) <= 6701691;
srom_1(40964) <= 6143270;
srom_1(40965) <= 5595377;
srom_1(40966) <= 5060584;
srom_1(40967) <= 4541396;
srom_1(40968) <= 4040249;
srom_1(40969) <= 3559493;
srom_1(40970) <= 3101383;
srom_1(40971) <= 2668066;
srom_1(40972) <= 2261575;
srom_1(40973) <= 1883815;
srom_1(40974) <= 1536559;
srom_1(40975) <= 1221435;
srom_1(40976) <= 939919;
srom_1(40977) <= 693333;
srom_1(40978) <= 482833;
srom_1(40979) <= 309406;
srom_1(40980) <= 173865;
srom_1(40981) <= 76846;
srom_1(40982) <= 18803;
srom_1(40983) <= 9;
srom_1(40984) <= 20553;
srom_1(40985) <= 80336;
srom_1(40986) <= 179081;
srom_1(40987) <= 316322;
srom_1(40988) <= 491418;
srom_1(40989) <= 703546;
srom_1(40990) <= 951711;
srom_1(40991) <= 1234751;
srom_1(40992) <= 1551338;
srom_1(40993) <= 1899987;
srom_1(40994) <= 2279064;
srom_1(40995) <= 2686790;
srom_1(40996) <= 3121254;
srom_1(40997) <= 3580419;
srom_1(40998) <= 4062130;
srom_1(40999) <= 4564130;
srom_1(41000) <= 5084065;
srom_1(41001) <= 5619495;
srom_1(41002) <= 6167911;
srom_1(41003) <= 6726740;
srom_1(41004) <= 7293363;
srom_1(41005) <= 7865121;
srom_1(41006) <= 8439334;
srom_1(41007) <= 9013310;
srom_1(41008) <= 9584356;
srom_1(41009) <= 10149794;
srom_1(41010) <= 10706974;
srom_1(41011) <= 11253282;
srom_1(41012) <= 11786157;
srom_1(41013) <= 12303099;
srom_1(41014) <= 12801685;
srom_1(41015) <= 13279577;
srom_1(41016) <= 13734533;
srom_1(41017) <= 14164420;
srom_1(41018) <= 14567223;
srom_1(41019) <= 14941052;
srom_1(41020) <= 15284154;
srom_1(41021) <= 15594920;
srom_1(41022) <= 15871894;
srom_1(41023) <= 16113776;
srom_1(41024) <= 16319432;
srom_1(41025) <= 16487898;
srom_1(41026) <= 16618383;
srom_1(41027) <= 16710276;
srom_1(41028) <= 16763146;
srom_1(41029) <= 16776745;
srom_1(41030) <= 16751009;
srom_1(41031) <= 16686058;
srom_1(41032) <= 16582199;
srom_1(41033) <= 16439916;
srom_1(41034) <= 16259878;
srom_1(41035) <= 16042930;
srom_1(41036) <= 15790087;
srom_1(41037) <= 15502536;
srom_1(41038) <= 15181626;
srom_1(41039) <= 14828861;
srom_1(41040) <= 14445895;
srom_1(41041) <= 14034524;
srom_1(41042) <= 13596678;
srom_1(41043) <= 13134410;
srom_1(41044) <= 12649886;
srom_1(41045) <= 12145381;
srom_1(41046) <= 11623258;
srom_1(41047) <= 11085967;
srom_1(41048) <= 10536027;
srom_1(41049) <= 9976017;
srom_1(41050) <= 9408563;
srom_1(41051) <= 8836327;
srom_1(41052) <= 8261990;
srom_1(41053) <= 7688248;
srom_1(41054) <= 7117790;
srom_1(41055) <= 6553291;
srom_1(41056) <= 5997398;
srom_1(41057) <= 5452719;
srom_1(41058) <= 4921807;
srom_1(41059) <= 4407152;
srom_1(41060) <= 3911167;
srom_1(41061) <= 3436179;
srom_1(41062) <= 2984414;
srom_1(41063) <= 2557992;
srom_1(41064) <= 2158911;
srom_1(41065) <= 1789043;
srom_1(41066) <= 1450123;
srom_1(41067) <= 1143740;
srom_1(41068) <= 871331;
srom_1(41069) <= 634173;
srom_1(41070) <= 433378;
srom_1(41071) <= 269887;
srom_1(41072) <= 144468;
srom_1(41073) <= 57709;
srom_1(41074) <= 10016;
srom_1(41075) <= 1614;
srom_1(41076) <= 32540;
srom_1(41077) <= 102652;
srom_1(41078) <= 211619;
srom_1(41079) <= 358930;
srom_1(41080) <= 543896;
srom_1(41081) <= 765648;
srom_1(41082) <= 1023147;
srom_1(41083) <= 1315185;
srom_1(41084) <= 1640392;
srom_1(41085) <= 1997245;
srom_1(41086) <= 2384068;
srom_1(41087) <= 2799049;
srom_1(41088) <= 3240242;
srom_1(41089) <= 3705576;
srom_1(41090) <= 4192871;
srom_1(41091) <= 4699842;
srom_1(41092) <= 5224110;
srom_1(41093) <= 5763218;
srom_1(41094) <= 6314637;
srom_1(41095) <= 6875781;
srom_1(41096) <= 7444020;
srom_1(41097) <= 8016688;
srom_1(41098) <= 8591100;
srom_1(41099) <= 9164563;
srom_1(41100) <= 9734387;
srom_1(41101) <= 10297900;
srom_1(41102) <= 10852460;
srom_1(41103) <= 11395466;
srom_1(41104) <= 11924372;
srom_1(41105) <= 12436697;
srom_1(41106) <= 12930040;
srom_1(41107) <= 13402086;
srom_1(41108) <= 13850622;
srom_1(41109) <= 14273545;
srom_1(41110) <= 14668871;
srom_1(41111) <= 15034747;
srom_1(41112) <= 15369457;
srom_1(41113) <= 15671432;
srom_1(41114) <= 15939255;
srom_1(41115) <= 16171670;
srom_1(41116) <= 16367588;
srom_1(41117) <= 16526089;
srom_1(41118) <= 16646431;
srom_1(41119) <= 16728050;
srom_1(41120) <= 16770561;
srom_1(41121) <= 16773767;
srom_1(41122) <= 16737652;
srom_1(41123) <= 16662386;
srom_1(41124) <= 16548321;
srom_1(41125) <= 16395992;
srom_1(41126) <= 16206114;
srom_1(41127) <= 15979577;
srom_1(41128) <= 15717443;
srom_1(41129) <= 15420942;
srom_1(41130) <= 15091463;
srom_1(41131) <= 14730553;
srom_1(41132) <= 14339903;
srom_1(41133) <= 13921346;
srom_1(41134) <= 13476843;
srom_1(41135) <= 13008480;
srom_1(41136) <= 12518453;
srom_1(41137) <= 12009060;
srom_1(41138) <= 11482689;
srom_1(41139) <= 10941809;
srom_1(41140) <= 10388956;
srom_1(41141) <= 9826722;
srom_1(41142) <= 9257745;
srom_1(41143) <= 8684693;
srom_1(41144) <= 8110251;
srom_1(41145) <= 7537115;
srom_1(41146) <= 6967972;
srom_1(41147) <= 6405491;
srom_1(41148) <= 5852309;
srom_1(41149) <= 5311021;
srom_1(41150) <= 4784165;
srom_1(41151) <= 4274211;
srom_1(41152) <= 3783551;
srom_1(41153) <= 3314486;
srom_1(41154) <= 2869215;
srom_1(41155) <= 2449826;
srom_1(41156) <= 2058287;
srom_1(41157) <= 1696432;
srom_1(41158) <= 1365959;
srom_1(41159) <= 1068418;
srom_1(41160) <= 805204;
srom_1(41161) <= 577551;
srom_1(41162) <= 386526;
srom_1(41163) <= 233027;
srom_1(41164) <= 117771;
srom_1(41165) <= 41300;
srom_1(41166) <= 3973;
srom_1(41167) <= 5964;
srom_1(41168) <= 47264;
srom_1(41169) <= 127680;
srom_1(41170) <= 246834;
srom_1(41171) <= 404167;
srom_1(41172) <= 598942;
srom_1(41173) <= 830246;
srom_1(41174) <= 1096993;
srom_1(41175) <= 1397934;
srom_1(41176) <= 1731656;
srom_1(41177) <= 2096594;
srom_1(41178) <= 2491038;
srom_1(41179) <= 2913138;
srom_1(41180) <= 3360914;
srom_1(41181) <= 3832267;
srom_1(41182) <= 4324986;
srom_1(41183) <= 4836761;
srom_1(41184) <= 5365191;
srom_1(41185) <= 5907800;
srom_1(41186) <= 6462041;
srom_1(41187) <= 7025317;
srom_1(41188) <= 7594986;
srom_1(41189) <= 8168377;
srom_1(41190) <= 8742800;
srom_1(41191) <= 9315563;
srom_1(41192) <= 9883978;
srom_1(41193) <= 10445381;
srom_1(41194) <= 10997140;
srom_1(41195) <= 11536665;
srom_1(41196) <= 12061429;
srom_1(41197) <= 12568970;
srom_1(41198) <= 13056907;
srom_1(41199) <= 13522953;
srom_1(41200) <= 13964922;
srom_1(41201) <= 14380743;
srom_1(41202) <= 14768463;
srom_1(41203) <= 15126267;
srom_1(41204) <= 15452475;
srom_1(41205) <= 15745559;
srom_1(41206) <= 16004143;
srom_1(41207) <= 16227015;
srom_1(41208) <= 16413131;
srom_1(41209) <= 16561616;
srom_1(41210) <= 16671776;
srom_1(41211) <= 16743093;
srom_1(41212) <= 16775233;
srom_1(41213) <= 16768045;
srom_1(41214) <= 16721563;
srom_1(41215) <= 16636005;
srom_1(41216) <= 16511772;
srom_1(41217) <= 16349446;
srom_1(41218) <= 16149790;
srom_1(41219) <= 15913739;
srom_1(41220) <= 15642399;
srom_1(41221) <= 15337045;
srom_1(41222) <= 14999106;
srom_1(41223) <= 14630169;
srom_1(41224) <= 14231963;
srom_1(41225) <= 13806356;
srom_1(41226) <= 13355342;
srom_1(41227) <= 12881038;
srom_1(41228) <= 12385668;
srom_1(41229) <= 11871554;
srom_1(41230) <= 11341107;
srom_1(41231) <= 10796815;
srom_1(41232) <= 10241230;
srom_1(41233) <= 9676957;
srom_1(41234) <= 9106643;
srom_1(41235) <= 8532961;
srom_1(41236) <= 7958603;
srom_1(41237) <= 7386261;
srom_1(41238) <= 6818620;
srom_1(41239) <= 6258341;
srom_1(41240) <= 5708051;
srom_1(41241) <= 5170331;
srom_1(41242) <= 4647703;
srom_1(41243) <= 4142618;
srom_1(41244) <= 3657443;
srom_1(41245) <= 3194454;
srom_1(41246) <= 2755823;
srom_1(41247) <= 2343605;
srom_1(41248) <= 1959735;
srom_1(41249) <= 1606012;
srom_1(41250) <= 1284094;
srom_1(41251) <= 995492;
srom_1(41252) <= 741559;
srom_1(41253) <= 523486;
srom_1(41254) <= 342295;
srom_1(41255) <= 198836;
srom_1(41256) <= 93781;
srom_1(41257) <= 27624;
srom_1(41258) <= 674;
srom_1(41259) <= 13059;
srom_1(41260) <= 64719;
srom_1(41261) <= 155412;
srom_1(41262) <= 284714;
srom_1(41263) <= 452018;
srom_1(41264) <= 656539;
srom_1(41265) <= 897319;
srom_1(41266) <= 1173227;
srom_1(41267) <= 1482971;
srom_1(41268) <= 1825098;
srom_1(41269) <= 2198004;
srom_1(41270) <= 2599939;
srom_1(41271) <= 3029020;
srom_1(41272) <= 3483233;
srom_1(41273) <= 3960450;
srom_1(41274) <= 4458431;
srom_1(41275) <= 4974843;
srom_1(41276) <= 5507263;
srom_1(41277) <= 6053194;
srom_1(41278) <= 6610077;
srom_1(41279) <= 7175300;
srom_1(41280) <= 7746213;
srom_1(41281) <= 8320138;
srom_1(41282) <= 8894384;
srom_1(41283) <= 9466258;
srom_1(41284) <= 10033079;
srom_1(41285) <= 10592189;
srom_1(41286) <= 11140965;
srom_1(41287) <= 11676834;
srom_1(41288) <= 12197284;
srom_1(41289) <= 12699873;
srom_1(41290) <= 13182246;
srom_1(41291) <= 13642139;
srom_1(41292) <= 14077397;
srom_1(41293) <= 14485978;
srom_1(41294) <= 14865967;
srom_1(41295) <= 15215581;
srom_1(41296) <= 15533181;
srom_1(41297) <= 15817277;
srom_1(41298) <= 16066538;
srom_1(41299) <= 16279795;
srom_1(41300) <= 16456047;
srom_1(41301) <= 16594468;
srom_1(41302) <= 16694408;
srom_1(41303) <= 16755401;
srom_1(41304) <= 16777158;
srom_1(41305) <= 16759579;
srom_1(41306) <= 16702745;
srom_1(41307) <= 16606923;
srom_1(41308) <= 16472563;
srom_1(41309) <= 16300294;
srom_1(41310) <= 16090925;
srom_1(41311) <= 15845437;
srom_1(41312) <= 15564981;
srom_1(41313) <= 15250873;
srom_1(41314) <= 14904585;
srom_1(41315) <= 14527742;
srom_1(41316) <= 14122110;
srom_1(41317) <= 13689592;
srom_1(41318) <= 13232215;
srom_1(41319) <= 12752126;
srom_1(41320) <= 12251574;
srom_1(41321) <= 11732907;
srom_1(41322) <= 11198558;
srom_1(41323) <= 10651032;
srom_1(41324) <= 10092897;
srom_1(41325) <= 9526770;
srom_1(41326) <= 8955305;
srom_1(41327) <= 8381183;
srom_1(41328) <= 7807096;
srom_1(41329) <= 7235736;
srom_1(41330) <= 6669782;
srom_1(41331) <= 6111888;
srom_1(41332) <= 5564670;
srom_1(41333) <= 5030695;
srom_1(41334) <= 4512466;
srom_1(41335) <= 4012414;
srom_1(41336) <= 3532884;
srom_1(41337) <= 3076123;
srom_1(41338) <= 2644274;
srom_1(41339) <= 2239363;
srom_1(41340) <= 1863288;
srom_1(41341) <= 1517812;
srom_1(41342) <= 1204555;
srom_1(41343) <= 924987;
srom_1(41344) <= 680419;
srom_1(41345) <= 471996;
srom_1(41346) <= 300698;
srom_1(41347) <= 167327;
srom_1(41348) <= 72507;
srom_1(41349) <= 16685;
srom_1(41350) <= 122;
srom_1(41351) <= 22895;
srom_1(41352) <= 84898;
srom_1(41353) <= 185840;
srom_1(41354) <= 325248;
srom_1(41355) <= 502467;
srom_1(41356) <= 716667;
srom_1(41357) <= 966844;
srom_1(41358) <= 1251824;
srom_1(41359) <= 1570270;
srom_1(41360) <= 1920690;
srom_1(41361) <= 2301441;
srom_1(41362) <= 2710736;
srom_1(41363) <= 3146656;
srom_1(41364) <= 3607158;
srom_1(41365) <= 4090082;
srom_1(41366) <= 4593163;
srom_1(41367) <= 5114042;
srom_1(41368) <= 5650277;
srom_1(41369) <= 6199353;
srom_1(41370) <= 6758695;
srom_1(41371) <= 7325680;
srom_1(41372) <= 7897649;
srom_1(41373) <= 8471921;
srom_1(41374) <= 9045802;
srom_1(41375) <= 9616602;
srom_1(41376) <= 10181642;
srom_1(41377) <= 10738275;
srom_1(41378) <= 11283889;
srom_1(41379) <= 11815927;
srom_1(41380) <= 12331892;
srom_1(41381) <= 12829366;
srom_1(41382) <= 13306016;
srom_1(41383) <= 13759606;
srom_1(41384) <= 14188010;
srom_1(41385) <= 14589218;
srom_1(41386) <= 14961350;
srom_1(41387) <= 15302660;
srom_1(41388) <= 15611547;
srom_1(41389) <= 15886564;
srom_1(41390) <= 16126420;
srom_1(41391) <= 16329990;
srom_1(41392) <= 16496321;
srom_1(41393) <= 16624632;
srom_1(41394) <= 16714322;
srom_1(41395) <= 16764969;
srom_1(41396) <= 16776337;
srom_1(41397) <= 16748372;
srom_1(41398) <= 16681205;
srom_1(41399) <= 16575151;
srom_1(41400) <= 16430708;
srom_1(41401) <= 16248552;
srom_1(41402) <= 16029538;
srom_1(41403) <= 15774694;
srom_1(41404) <= 15485214;
srom_1(41405) <= 15162455;
srom_1(41406) <= 14807931;
srom_1(41407) <= 14423305;
srom_1(41408) <= 14010380;
srom_1(41409) <= 13571092;
srom_1(41410) <= 13107503;
srom_1(41411) <= 12621784;
srom_1(41412) <= 12116215;
srom_1(41413) <= 11593166;
srom_1(41414) <= 11055090;
srom_1(41415) <= 10504509;
srom_1(41416) <= 9944006;
srom_1(41417) <= 9376210;
srom_1(41418) <= 8803782;
srom_1(41419) <= 8229407;
srom_1(41420) <= 7655779;
srom_1(41421) <= 7085588;
srom_1(41422) <= 6521506;
srom_1(41423) <= 5966180;
srom_1(41424) <= 5422214;
srom_1(41425) <= 4892158;
srom_1(41426) <= 4378499;
srom_1(41427) <= 3883644;
srom_1(41428) <= 3409914;
srom_1(41429) <= 2959531;
srom_1(41430) <= 2534607;
srom_1(41431) <= 2137134;
srom_1(41432) <= 1768977;
srom_1(41433) <= 1431861;
srom_1(41434) <= 1127368;
srom_1(41435) <= 856925;
srom_1(41436) <= 621801;
srom_1(41437) <= 423099;
srom_1(41438) <= 261749;
srom_1(41439) <= 138509;
srom_1(41440) <= 53956;
srom_1(41441) <= 8488;
srom_1(41442) <= 2316;
srom_1(41443) <= 35471;
srom_1(41444) <= 107797;
srom_1(41445) <= 218954;
srom_1(41446) <= 368421;
srom_1(41447) <= 555498;
srom_1(41448) <= 779307;
srom_1(41449) <= 1038799;
srom_1(41450) <= 1332756;
srom_1(41451) <= 1659801;
srom_1(41452) <= 2018399;
srom_1(41453) <= 2406870;
srom_1(41454) <= 2823391;
srom_1(41455) <= 3266009;
srom_1(41456) <= 3732649;
srom_1(41457) <= 4221122;
srom_1(41458) <= 4729138;
srom_1(41459) <= 5254314;
srom_1(41460) <= 5794188;
srom_1(41461) <= 6346228;
srom_1(41462) <= 6907846;
srom_1(41463) <= 7476408;
srom_1(41464) <= 8049247;
srom_1(41465) <= 8623677;
srom_1(41466) <= 9197005;
srom_1(41467) <= 9766543;
srom_1(41468) <= 10329618;
srom_1(41469) <= 10883592;
srom_1(41470) <= 11425866;
srom_1(41471) <= 11953897;
srom_1(41472) <= 12465209;
srom_1(41473) <= 12957404;
srom_1(41474) <= 13428175;
srom_1(41475) <= 13875314;
srom_1(41476) <= 14296723;
srom_1(41477) <= 14690428;
srom_1(41478) <= 15054581;
srom_1(41479) <= 15387475;
srom_1(41480) <= 15687549;
srom_1(41481) <= 15953395;
srom_1(41482) <= 16183768;
srom_1(41483) <= 16377586;
srom_1(41484) <= 16533942;
srom_1(41485) <= 16652101;
srom_1(41486) <= 16731510;
srom_1(41487) <= 16771796;
srom_1(41488) <= 16772770;
srom_1(41489) <= 16734428;
srom_1(41490) <= 16656950;
srom_1(41491) <= 16540699;
srom_1(41492) <= 16386219;
srom_1(41493) <= 16194236;
srom_1(41494) <= 15965650;
srom_1(41495) <= 15701533;
srom_1(41496) <= 15403122;
srom_1(41497) <= 15071819;
srom_1(41498) <= 14709175;
srom_1(41499) <= 14316892;
srom_1(41500) <= 13896809;
srom_1(41501) <= 13450896;
srom_1(41502) <= 12981245;
srom_1(41503) <= 12490057;
srom_1(41504) <= 11979636;
srom_1(41505) <= 11452376;
srom_1(41506) <= 10910748;
srom_1(41507) <= 10357293;
srom_1(41508) <= 9794606;
srom_1(41509) <= 9225326;
srom_1(41510) <= 8652123;
srom_1(41511) <= 8077684;
srom_1(41512) <= 7504702;
srom_1(41513) <= 6935866;
srom_1(41514) <= 6373842;
srom_1(41515) <= 5821266;
srom_1(41516) <= 5280729;
srom_1(41517) <= 4754766;
srom_1(41518) <= 4245844;
srom_1(41519) <= 3756348;
srom_1(41520) <= 3288574;
srom_1(41521) <= 2844716;
srom_1(41522) <= 2426856;
srom_1(41523) <= 2036952;
srom_1(41524) <= 1676833;
srom_1(41525) <= 1348188;
srom_1(41526) <= 1052558;
srom_1(41527) <= 791330;
srom_1(41528) <= 565727;
srom_1(41529) <= 376809;
srom_1(41530) <= 225460;
srom_1(41531) <= 112392;
srom_1(41532) <= 38134;
srom_1(41533) <= 3033;
srom_1(41534) <= 7256;
srom_1(41535) <= 50782;
srom_1(41536) <= 133406;
srom_1(41537) <= 254742;
srom_1(41538) <= 414221;
srom_1(41539) <= 611094;
srom_1(41540) <= 844438;
srom_1(41541) <= 1113160;
srom_1(41542) <= 1415999;
srom_1(41543) <= 1751535;
srom_1(41544) <= 2118194;
srom_1(41545) <= 2514258;
srom_1(41546) <= 2937868;
srom_1(41547) <= 3387039;
srom_1(41548) <= 3859663;
srom_1(41549) <= 4353526;
srom_1(41550) <= 4866310;
srom_1(41551) <= 5395612;
srom_1(41552) <= 5938949;
srom_1(41553) <= 6493773;
srom_1(41554) <= 7057482;
srom_1(41555) <= 7627434;
srom_1(41556) <= 8200955;
srom_1(41557) <= 8775356;
srom_1(41558) <= 9347944;
srom_1(41559) <= 9916033;
srom_1(41560) <= 10476959;
srom_1(41561) <= 11028092;
srom_1(41562) <= 11566848;
srom_1(41563) <= 12090700;
srom_1(41564) <= 12597191;
srom_1(41565) <= 13083947;
srom_1(41566) <= 13548685;
srom_1(41567) <= 13989226;
srom_1(41568) <= 14403503;
srom_1(41569) <= 14789574;
srom_1(41570) <= 15145629;
srom_1(41571) <= 15469998;
srom_1(41572) <= 15761160;
srom_1(41573) <= 16017750;
srom_1(41574) <= 16238564;
srom_1(41575) <= 16422567;
srom_1(41576) <= 16568895;
srom_1(41577) <= 16676864;
srom_1(41578) <= 16745966;
srom_1(41579) <= 16775877;
srom_1(41580) <= 16766458;
srom_1(41581) <= 16717752;
srom_1(41582) <= 16629988;
srom_1(41583) <= 16503577;
srom_1(41584) <= 16339113;
srom_1(41585) <= 16137365;
srom_1(41586) <= 15899281;
srom_1(41587) <= 15625977;
srom_1(41588) <= 15318735;
srom_1(41589) <= 14978994;
srom_1(41590) <= 14608350;
srom_1(41591) <= 14208538;
srom_1(41592) <= 13781435;
srom_1(41593) <= 13329043;
srom_1(41594) <= 12853484;
srom_1(41595) <= 12356987;
srom_1(41596) <= 11841881;
srom_1(41597) <= 11310582;
srom_1(41598) <= 10765581;
srom_1(41599) <= 10209433;
srom_1(41600) <= 9644746;
srom_1(41601) <= 9074169;
srom_1(41602) <= 8500377;
srom_1(41603) <= 7926062;
srom_1(41604) <= 7353915;
srom_1(41605) <= 6786620;
srom_1(41606) <= 6226837;
srom_1(41607) <= 5677192;
srom_1(41608) <= 5140262;
srom_1(41609) <= 4618564;
srom_1(41610) <= 4114545;
srom_1(41611) <= 3630568;
srom_1(41612) <= 3168904;
srom_1(41613) <= 2731717;
srom_1(41614) <= 2321057;
srom_1(41615) <= 1938849;
srom_1(41616) <= 1586887;
srom_1(41617) <= 1266820;
srom_1(41618) <= 980150;
srom_1(41619) <= 728221;
srom_1(41620) <= 512214;
srom_1(41621) <= 333142;
srom_1(41622) <= 191845;
srom_1(41623) <= 88985;
srom_1(41624) <= 25045;
srom_1(41625) <= 324;
srom_1(41626) <= 14940;
srom_1(41627) <= 68822;
srom_1(41628) <= 161718;
srom_1(41629) <= 293193;
srom_1(41630) <= 462631;
srom_1(41631) <= 669236;
srom_1(41632) <= 912039;
srom_1(41633) <= 1189903;
srom_1(41634) <= 1501525;
srom_1(41635) <= 1845442;
srom_1(41636) <= 2220042;
srom_1(41637) <= 2623569;
srom_1(41638) <= 3054129;
srom_1(41639) <= 3509706;
srom_1(41640) <= 3988161;
srom_1(41641) <= 4487251;
srom_1(41642) <= 5004636;
srom_1(41643) <= 5537889;
srom_1(41644) <= 6084511;
srom_1(41645) <= 6641937;
srom_1(41646) <= 7207554;
srom_1(41647) <= 7778710;
srom_1(41648) <= 8352725;
srom_1(41649) <= 8926909;
srom_1(41650) <= 9498568;
srom_1(41651) <= 10065022;
srom_1(41652) <= 10623616;
srom_1(41653) <= 11171728;
srom_1(41654) <= 11706789;
srom_1(41655) <= 12226290;
srom_1(41656) <= 12727795;
srom_1(41657) <= 13208953;
srom_1(41658) <= 13667505;
srom_1(41659) <= 14101304;
srom_1(41660) <= 14508313;
srom_1(41661) <= 14886625;
srom_1(41662) <= 15234466;
srom_1(41663) <= 15550204;
srom_1(41664) <= 15832359;
srom_1(41665) <= 16079607;
srom_1(41666) <= 16290790;
srom_1(41667) <= 16464917;
srom_1(41668) <= 16601171;
srom_1(41669) <= 16698913;
srom_1(41670) <= 16757686;
srom_1(41671) <= 16777213;
srom_1(41672) <= 16757403;
srom_1(41673) <= 16698349;
srom_1(41674) <= 16600328;
srom_1(41675) <= 16463799;
srom_1(41676) <= 16289403;
srom_1(41677) <= 16077957;
srom_1(41678) <= 15830454;
srom_1(41679) <= 15548053;
srom_1(41680) <= 15232078;
srom_1(41681) <= 14884013;
srom_1(41682) <= 14505488;
srom_1(41683) <= 14098279;
srom_1(41684) <= 13664295;
srom_1(41685) <= 13205572;
srom_1(41686) <= 12724261;
srom_1(41687) <= 12222618;
srom_1(41688) <= 11702996;
srom_1(41689) <= 11167832;
srom_1(41690) <= 10619635;
srom_1(41691) <= 10060976;
srom_1(41692) <= 9494475;
srom_1(41693) <= 8922788;
srom_1(41694) <= 8348596;
srom_1(41695) <= 7774591;
srom_1(41696) <= 7203466;
srom_1(41697) <= 6637898;
srom_1(41698) <= 6080541;
srom_1(41699) <= 5534006;
srom_1(41700) <= 5000858;
srom_1(41701) <= 4483595;
srom_1(41702) <= 3984645;
srom_1(41703) <= 3506347;
srom_1(41704) <= 3050943;
srom_1(41705) <= 2620569;
srom_1(41706) <= 2217244;
srom_1(41707) <= 1842858;
srom_1(41708) <= 1499168;
srom_1(41709) <= 1187784;
srom_1(41710) <= 910168;
srom_1(41711) <= 667620;
srom_1(41712) <= 461279;
srom_1(41713) <= 292112;
srom_1(41714) <= 160912;
srom_1(41715) <= 68295;
srom_1(41716) <= 14694;
srom_1(41717) <= 362;
srom_1(41718) <= 25365;
srom_1(41719) <= 89586;
srom_1(41720) <= 192724;
srom_1(41721) <= 334295;
srom_1(41722) <= 513636;
srom_1(41723) <= 729905;
srom_1(41724) <= 982088;
srom_1(41725) <= 1269003;
srom_1(41726) <= 1589305;
srom_1(41727) <= 1941491;
srom_1(41728) <= 2323909;
srom_1(41729) <= 2734767;
srom_1(41730) <= 3172138;
srom_1(41731) <= 3633970;
srom_1(41732) <= 4118099;
srom_1(41733) <= 4622253;
srom_1(41734) <= 5144069;
srom_1(41735) <= 5681100;
srom_1(41736) <= 6230828;
srom_1(41737) <= 6790674;
srom_1(41738) <= 7358013;
srom_1(41739) <= 7930185;
srom_1(41740) <= 8504507;
srom_1(41741) <= 9078285;
srom_1(41742) <= 9648829;
srom_1(41743) <= 10213463;
srom_1(41744) <= 10769541;
srom_1(41745) <= 11314453;
srom_1(41746) <= 11845644;
srom_1(41747) <= 12360625;
srom_1(41748) <= 12856979;
srom_1(41749) <= 13332380;
srom_1(41750) <= 13784598;
srom_1(41751) <= 14211511;
srom_1(41752) <= 14611120;
srom_1(41753) <= 14981549;
srom_1(41754) <= 15321061;
srom_1(41755) <= 15628064;
srom_1(41756) <= 15901120;
srom_1(41757) <= 16138946;
srom_1(41758) <= 16340429;
srom_1(41759) <= 16504623;
srom_1(41760) <= 16630757;
srom_1(41761) <= 16718242;
srom_1(41762) <= 16766666;
srom_1(41763) <= 16775803;
srom_1(41764) <= 16745609;
srom_1(41765) <= 16676226;
srom_1(41766) <= 16567980;
srom_1(41767) <= 16421378;
srom_1(41768) <= 16237107;
srom_1(41769) <= 16016032;
srom_1(41770) <= 15759190;
srom_1(41771) <= 15467784;
srom_1(41772) <= 15143181;
srom_1(41773) <= 14786904;
srom_1(41774) <= 14400624;
srom_1(41775) <= 13986150;
srom_1(41776) <= 13545429;
srom_1(41777) <= 13080524;
srom_1(41778) <= 12593618;
srom_1(41779) <= 12086993;
srom_1(41780) <= 11563026;
srom_1(41781) <= 11024172;
srom_1(41782) <= 10472959;
srom_1(41783) <= 9911972;
srom_1(41784) <= 9343841;
srom_1(41785) <= 8771231;
srom_1(41786) <= 8196827;
srom_1(41787) <= 7623322;
srom_1(41788) <= 7053405;
srom_1(41789) <= 6489750;
srom_1(41790) <= 5934999;
srom_1(41791) <= 5391754;
srom_1(41792) <= 4862563;
srom_1(41793) <= 4349906;
srom_1(41794) <= 3856188;
srom_1(41795) <= 3383724;
srom_1(41796) <= 2934730;
srom_1(41797) <= 2511310;
srom_1(41798) <= 2115452;
srom_1(41799) <= 1749010;
srom_1(41800) <= 1413704;
srom_1(41801) <= 1111105;
srom_1(41802) <= 842634;
srom_1(41803) <= 609547;
srom_1(41804) <= 412940;
srom_1(41805) <= 253733;
srom_1(41806) <= 132674;
srom_1(41807) <= 50329;
srom_1(41808) <= 7085;
srom_1(41809) <= 3145;
srom_1(41810) <= 38528;
srom_1(41811) <= 113067;
srom_1(41812) <= 226412;
srom_1(41813) <= 378033;
srom_1(41814) <= 567219;
srom_1(41815) <= 793081;
srom_1(41816) <= 1054562;
srom_1(41817) <= 1350434;
srom_1(41818) <= 1679311;
srom_1(41819) <= 2039650;
srom_1(41820) <= 2429762;
srom_1(41821) <= 2847816;
srom_1(41822) <= 3291853;
srom_1(41823) <= 3759791;
srom_1(41824) <= 4249435;
srom_1(41825) <= 4758489;
srom_1(41826) <= 5284565;
srom_1(41827) <= 5825198;
srom_1(41828) <= 6377851;
srom_1(41829) <= 6939933;
srom_1(41830) <= 7508809;
srom_1(41831) <= 8081810;
srom_1(41832) <= 8656250;
srom_1(41833) <= 9229435;
srom_1(41834) <= 9798677;
srom_1(41835) <= 10361307;
srom_1(41836) <= 10914686;
srom_1(41837) <= 11456219;
srom_1(41838) <= 11983368;
srom_1(41839) <= 12493659;
srom_1(41840) <= 12984700;
srom_1(41841) <= 13454189;
srom_1(41842) <= 13899923;
srom_1(41843) <= 14319813;
srom_1(41844) <= 14711889;
srom_1(41845) <= 15074314;
srom_1(41846) <= 15405386;
srom_1(41847) <= 15703555;
srom_1(41848) <= 15967421;
srom_1(41849) <= 16195748;
srom_1(41850) <= 16387464;
srom_1(41851) <= 16541671;
srom_1(41852) <= 16657646;
srom_1(41853) <= 16734844;
srom_1(41854) <= 16772903;
srom_1(41855) <= 16771646;
srom_1(41856) <= 16731078;
srom_1(41857) <= 16651389;
srom_1(41858) <= 16532953;
srom_1(41859) <= 16376326;
srom_1(41860) <= 16182241;
srom_1(41861) <= 15951609;
srom_1(41862) <= 15685512;
srom_1(41863) <= 15385197;
srom_1(41864) <= 15052073;
srom_1(41865) <= 14687701;
srom_1(41866) <= 14293791;
srom_1(41867) <= 13872189;
srom_1(41868) <= 13424873;
srom_1(41869) <= 12953940;
srom_1(41870) <= 12461599;
srom_1(41871) <= 11950158;
srom_1(41872) <= 11422016;
srom_1(41873) <= 10879649;
srom_1(41874) <= 10325601;
srom_1(41875) <= 9762469;
srom_1(41876) <= 9192895;
srom_1(41877) <= 8619549;
srom_1(41878) <= 8045121;
srom_1(41879) <= 7472303;
srom_1(41880) <= 6903782;
srom_1(41881) <= 6342223;
srom_1(41882) <= 5790261;
srom_1(41883) <= 5250484;
srom_1(41884) <= 4725422;
srom_1(41885) <= 4217538;
srom_1(41886) <= 3729214;
srom_1(41887) <= 3262739;
srom_1(41888) <= 2820302;
srom_1(41889) <= 2403975;
srom_1(41890) <= 2015713;
srom_1(41891) <= 1657336;
srom_1(41892) <= 1330524;
srom_1(41893) <= 1036809;
srom_1(41894) <= 777570;
srom_1(41895) <= 554021;
srom_1(41896) <= 367212;
srom_1(41897) <= 218018;
srom_1(41898) <= 107138;
srom_1(41899) <= 35093;
srom_1(41900) <= 2220;
srom_1(41901) <= 8674;
srom_1(41902) <= 54425;
srom_1(41903) <= 139257;
srom_1(41904) <= 262773;
srom_1(41905) <= 424395;
srom_1(41906) <= 623363;
srom_1(41907) <= 858745;
srom_1(41908) <= 1129437;
srom_1(41909) <= 1434170;
srom_1(41910) <= 1771514;
srom_1(41911) <= 2139889;
srom_1(41912) <= 2537565;
srom_1(41913) <= 2962680;
srom_1(41914) <= 3413238;
srom_1(41915) <= 3887128;
srom_1(41916) <= 4382126;
srom_1(41917) <= 4895913;
srom_1(41918) <= 5426077;
srom_1(41919) <= 5970134;
srom_1(41920) <= 6525532;
srom_1(41921) <= 7089667;
srom_1(41922) <= 7659893;
srom_1(41923) <= 8233536;
srom_1(41924) <= 8807906;
srom_1(41925) <= 9380310;
srom_1(41926) <= 9948064;
srom_1(41927) <= 10508505;
srom_1(41928) <= 11059005;
srom_1(41929) <= 11596982;
srom_1(41930) <= 12119914;
srom_1(41931) <= 12625349;
srom_1(41932) <= 13110916;
srom_1(41933) <= 13574339;
srom_1(41934) <= 14013444;
srom_1(41935) <= 14426172;
srom_1(41936) <= 14810589;
srom_1(41937) <= 15164890;
srom_1(41938) <= 15487415;
srom_1(41939) <= 15776651;
srom_1(41940) <= 16031242;
srom_1(41941) <= 16249994;
srom_1(41942) <= 16431881;
srom_1(41943) <= 16576051;
srom_1(41944) <= 16681827;
srom_1(41945) <= 16748713;
srom_1(41946) <= 16776396;
srom_1(41947) <= 16764745;
srom_1(41948) <= 16713816;
srom_1(41949) <= 16623847;
srom_1(41950) <= 16495261;
srom_1(41951) <= 16328659;
srom_1(41952) <= 16124824;
srom_1(41953) <= 15884711;
srom_1(41954) <= 15609446;
srom_1(41955) <= 15300320;
srom_1(41956) <= 14958783;
srom_1(41957) <= 14586436;
srom_1(41958) <= 14185025;
srom_1(41959) <= 13756433;
srom_1(41960) <= 13302669;
srom_1(41961) <= 12825862;
srom_1(41962) <= 12328247;
srom_1(41963) <= 11812157;
srom_1(41964) <= 11280013;
srom_1(41965) <= 10734310;
srom_1(41966) <= 10177608;
srom_1(41967) <= 9612516;
srom_1(41968) <= 9041685;
srom_1(41969) <= 8467792;
srom_1(41970) <= 7893527;
srom_1(41971) <= 7321584;
srom_1(41972) <= 6754644;
srom_1(41973) <= 6195367;
srom_1(41974) <= 5646374;
srom_1(41975) <= 5110241;
srom_1(41976) <= 4589481;
srom_1(41977) <= 4086536;
srom_1(41978) <= 3603766;
srom_1(41979) <= 3143433;
srom_1(41980) <= 2707697;
srom_1(41981) <= 2298600;
srom_1(41982) <= 1918061;
srom_1(41983) <= 1567865;
srom_1(41984) <= 1249654;
srom_1(41985) <= 964920;
srom_1(41986) <= 714998;
srom_1(41987) <= 501060;
srom_1(41988) <= 324110;
srom_1(41989) <= 184977;
srom_1(41990) <= 84313;
srom_1(41991) <= 22592;
srom_1(41992) <= 101;
srom_1(41993) <= 16947;
srom_1(41994) <= 73050;
srom_1(41995) <= 168148;
srom_1(41996) <= 301795;
srom_1(41997) <= 473363;
srom_1(41998) <= 682049;
srom_1(41999) <= 926873;
srom_1(42000) <= 1206688;
srom_1(42001) <= 1520182;
srom_1(42002) <= 1865883;
srom_1(42003) <= 2242173;
srom_1(42004) <= 2647285;
srom_1(42005) <= 3079320;
srom_1(42006) <= 3536252;
srom_1(42007) <= 4015938;
srom_1(42008) <= 4516129;
srom_1(42009) <= 5034480;
srom_1(42010) <= 5568559;
srom_1(42011) <= 6115863;
srom_1(42012) <= 6673824;
srom_1(42013) <= 7239826;
srom_1(42014) <= 7811216;
srom_1(42015) <= 8385313;
srom_1(42016) <= 8959425;
srom_1(42017) <= 9530861;
srom_1(42018) <= 10096940;
srom_1(42019) <= 10655008;
srom_1(42020) <= 11202449;
srom_1(42021) <= 11736694;
srom_1(42022) <= 12255239;
srom_1(42023) <= 12755652;
srom_1(42024) <= 13235586;
srom_1(42025) <= 13692792;
srom_1(42026) <= 14125124;
srom_1(42027) <= 14530555;
srom_1(42028) <= 14907185;
srom_1(42029) <= 15253247;
srom_1(42030) <= 15567119;
srom_1(42031) <= 15847328;
srom_1(42032) <= 16092560;
srom_1(42033) <= 16301666;
srom_1(42034) <= 16473665;
srom_1(42035) <= 16607750;
srom_1(42036) <= 16703293;
srom_1(42037) <= 16759845;
srom_1(42038) <= 16777142;
srom_1(42039) <= 16755102;
srom_1(42040) <= 16693829;
srom_1(42041) <= 16593609;
srom_1(42042) <= 16454914;
srom_1(42043) <= 16278393;
srom_1(42044) <= 16064874;
srom_1(42045) <= 15815358;
srom_1(42046) <= 15531016;
srom_1(42047) <= 15213180;
srom_1(42048) <= 14863342;
srom_1(42049) <= 14483142;
srom_1(42050) <= 14074362;
srom_1(42051) <= 13638919;
srom_1(42052) <= 13178856;
srom_1(42053) <= 12696330;
srom_1(42054) <= 12193604;
srom_1(42055) <= 11673035;
srom_1(42056) <= 11137064;
srom_1(42057) <= 10588204;
srom_1(42058) <= 10029030;
srom_1(42059) <= 9462163;
srom_1(42060) <= 8890262;
srom_1(42061) <= 8316008;
srom_1(42062) <= 7742095;
srom_1(42063) <= 7171214;
srom_1(42064) <= 6606041;
srom_1(42065) <= 6049228;
srom_1(42066) <= 5503385;
srom_1(42067) <= 4971071;
srom_1(42068) <= 4454783;
srom_1(42069) <= 3956943;
srom_1(42070) <= 3479884;
srom_1(42071) <= 3025844;
srom_1(42072) <= 2596951;
srom_1(42073) <= 2195218;
srom_1(42074) <= 1822528;
srom_1(42075) <= 1480628;
srom_1(42076) <= 1171122;
srom_1(42077) <= 895461;
srom_1(42078) <= 654939;
srom_1(42079) <= 450682;
srom_1(42080) <= 283648;
srom_1(42081) <= 154622;
srom_1(42082) <= 64208;
srom_1(42083) <= 12829;
srom_1(42084) <= 728;
srom_1(42085) <= 27960;
srom_1(42086) <= 94398;
srom_1(42087) <= 199731;
srom_1(42088) <= 343464;
srom_1(42089) <= 524923;
srom_1(42090) <= 743258;
srom_1(42091) <= 997445;
srom_1(42092) <= 1286291;
srom_1(42093) <= 1608442;
srom_1(42094) <= 1962388;
srom_1(42095) <= 2346469;
srom_1(42096) <= 2758883;
srom_1(42097) <= 3197698;
srom_1(42098) <= 3660854;
srom_1(42099) <= 4146180;
srom_1(42100) <= 4651400;
srom_1(42101) <= 5174145;
srom_1(42102) <= 5711964;
srom_1(42103) <= 6262335;
srom_1(42104) <= 6822677;
srom_1(42105) <= 7390362;
srom_1(42106) <= 7962727;
srom_1(42107) <= 8537090;
srom_1(42108) <= 9110757;
srom_1(42109) <= 9681037;
srom_1(42110) <= 10245257;
srom_1(42111) <= 10800770;
srom_1(42112) <= 11344972;
srom_1(42113) <= 11875310;
srom_1(42114) <= 12389298;
srom_1(42115) <= 12884525;
srom_1(42116) <= 13358670;
srom_1(42117) <= 13809508;
srom_1(42118) <= 14234925;
srom_1(42119) <= 14632928;
srom_1(42120) <= 15001648;
srom_1(42121) <= 15339358;
srom_1(42122) <= 15644473;
srom_1(42123) <= 15915563;
srom_1(42124) <= 16151356;
srom_1(42125) <= 16350747;
srom_1(42126) <= 16512801;
srom_1(42127) <= 16636758;
srom_1(42128) <= 16722036;
srom_1(42129) <= 16768237;
srom_1(42130) <= 16775142;
srom_1(42131) <= 16742720;
srom_1(42132) <= 16671122;
srom_1(42133) <= 16560685;
srom_1(42134) <= 16411926;
srom_1(42135) <= 16225543;
srom_1(42136) <= 16002411;
srom_1(42137) <= 15743574;
srom_1(42138) <= 15450247;
srom_1(42139) <= 15123806;
srom_1(42140) <= 14765781;
srom_1(42141) <= 14377852;
srom_1(42142) <= 13961837;
srom_1(42143) <= 13519687;
srom_1(42144) <= 13053475;
srom_1(42145) <= 12565389;
srom_1(42146) <= 12057716;
srom_1(42147) <= 11532837;
srom_1(42148) <= 10993214;
srom_1(42149) <= 10441377;
srom_1(42150) <= 9879914;
srom_1(42151) <= 9311458;
srom_1(42152) <= 8738674;
srom_1(42153) <= 8164249;
srom_1(42154) <= 7590875;
srom_1(42155) <= 7021243;
srom_1(42156) <= 6458022;
srom_1(42157) <= 5903855;
srom_1(42158) <= 5361340;
srom_1(42159) <= 4833020;
srom_1(42160) <= 4321374;
srom_1(42161) <= 3828800;
srom_1(42162) <= 3357609;
srom_1(42163) <= 2910010;
srom_1(42164) <= 2488102;
srom_1(42165) <= 2093864;
srom_1(42166) <= 1729144;
srom_1(42167) <= 1395652;
srom_1(42168) <= 1094953;
srom_1(42169) <= 828456;
srom_1(42170) <= 597411;
srom_1(42171) <= 402902;
srom_1(42172) <= 245840;
srom_1(42173) <= 126963;
srom_1(42174) <= 46827;
srom_1(42175) <= 5809;
srom_1(42176) <= 4101;
srom_1(42177) <= 41711;
srom_1(42178) <= 118462;
srom_1(42179) <= 233994;
srom_1(42180) <= 387766;
srom_1(42181) <= 579057;
srom_1(42182) <= 806970;
srom_1(42183) <= 1070436;
srom_1(42184) <= 1368219;
srom_1(42185) <= 1698923;
srom_1(42186) <= 2060997;
srom_1(42187) <= 2452744;
srom_1(42188) <= 2872325;
srom_1(42189) <= 3317775;
srom_1(42190) <= 3787004;
srom_1(42191) <= 4277810;
srom_1(42192) <= 4787894;
srom_1(42193) <= 5314863;
srom_1(42194) <= 5856246;
srom_1(42195) <= 6409504;
srom_1(42196) <= 6972042;
srom_1(42197) <= 7541224;
srom_1(42198) <= 8114379;
srom_1(42199) <= 8688819;
srom_1(42200) <= 9261853;
srom_1(42201) <= 9830791;
srom_1(42202) <= 10392966;
srom_1(42203) <= 10945742;
srom_1(42204) <= 11486527;
srom_1(42205) <= 12012785;
srom_1(42206) <= 12522047;
srom_1(42207) <= 13011927;
srom_1(42208) <= 13480126;
srom_1(42209) <= 13924449;
srom_1(42210) <= 14342813;
srom_1(42211) <= 14733255;
srom_1(42212) <= 15093946;
srom_1(42213) <= 15423192;
srom_1(42214) <= 15719451;
srom_1(42215) <= 15981333;
srom_1(42216) <= 16207611;
srom_1(42217) <= 16397222;
srom_1(42218) <= 16549278;
srom_1(42219) <= 16663066;
srom_1(42220) <= 16738052;
srom_1(42221) <= 16773885;
srom_1(42222) <= 16770396;
srom_1(42223) <= 16727602;
srom_1(42224) <= 16645704;
srom_1(42225) <= 16525085;
srom_1(42226) <= 16366312;
srom_1(42227) <= 16170128;
srom_1(42228) <= 15937455;
srom_1(42229) <= 15669382;
srom_1(42230) <= 15367167;
srom_1(42231) <= 15032227;
srom_1(42232) <= 14666133;
srom_1(42233) <= 14270601;
srom_1(42234) <= 13847487;
srom_1(42235) <= 13398774;
srom_1(42236) <= 12926567;
srom_1(42237) <= 12433080;
srom_1(42238) <= 11920627;
srom_1(42239) <= 11391611;
srom_1(42240) <= 10848512;
srom_1(42241) <= 10293879;
srom_1(42242) <= 9730311;
srom_1(42243) <= 9160451;
srom_1(42244) <= 8586972;
srom_1(42245) <= 8012563;
srom_1(42246) <= 7439917;
srom_1(42247) <= 6871720;
srom_1(42248) <= 6310636;
srom_1(42249) <= 5759296;
srom_1(42250) <= 5220286;
srom_1(42251) <= 4696133;
srom_1(42252) <= 4189296;
srom_1(42253) <= 3702151;
srom_1(42254) <= 3236982;
srom_1(42255) <= 2795971;
srom_1(42256) <= 2381185;
srom_1(42257) <= 1994571;
srom_1(42258) <= 1637940;
srom_1(42259) <= 1312966;
srom_1(42260) <= 1021171;
srom_1(42261) <= 763925;
srom_1(42262) <= 542434;
srom_1(42263) <= 357736;
srom_1(42264) <= 210698;
srom_1(42265) <= 102009;
srom_1(42266) <= 32178;
srom_1(42267) <= 1534;
srom_1(42268) <= 10219;
srom_1(42269) <= 58194;
srom_1(42270) <= 145233;
srom_1(42271) <= 270927;
srom_1(42272) <= 434689;
srom_1(42273) <= 635749;
srom_1(42274) <= 873165;
srom_1(42275) <= 1145823;
srom_1(42276) <= 1452445;
srom_1(42277) <= 1791593;
srom_1(42278) <= 2161677;
srom_1(42279) <= 2560961;
srom_1(42280) <= 2987573;
srom_1(42281) <= 3439513;
srom_1(42282) <= 3914660;
srom_1(42283) <= 4410787;
srom_1(42284) <= 4925568;
srom_1(42285) <= 5456588;
srom_1(42286) <= 6001357;
srom_1(42287) <= 6557320;
srom_1(42288) <= 7121872;
srom_1(42289) <= 7692363;
srom_1(42290) <= 8266120;
srom_1(42291) <= 8840450;
srom_1(42292) <= 9412662;
srom_1(42293) <= 9980072;
srom_1(42294) <= 10540019;
srom_1(42295) <= 11089877;
srom_1(42296) <= 11627068;
srom_1(42297) <= 12149072;
srom_1(42298) <= 12653443;
srom_1(42299) <= 13137814;
srom_1(42300) <= 13599915;
srom_1(42301) <= 14037578;
srom_1(42302) <= 14448751;
srom_1(42303) <= 14831506;
srom_1(42304) <= 15184048;
srom_1(42305) <= 15504724;
srom_1(42306) <= 15792030;
srom_1(42307) <= 16044618;
srom_1(42308) <= 16261305;
srom_1(42309) <= 16441074;
srom_1(42310) <= 16583083;
srom_1(42311) <= 16686665;
srom_1(42312) <= 16751334;
srom_1(42313) <= 16776787;
srom_1(42314) <= 16762906;
srom_1(42315) <= 16709755;
srom_1(42316) <= 16617582;
srom_1(42317) <= 16486822;
srom_1(42318) <= 16318086;
srom_1(42319) <= 16112166;
srom_1(42320) <= 15870027;
srom_1(42321) <= 15592806;
srom_1(42322) <= 15281801;
srom_1(42323) <= 14938472;
srom_1(42324) <= 14564429;
srom_1(42325) <= 14161425;
srom_1(42326) <= 13731350;
srom_1(42327) <= 13276221;
srom_1(42328) <= 12798173;
srom_1(42329) <= 12299446;
srom_1(42330) <= 11782381;
srom_1(42331) <= 11249401;
srom_1(42332) <= 10703005;
srom_1(42333) <= 10145756;
srom_1(42334) <= 9580268;
srom_1(42335) <= 9009192;
srom_1(42336) <= 8435205;
srom_1(42337) <= 7861000;
srom_1(42338) <= 7289269;
srom_1(42339) <= 6722693;
srom_1(42340) <= 6163929;
srom_1(42341) <= 5615597;
srom_1(42342) <= 5080269;
srom_1(42343) <= 4560455;
srom_1(42344) <= 4058593;
srom_1(42345) <= 3577035;
srom_1(42346) <= 3118041;
srom_1(42347) <= 2683762;
srom_1(42348) <= 2276235;
srom_1(42349) <= 1897371;
srom_1(42350) <= 1548946;
srom_1(42351) <= 1232596;
srom_1(42352) <= 949802;
srom_1(42353) <= 701891;
srom_1(42354) <= 490026;
srom_1(42355) <= 315200;
srom_1(42356) <= 178233;
srom_1(42357) <= 79767;
srom_1(42358) <= 20265;
srom_1(42359) <= 4;
srom_1(42360) <= 19080;
srom_1(42361) <= 77404;
srom_1(42362) <= 174702;
srom_1(42363) <= 310518;
srom_1(42364) <= 484215;
srom_1(42365) <= 694978;
srom_1(42366) <= 941819;
srom_1(42367) <= 1223581;
srom_1(42368) <= 1538942;
srom_1(42369) <= 1886424;
srom_1(42370) <= 2264396;
srom_1(42371) <= 2671087;
srom_1(42372) <= 3104590;
srom_1(42373) <= 3562871;
srom_1(42374) <= 4043781;
srom_1(42375) <= 4545066;
srom_1(42376) <= 5064375;
srom_1(42377) <= 5599272;
srom_1(42378) <= 6147249;
srom_1(42379) <= 6705736;
srom_1(42380) <= 7272116;
srom_1(42381) <= 7843731;
srom_1(42382) <= 8417901;
srom_1(42383) <= 8991933;
srom_1(42384) <= 9563136;
srom_1(42385) <= 10128832;
srom_1(42386) <= 10686367;
srom_1(42387) <= 11233127;
srom_1(42388) <= 11766548;
srom_1(42389) <= 12284129;
srom_1(42390) <= 12783443;
srom_1(42391) <= 13262147;
srom_1(42392) <= 13717998;
srom_1(42393) <= 14148857;
srom_1(42394) <= 14552705;
srom_1(42395) <= 14927647;
srom_1(42396) <= 15271925;
srom_1(42397) <= 15583925;
srom_1(42398) <= 15862184;
srom_1(42399) <= 16105397;
srom_1(42400) <= 16312422;
srom_1(42401) <= 16482291;
srom_1(42402) <= 16614205;
srom_1(42403) <= 16707547;
srom_1(42404) <= 16761878;
srom_1(42405) <= 16776944;
srom_1(42406) <= 16752674;
srom_1(42407) <= 16689183;
srom_1(42408) <= 16586767;
srom_1(42409) <= 16445907;
srom_1(42410) <= 16267263;
srom_1(42411) <= 16051674;
srom_1(42412) <= 15800150;
srom_1(42413) <= 15513871;
srom_1(42414) <= 15194179;
srom_1(42415) <= 14842574;
srom_1(42416) <= 14460703;
srom_1(42417) <= 14050359;
srom_1(42418) <= 13613464;
srom_1(42419) <= 13152068;
srom_1(42420) <= 12668335;
srom_1(42421) <= 12164533;
srom_1(42422) <= 11643024;
srom_1(42423) <= 11106254;
srom_1(42424) <= 10556740;
srom_1(42425) <= 9997059;
srom_1(42426) <= 9429835;
srom_1(42427) <= 8857729;
srom_1(42428) <= 8283422;
srom_1(42429) <= 7709609;
srom_1(42430) <= 7138980;
srom_1(42431) <= 6574211;
srom_1(42432) <= 6017951;
srom_1(42433) <= 5472807;
srom_1(42434) <= 4941336;
srom_1(42435) <= 4426031;
srom_1(42436) <= 3929307;
srom_1(42437) <= 3453495;
srom_1(42438) <= 3000825;
srom_1(42439) <= 2573421;
srom_1(42440) <= 2173286;
srom_1(42441) <= 1802296;
srom_1(42442) <= 1462192;
srom_1(42443) <= 1154569;
srom_1(42444) <= 880868;
srom_1(42445) <= 642373;
srom_1(42446) <= 440204;
srom_1(42447) <= 275307;
srom_1(42448) <= 148456;
srom_1(42449) <= 60246;
srom_1(42450) <= 11091;
srom_1(42451) <= 1221;
srom_1(42452) <= 30682;
srom_1(42453) <= 99336;
srom_1(42454) <= 206861;
srom_1(42455) <= 352754;
srom_1(42456) <= 536329;
srom_1(42457) <= 756726;
srom_1(42458) <= 1012912;
srom_1(42459) <= 1303685;
srom_1(42460) <= 1627682;
srom_1(42461) <= 1983383;
srom_1(42462) <= 2369120;
srom_1(42463) <= 2783085;
srom_1(42464) <= 3223336;
srom_1(42465) <= 3687808;
srom_1(42466) <= 4174325;
srom_1(42467) <= 4680603;
srom_1(42468) <= 5204270;
srom_1(42469) <= 5742869;
srom_1(42470) <= 6293875;
srom_1(42471) <= 6854704;
srom_1(42472) <= 7422725;
srom_1(42473) <= 7995276;
srom_1(42474) <= 8569672;
srom_1(42475) <= 9143218;
srom_1(42476) <= 9713226;
srom_1(42477) <= 10277023;
srom_1(42478) <= 10831963;
srom_1(42479) <= 11375446;
srom_1(42480) <= 11904923;
srom_1(42481) <= 12417911;
srom_1(42482) <= 12912003;
srom_1(42483) <= 13384884;
srom_1(42484) <= 13834336;
srom_1(42485) <= 14258251;
srom_1(42486) <= 14654641;
srom_1(42487) <= 15021648;
srom_1(42488) <= 15357549;
srom_1(42489) <= 15660771;
srom_1(42490) <= 15929892;
srom_1(42491) <= 16163649;
srom_1(42492) <= 16360945;
srom_1(42493) <= 16520857;
srom_1(42494) <= 16642634;
srom_1(42495) <= 16725705;
srom_1(42496) <= 16769681;
srom_1(42497) <= 16774354;
srom_1(42498) <= 16739704;
srom_1(42499) <= 16665893;
srom_1(42500) <= 16553267;
srom_1(42501) <= 16402354;
srom_1(42502) <= 16213862;
srom_1(42503) <= 15988674;
srom_1(42504) <= 15727847;
srom_1(42505) <= 15432604;
srom_1(42506) <= 15104329;
srom_1(42507) <= 14744562;
srom_1(42508) <= 14354990;
srom_1(42509) <= 13937439;
srom_1(42510) <= 13493867;
srom_1(42511) <= 13026356;
srom_1(42512) <= 12537096;
srom_1(42513) <= 12028383;
srom_1(42514) <= 11502602;
srom_1(42515) <= 10962218;
srom_1(42516) <= 10409765;
srom_1(42517) <= 9847835;
srom_1(42518) <= 9279061;
srom_1(42519) <= 8706112;
srom_1(42520) <= 8131674;
srom_1(42521) <= 7558441;
srom_1(42522) <= 6989101;
srom_1(42523) <= 6426324;
srom_1(42524) <= 5872749;
srom_1(42525) <= 5330971;
srom_1(42526) <= 4803531;
srom_1(42527) <= 4292904;
srom_1(42528) <= 3801482;
srom_1(42529) <= 3331571;
srom_1(42530) <= 2885374;
srom_1(42531) <= 2464984;
srom_1(42532) <= 2072371;
srom_1(42533) <= 1709378;
srom_1(42534) <= 1377706;
srom_1(42535) <= 1078910;
srom_1(42536) <= 814392;
srom_1(42537) <= 585392;
srom_1(42538) <= 392984;
srom_1(42539) <= 238070;
srom_1(42540) <= 121377;
srom_1(42541) <= 43452;
srom_1(42542) <= 4660;
srom_1(42543) <= 5183;
srom_1(42544) <= 45019;
srom_1(42545) <= 123981;
srom_1(42546) <= 241699;
srom_1(42547) <= 397620;
srom_1(42548) <= 591014;
srom_1(42549) <= 820973;
srom_1(42550) <= 1086420;
srom_1(42551) <= 1386109;
srom_1(42552) <= 1718635;
srom_1(42553) <= 2082439;
srom_1(42554) <= 2475815;
srom_1(42555) <= 2896918;
srom_1(42556) <= 3343773;
srom_1(42557) <= 3814285;
srom_1(42558) <= 4306248;
srom_1(42559) <= 4817355;
srom_1(42560) <= 5345208;
srom_1(42561) <= 5887333;
srom_1(42562) <= 6441187;
srom_1(42563) <= 7004173;
srom_1(42564) <= 7573651;
srom_1(42565) <= 8146951;
srom_1(42566) <= 8721384;
srom_1(42567) <= 9294257;
srom_1(42568) <= 9862882;
srom_1(42569) <= 10424595;
srom_1(42570) <= 10976760;
srom_1(42571) <= 11516788;
srom_1(42572) <= 12042147;
srom_1(42573) <= 12550373;
srom_1(42574) <= 13039083;
srom_1(42575) <= 13505986;
srom_1(42576) <= 13948891;
srom_1(42577) <= 14365723;
srom_1(42578) <= 14754526;
srom_1(42579) <= 15113476;
srom_1(42580) <= 15440892;
srom_1(42581) <= 15735237;
srom_1(42582) <= 15995131;
srom_1(42583) <= 16219355;
srom_1(42584) <= 16406858;
srom_1(42585) <= 16556761;
srom_1(42586) <= 16668361;
srom_1(42587) <= 16741134;
srom_1(42588) <= 16774739;
srom_1(42589) <= 16769019;
srom_1(42590) <= 16724000;
srom_1(42591) <= 16639894;
srom_1(42592) <= 16517094;
srom_1(42593) <= 16356178;
srom_1(42594) <= 16157898;
srom_1(42595) <= 15923186;
srom_1(42596) <= 15653141;
srom_1(42597) <= 15349031;
srom_1(42598) <= 15012280;
srom_1(42599) <= 14644469;
srom_1(42600) <= 14247323;
srom_1(42601) <= 13822702;
srom_1(42602) <= 13372599;
srom_1(42603) <= 12899125;
srom_1(42604) <= 12404499;
srom_1(42605) <= 11891042;
srom_1(42606) <= 11361160;
srom_1(42607) <= 10817339;
srom_1(42608) <= 10262128;
srom_1(42609) <= 9698133;
srom_1(42610) <= 9127996;
srom_1(42611) <= 8554392;
srom_1(42612) <= 7980011;
srom_1(42613) <= 7407545;
srom_1(42614) <= 6839680;
srom_1(42615) <= 6279079;
srom_1(42616) <= 5728370;
srom_1(42617) <= 5190136;
srom_1(42618) <= 4666900;
srom_1(42619) <= 4161117;
srom_1(42620) <= 3675158;
srom_1(42621) <= 3211302;
srom_1(42622) <= 2771724;
srom_1(42623) <= 2358486;
srom_1(42624) <= 1973525;
srom_1(42625) <= 1618646;
srom_1(42626) <= 1295514;
srom_1(42627) <= 1005644;
srom_1(42628) <= 750396;
srom_1(42629) <= 530965;
srom_1(42630) <= 348382;
srom_1(42631) <= 203502;
srom_1(42632) <= 97005;
srom_1(42633) <= 29390;
srom_1(42634) <= 974;
srom_1(42635) <= 11890;
srom_1(42636) <= 62088;
srom_1(42637) <= 151332;
srom_1(42638) <= 279204;
srom_1(42639) <= 445103;
srom_1(42640) <= 648252;
srom_1(42641) <= 887698;
srom_1(42642) <= 1162318;
srom_1(42643) <= 1470825;
srom_1(42644) <= 1811772;
srom_1(42645) <= 2183560;
srom_1(42646) <= 2584445;
srom_1(42647) <= 3012549;
srom_1(42648) <= 3465862;
srom_1(42649) <= 3942260;
srom_1(42650) <= 4439508;
srom_1(42651) <= 4955275;
srom_1(42652) <= 5487142;
srom_1(42653) <= 6032615;
srom_1(42654) <= 6589136;
srom_1(42655) <= 7154095;
srom_1(42656) <= 7724844;
srom_1(42657) <= 8298705;
srom_1(42658) <= 8872987;
srom_1(42659) <= 9444998;
srom_1(42660) <= 10012056;
srom_1(42661) <= 10571500;
srom_1(42662) <= 11120708;
srom_1(42663) <= 11657105;
srom_1(42664) <= 12178174;
srom_1(42665) <= 12681473;
srom_1(42666) <= 13164641;
srom_1(42667) <= 13625412;
srom_1(42668) <= 14061626;
srom_1(42669) <= 14471238;
srom_1(42670) <= 14852326;
srom_1(42671) <= 15203103;
srom_1(42672) <= 15521925;
srom_1(42673) <= 15807297;
srom_1(42674) <= 16057879;
srom_1(42675) <= 16272498;
srom_1(42676) <= 16450146;
srom_1(42677) <= 16589991;
srom_1(42678) <= 16691377;
srom_1(42679) <= 16753829;
srom_1(42680) <= 16777053;
srom_1(42681) <= 16760940;
srom_1(42682) <= 16705567;
srom_1(42683) <= 16611193;
srom_1(42684) <= 16478260;
srom_1(42685) <= 16307393;
srom_1(42686) <= 16099391;
srom_1(42687) <= 15855231;
srom_1(42688) <= 15576057;
srom_1(42689) <= 15263179;
srom_1(42690) <= 14918063;
srom_1(42691) <= 14542329;
srom_1(42692) <= 14137737;
srom_1(42693) <= 13706187;
srom_1(42694) <= 13249700;
srom_1(42695) <= 12770417;
srom_1(42696) <= 12270587;
srom_1(42697) <= 11752553;
srom_1(42698) <= 11218745;
srom_1(42699) <= 10671665;
srom_1(42700) <= 10113878;
srom_1(42701) <= 9548002;
srom_1(42702) <= 8976688;
srom_1(42703) <= 8402617;
srom_1(42704) <= 7828480;
srom_1(42705) <= 7256970;
srom_1(42706) <= 6690767;
srom_1(42707) <= 6132525;
srom_1(42708) <= 5584863;
srom_1(42709) <= 5050348;
srom_1(42710) <= 4531488;
srom_1(42711) <= 4030715;
srom_1(42712) <= 3550377;
srom_1(42713) <= 3092728;
srom_1(42714) <= 2659913;
srom_1(42715) <= 2253962;
srom_1(42716) <= 1876778;
srom_1(42717) <= 1530131;
srom_1(42718) <= 1215645;
srom_1(42719) <= 934796;
srom_1(42720) <= 688900;
srom_1(42721) <= 479111;
srom_1(42722) <= 306412;
srom_1(42723) <= 171613;
srom_1(42724) <= 75347;
srom_1(42725) <= 18064;
srom_1(42726) <= 34;
srom_1(42727) <= 21340;
srom_1(42728) <= 81884;
srom_1(42729) <= 181380;
srom_1(42730) <= 319364;
srom_1(42731) <= 495186;
srom_1(42732) <= 708024;
srom_1(42733) <= 956878;
srom_1(42734) <= 1240582;
srom_1(42735) <= 1557806;
srom_1(42736) <= 1907062;
srom_1(42737) <= 2286712;
srom_1(42738) <= 2694976;
srom_1(42739) <= 3129940;
srom_1(42740) <= 3589563;
srom_1(42741) <= 4071690;
srom_1(42742) <= 4574061;
srom_1(42743) <= 5094319;
srom_1(42744) <= 5630026;
srom_1(42745) <= 6178669;
srom_1(42746) <= 6737674;
srom_1(42747) <= 7304422;
srom_1(42748) <= 7876254;
srom_1(42749) <= 8450488;
srom_1(42750) <= 9024432;
srom_1(42751) <= 9595394;
srom_1(42752) <= 10160698;
srom_1(42753) <= 10717691;
srom_1(42754) <= 11263763;
srom_1(42755) <= 11796352;
srom_1(42756) <= 12312961;
srom_1(42757) <= 12811167;
srom_1(42758) <= 13288634;
srom_1(42759) <= 13743124;
srom_1(42760) <= 14172504;
srom_1(42761) <= 14574762;
srom_1(42762) <= 14948010;
srom_1(42763) <= 15290499;
srom_1(42764) <= 15600623;
srom_1(42765) <= 15876928;
srom_1(42766) <= 16118117;
srom_1(42767) <= 16323059;
srom_1(42768) <= 16490795;
srom_1(42769) <= 16620536;
srom_1(42770) <= 16711675;
srom_1(42771) <= 16763784;
srom_1(42772) <= 16776620;
srom_1(42773) <= 16750120;
srom_1(42774) <= 16684411;
srom_1(42775) <= 16579800;
srom_1(42776) <= 16436778;
srom_1(42777) <= 16256015;
srom_1(42778) <= 16038359;
srom_1(42779) <= 15784831;
srom_1(42780) <= 15496619;
srom_1(42781) <= 15175076;
srom_1(42782) <= 14821708;
srom_1(42783) <= 14438173;
srom_1(42784) <= 14026270;
srom_1(42785) <= 13587930;
srom_1(42786) <= 13125208;
srom_1(42787) <= 12640275;
srom_1(42788) <= 12135405;
srom_1(42789) <= 11612964;
srom_1(42790) <= 11075403;
srom_1(42791) <= 10525243;
srom_1(42792) <= 9965064;
srom_1(42793) <= 9397491;
srom_1(42794) <= 8825188;
srom_1(42795) <= 8250838;
srom_1(42796) <= 7677134;
srom_1(42797) <= 7106766;
srom_1(42798) <= 6542409;
srom_1(42799) <= 5986709;
srom_1(42800) <= 5442273;
srom_1(42801) <= 4911653;
srom_1(42802) <= 4397338;
srom_1(42803) <= 3901739;
srom_1(42804) <= 3427181;
srom_1(42805) <= 2975888;
srom_1(42806) <= 2549978;
srom_1(42807) <= 2151447;
srom_1(42808) <= 1782164;
srom_1(42809) <= 1443861;
srom_1(42810) <= 1138124;
srom_1(42811) <= 866388;
srom_1(42812) <= 629925;
srom_1(42813) <= 429846;
srom_1(42814) <= 267088;
srom_1(42815) <= 142415;
srom_1(42816) <= 56410;
srom_1(42817) <= 9479;
srom_1(42818) <= 1840;
srom_1(42819) <= 33529;
srom_1(42820) <= 104399;
srom_1(42821) <= 214115;
srom_1(42822) <= 362165;
srom_1(42823) <= 547854;
srom_1(42824) <= 770310;
srom_1(42825) <= 1028491;
srom_1(42826) <= 1321187;
srom_1(42827) <= 1647024;
srom_1(42828) <= 2004474;
srom_1(42829) <= 2391862;
srom_1(42830) <= 2807371;
srom_1(42831) <= 3249052;
srom_1(42832) <= 3714834;
srom_1(42833) <= 4202533;
srom_1(42834) <= 4709863;
srom_1(42835) <= 5234442;
srom_1(42836) <= 5773813;
srom_1(42837) <= 6325446;
srom_1(42838) <= 6886753;
srom_1(42839) <= 7455104;
srom_1(42840) <= 8027831;
srom_1(42841) <= 8602251;
srom_1(42842) <= 9175668;
srom_1(42843) <= 9745395;
srom_1(42844) <= 10308760;
srom_1(42845) <= 10863120;
srom_1(42846) <= 11405876;
srom_1(42847) <= 11934483;
srom_1(42848) <= 12446463;
srom_1(42849) <= 12939413;
srom_1(42850) <= 13411024;
srom_1(42851) <= 13859082;
srom_1(42852) <= 14281488;
srom_1(42853) <= 14676260;
srom_1(42854) <= 15041547;
srom_1(42855) <= 15375636;
srom_1(42856) <= 15676960;
srom_1(42857) <= 15944107;
srom_1(42858) <= 16175824;
srom_1(42859) <= 16371023;
srom_1(42860) <= 16528791;
srom_1(42861) <= 16648386;
srom_1(42862) <= 16729248;
srom_1(42863) <= 16770998;
srom_1(42864) <= 16773440;
srom_1(42865) <= 16736563;
srom_1(42866) <= 16660539;
srom_1(42867) <= 16545726;
srom_1(42868) <= 16392661;
srom_1(42869) <= 16202062;
srom_1(42870) <= 15974823;
srom_1(42871) <= 15712010;
srom_1(42872) <= 15414855;
srom_1(42873) <= 15084751;
srom_1(42874) <= 14723247;
srom_1(42875) <= 14332037;
srom_1(42876) <= 13912957;
srom_1(42877) <= 13467971;
srom_1(42878) <= 12999166;
srom_1(42879) <= 12508741;
srom_1(42880) <= 11998995;
srom_1(42881) <= 11472319;
srom_1(42882) <= 10931182;
srom_1(42883) <= 10378122;
srom_1(42884) <= 9815733;
srom_1(42885) <= 9246651;
srom_1(42886) <= 8673545;
srom_1(42887) <= 8099104;
srom_1(42888) <= 7526020;
srom_1(42889) <= 6956981;
srom_1(42890) <= 6394655;
srom_1(42891) <= 5841680;
srom_1(42892) <= 5300648;
srom_1(42893) <= 4774097;
srom_1(42894) <= 4264495;
srom_1(42895) <= 3774233;
srom_1(42896) <= 3305609;
srom_1(42897) <= 2860821;
srom_1(42898) <= 2441954;
srom_1(42899) <= 2050974;
srom_1(42900) <= 1689713;
srom_1(42901) <= 1359865;
srom_1(42902) <= 1062977;
srom_1(42903) <= 800442;
srom_1(42904) <= 573491;
srom_1(42905) <= 383187;
srom_1(42906) <= 230423;
srom_1(42907) <= 115916;
srom_1(42908) <= 40202;
srom_1(42909) <= 3637;
srom_1(42910) <= 6392;
srom_1(42911) <= 48454;
srom_1(42912) <= 129626;
srom_1(42913) <= 249527;
srom_1(42914) <= 407595;
srom_1(42915) <= 603088;
srom_1(42916) <= 835091;
srom_1(42917) <= 1102514;
srom_1(42918) <= 1404105;
srom_1(42919) <= 1738448;
srom_1(42920) <= 2103977;
srom_1(42921) <= 2498976;
srom_1(42922) <= 2921593;
srom_1(42923) <= 3369847;
srom_1(42924) <= 3841636;
srom_1(42925) <= 4334747;
srom_1(42926) <= 4846869;
srom_1(42927) <= 5375598;
srom_1(42928) <= 5918457;
srom_1(42929) <= 6472899;
srom_1(42930) <= 7036324;
srom_1(42931) <= 7606091;
srom_1(42932) <= 8179527;
srom_1(42933) <= 8753944;
srom_1(42934) <= 9326647;
srom_1(42935) <= 9894952;
srom_1(42936) <= 10456193;
srom_1(42937) <= 11007738;
srom_1(42938) <= 11547001;
srom_1(42939) <= 12071454;
srom_1(42940) <= 12578636;
srom_1(42941) <= 13066170;
srom_1(42942) <= 13531769;
srom_1(42943) <= 13973250;
srom_1(42944) <= 14388543;
srom_1(42945) <= 14775700;
srom_1(42946) <= 15132906;
srom_1(42947) <= 15458485;
srom_1(42948) <= 15750911;
srom_1(42949) <= 16008813;
srom_1(42950) <= 16230981;
srom_1(42951) <= 16416374;
srom_1(42952) <= 16564122;
srom_1(42953) <= 16673531;
srom_1(42954) <= 16744090;
srom_1(42955) <= 16775468;
srom_1(42956) <= 16767516;
srom_1(42957) <= 16720273;
srom_1(42958) <= 16633959;
srom_1(42959) <= 16508981;
srom_1(42960) <= 16345923;
srom_1(42961) <= 16145551;
srom_1(42962) <= 15908803;
srom_1(42963) <= 15636791;
srom_1(42964) <= 15330790;
srom_1(42965) <= 14992234;
srom_1(42966) <= 14622712;
srom_1(42967) <= 14223955;
srom_1(42968) <= 13797835;
srom_1(42969) <= 13346349;
srom_1(42970) <= 12871615;
srom_1(42971) <= 12375858;
srom_1(42972) <= 11861404;
srom_1(42973) <= 11330664;
srom_1(42974) <= 10786128;
srom_1(42975) <= 10230350;
srom_1(42976) <= 9665934;
srom_1(42977) <= 9095529;
srom_1(42978) <= 8521809;
srom_1(42979) <= 7947465;
srom_1(42980) <= 7375189;
srom_1(42981) <= 6807665;
srom_1(42982) <= 6247555;
srom_1(42983) <= 5697485;
srom_1(42984) <= 5160034;
srom_1(42985) <= 4637723;
srom_1(42986) <= 4133002;
srom_1(42987) <= 3648237;
srom_1(42988) <= 3185700;
srom_1(42989) <= 2747562;
srom_1(42990) <= 2335877;
srom_1(42991) <= 1952575;
srom_1(42992) <= 1599454;
srom_1(42993) <= 1278170;
srom_1(42994) <= 990229;
srom_1(42995) <= 736981;
srom_1(42996) <= 519615;
srom_1(42997) <= 339149;
srom_1(42998) <= 196429;
srom_1(42999) <= 92126;
srom_1(43000) <= 26727;
srom_1(43001) <= 540;
srom_1(43002) <= 13688;
srom_1(43003) <= 66109;
srom_1(43004) <= 157557;
srom_1(43005) <= 287603;
srom_1(43006) <= 455637;
srom_1(43007) <= 660872;
srom_1(43008) <= 902344;
srom_1(43009) <= 1178923;
srom_1(43010) <= 1489310;
srom_1(43011) <= 1832050;
srom_1(43012) <= 2205536;
srom_1(43013) <= 2608017;
srom_1(43014) <= 3037605;
srom_1(43015) <= 3492286;
srom_1(43016) <= 3969927;
srom_1(43017) <= 4468289;
srom_1(43018) <= 4985034;
srom_1(43019) <= 5517740;
srom_1(43020) <= 6063909;
srom_1(43021) <= 6620979;
srom_1(43022) <= 7186338;
srom_1(43023) <= 7757334;
srom_1(43024) <= 8331291;
srom_1(43025) <= 8905517;
srom_1(43026) <= 9477319;
srom_1(43027) <= 10044015;
srom_1(43028) <= 10602949;
srom_1(43029) <= 11151499;
srom_1(43030) <= 11687092;
srom_1(43031) <= 12207218;
srom_1(43032) <= 12709438;
srom_1(43033) <= 13191395;
srom_1(43034) <= 13650830;
srom_1(43035) <= 14085589;
srom_1(43036) <= 14493633;
srom_1(43037) <= 14873049;
srom_1(43038) <= 15222056;
srom_1(43039) <= 15539019;
srom_1(43040) <= 15822452;
srom_1(43041) <= 16071024;
srom_1(43042) <= 16283571;
srom_1(43043) <= 16459096;
srom_1(43044) <= 16596776;
srom_1(43045) <= 16695964;
srom_1(43046) <= 16756197;
srom_1(43047) <= 16777191;
srom_1(43048) <= 16758848;
srom_1(43049) <= 16701254;
srom_1(43050) <= 16604680;
srom_1(43051) <= 16469577;
srom_1(43052) <= 16296580;
srom_1(43053) <= 16086500;
srom_1(43054) <= 15840321;
srom_1(43055) <= 15559199;
srom_1(43056) <= 15244452;
srom_1(43057) <= 14897555;
srom_1(43058) <= 14520136;
srom_1(43059) <= 14113963;
srom_1(43060) <= 13680943;
srom_1(43061) <= 13223105;
srom_1(43062) <= 12742596;
srom_1(43063) <= 12241670;
srom_1(43064) <= 11722675;
srom_1(43065) <= 11188046;
srom_1(43066) <= 10640290;
srom_1(43067) <= 10081974;
srom_1(43068) <= 9515718;
srom_1(43069) <= 8944176;
srom_1(43070) <= 8370029;
srom_1(43071) <= 7795970;
srom_1(43072) <= 7224689;
srom_1(43073) <= 6658866;
srom_1(43074) <= 6101155;
srom_1(43075) <= 5554170;
srom_1(43076) <= 5020477;
srom_1(43077) <= 4502578;
srom_1(43078) <= 4002902;
srom_1(43079) <= 3523793;
srom_1(43080) <= 3067496;
srom_1(43081) <= 2636151;
srom_1(43082) <= 2231782;
srom_1(43083) <= 1856284;
srom_1(43084) <= 1511419;
srom_1(43085) <= 1198803;
srom_1(43086) <= 919902;
srom_1(43087) <= 676025;
srom_1(43088) <= 468315;
srom_1(43089) <= 297746;
srom_1(43090) <= 165117;
srom_1(43091) <= 71051;
srom_1(43092) <= 15990;
srom_1(43093) <= 190;
srom_1(43094) <= 23726;
srom_1(43095) <= 86489;
srom_1(43096) <= 188182;
srom_1(43097) <= 328331;
srom_1(43098) <= 506276;
srom_1(43099) <= 721185;
srom_1(43100) <= 972049;
srom_1(43101) <= 1257692;
srom_1(43102) <= 1576774;
srom_1(43103) <= 1927798;
srom_1(43104) <= 2309120;
srom_1(43105) <= 2718951;
srom_1(43106) <= 3155369;
srom_1(43107) <= 3616327;
srom_1(43108) <= 4099664;
srom_1(43109) <= 4603113;
srom_1(43110) <= 5124314;
srom_1(43111) <= 5660822;
srom_1(43112) <= 6210122;
srom_1(43113) <= 6769637;
srom_1(43114) <= 7336745;
srom_1(43115) <= 7908784;
srom_1(43116) <= 8483074;
srom_1(43117) <= 9056921;
srom_1(43118) <= 9627634;
srom_1(43119) <= 10192537;
srom_1(43120) <= 10748980;
srom_1(43121) <= 11294355;
srom_1(43122) <= 11826104;
srom_1(43123) <= 12341733;
srom_1(43124) <= 12838825;
srom_1(43125) <= 13315048;
srom_1(43126) <= 13768169;
srom_1(43127) <= 14196063;
srom_1(43128) <= 14596725;
srom_1(43129) <= 14968274;
srom_1(43130) <= 15308969;
srom_1(43131) <= 15617213;
srom_1(43132) <= 15891558;
srom_1(43133) <= 16130720;
srom_1(43134) <= 16333577;
srom_1(43135) <= 16499176;
srom_1(43136) <= 16626743;
srom_1(43137) <= 16715678;
srom_1(43138) <= 16765564;
srom_1(43139) <= 16776168;
srom_1(43140) <= 16747440;
srom_1(43141) <= 16679515;
srom_1(43142) <= 16572710;
srom_1(43143) <= 16427528;
srom_1(43144) <= 16244648;
srom_1(43145) <= 16024929;
srom_1(43146) <= 15769400;
srom_1(43147) <= 15479260;
srom_1(43148) <= 15155870;
srom_1(43149) <= 14800745;
srom_1(43150) <= 14415552;
srom_1(43151) <= 14002096;
srom_1(43152) <= 13562317;
srom_1(43153) <= 13098277;
srom_1(43154) <= 12612151;
srom_1(43155) <= 12106220;
srom_1(43156) <= 11582855;
srom_1(43157) <= 11044512;
srom_1(43158) <= 10493714;
srom_1(43159) <= 9933045;
srom_1(43160) <= 9365133;
srom_1(43161) <= 8792642;
srom_1(43162) <= 8218256;
srom_1(43163) <= 7644669;
srom_1(43164) <= 7074570;
srom_1(43165) <= 6510634;
srom_1(43166) <= 5955504;
srom_1(43167) <= 5411784;
srom_1(43168) <= 4882023;
srom_1(43169) <= 4368705;
srom_1(43170) <= 3874239;
srom_1(43171) <= 3400941;
srom_1(43172) <= 2951033;
srom_1(43173) <= 2526623;
srom_1(43174) <= 2129702;
srom_1(43175) <= 1762132;
srom_1(43176) <= 1425635;
srom_1(43177) <= 1121790;
srom_1(43178) <= 852021;
srom_1(43179) <= 617594;
srom_1(43180) <= 419608;
srom_1(43181) <= 258992;
srom_1(43182) <= 136498;
srom_1(43183) <= 52700;
srom_1(43184) <= 7993;
srom_1(43185) <= 2586;
srom_1(43186) <= 36503;
srom_1(43187) <= 109586;
srom_1(43188) <= 221493;
srom_1(43189) <= 371698;
srom_1(43190) <= 559497;
srom_1(43191) <= 784009;
srom_1(43192) <= 1044182;
srom_1(43193) <= 1338795;
srom_1(43194) <= 1666467;
srom_1(43195) <= 2025662;
srom_1(43196) <= 2414695;
srom_1(43197) <= 2831741;
srom_1(43198) <= 3274846;
srom_1(43199) <= 3741931;
srom_1(43200) <= 4230805;
srom_1(43201) <= 4739177;
srom_1(43202) <= 5264663;
srom_1(43203) <= 5804797;
srom_1(43204) <= 6357048;
srom_1(43205) <= 6918826;
srom_1(43206) <= 7487496;
srom_1(43207) <= 8060392;
srom_1(43208) <= 8634826;
srom_1(43209) <= 9208106;
srom_1(43210) <= 9777544;
srom_1(43211) <= 10340468;
srom_1(43212) <= 10894239;
srom_1(43213) <= 11436260;
srom_1(43214) <= 11963990;
srom_1(43215) <= 12474953;
srom_1(43216) <= 12966755;
srom_1(43217) <= 13437087;
srom_1(43218) <= 13883746;
srom_1(43219) <= 14304636;
srom_1(43220) <= 14697784;
srom_1(43221) <= 15061346;
srom_1(43222) <= 15393617;
srom_1(43223) <= 15693039;
srom_1(43224) <= 15958209;
srom_1(43225) <= 16187881;
srom_1(43226) <= 16380981;
srom_1(43227) <= 16536601;
srom_1(43228) <= 16654013;
srom_1(43229) <= 16732665;
srom_1(43230) <= 16772189;
srom_1(43231) <= 16772400;
srom_1(43232) <= 16733296;
srom_1(43233) <= 16655061;
srom_1(43234) <= 16538062;
srom_1(43235) <= 16382847;
srom_1(43236) <= 16190144;
srom_1(43237) <= 15960857;
srom_1(43238) <= 15696062;
srom_1(43239) <= 15396999;
srom_1(43240) <= 15065072;
srom_1(43241) <= 14701836;
srom_1(43242) <= 14308995;
srom_1(43243) <= 13888392;
srom_1(43244) <= 13441998;
srom_1(43245) <= 12971907;
srom_1(43246) <= 12480324;
srom_1(43247) <= 11969553;
srom_1(43248) <= 11441990;
srom_1(43249) <= 10900108;
srom_1(43250) <= 10346449;
srom_1(43251) <= 9783609;
srom_1(43252) <= 9214228;
srom_1(43253) <= 8640974;
srom_1(43254) <= 8066538;
srom_1(43255) <= 7493611;
srom_1(43256) <= 6924882;
srom_1(43257) <= 6363017;
srom_1(43258) <= 5810650;
srom_1(43259) <= 5270372;
srom_1(43260) <= 4744716;
srom_1(43261) <= 4236149;
srom_1(43262) <= 3747053;
srom_1(43263) <= 3279723;
srom_1(43264) <= 2836351;
srom_1(43265) <= 2419015;
srom_1(43266) <= 2029672;
srom_1(43267) <= 1670149;
srom_1(43268) <= 1342130;
srom_1(43269) <= 1047155;
srom_1(43270) <= 786607;
srom_1(43271) <= 561707;
srom_1(43272) <= 373510;
srom_1(43273) <= 222899;
srom_1(43274) <= 110580;
srom_1(43275) <= 37079;
srom_1(43276) <= 2741;
srom_1(43277) <= 7727;
srom_1(43278) <= 52014;
srom_1(43279) <= 135395;
srom_1(43280) <= 257477;
srom_1(43281) <= 417689;
srom_1(43282) <= 615280;
srom_1(43283) <= 849322;
srom_1(43284) <= 1118719;
srom_1(43285) <= 1422206;
srom_1(43286) <= 1758362;
srom_1(43287) <= 2125609;
srom_1(43288) <= 2522225;
srom_1(43289) <= 2946351;
srom_1(43290) <= 3395997;
srom_1(43291) <= 3869056;
srom_1(43292) <= 4363308;
srom_1(43293) <= 4876436;
srom_1(43294) <= 5406034;
srom_1(43295) <= 5949618;
srom_1(43296) <= 6504640;
srom_1(43297) <= 7068496;
srom_1(43298) <= 7638542;
srom_1(43299) <= 8212106;
srom_1(43300) <= 8786498;
srom_1(43301) <= 9359023;
srom_1(43302) <= 9926998;
srom_1(43303) <= 10487759;
srom_1(43304) <= 11038677;
srom_1(43305) <= 11577167;
srom_1(43306) <= 12100705;
srom_1(43307) <= 12606836;
srom_1(43308) <= 13093186;
srom_1(43309) <= 13557474;
srom_1(43310) <= 13997524;
srom_1(43311) <= 14411272;
srom_1(43312) <= 14796778;
srom_1(43313) <= 15152233;
srom_1(43314) <= 15475971;
srom_1(43315) <= 15766475;
srom_1(43316) <= 16022381;
srom_1(43317) <= 16242489;
srom_1(43318) <= 16425768;
srom_1(43319) <= 16571358;
srom_1(43320) <= 16678577;
srom_1(43321) <= 16746920;
srom_1(43322) <= 16776069;
srom_1(43323) <= 16765886;
srom_1(43324) <= 16716419;
srom_1(43325) <= 16627900;
srom_1(43326) <= 16500745;
srom_1(43327) <= 16335548;
srom_1(43328) <= 16133086;
srom_1(43329) <= 15894307;
srom_1(43330) <= 15620332;
srom_1(43331) <= 15312444;
srom_1(43332) <= 14972088;
srom_1(43333) <= 14600860;
srom_1(43334) <= 14200500;
srom_1(43335) <= 13772887;
srom_1(43336) <= 13320025;
srom_1(43337) <= 12844037;
srom_1(43338) <= 12347157;
srom_1(43339) <= 11831714;
srom_1(43340) <= 11300124;
srom_1(43341) <= 10754882;
srom_1(43342) <= 10198543;
srom_1(43343) <= 9633717;
srom_1(43344) <= 9063052;
srom_1(43345) <= 8489225;
srom_1(43346) <= 7914925;
srom_1(43347) <= 7342847;
srom_1(43348) <= 6775673;
srom_1(43349) <= 6216062;
srom_1(43350) <= 5666640;
srom_1(43351) <= 5129981;
srom_1(43352) <= 4608603;
srom_1(43353) <= 4104951;
srom_1(43354) <= 3621387;
srom_1(43355) <= 3160177;
srom_1(43356) <= 2723486;
srom_1(43357) <= 2313360;
srom_1(43358) <= 1931723;
srom_1(43359) <= 1580365;
srom_1(43360) <= 1260933;
srom_1(43361) <= 974925;
srom_1(43362) <= 723682;
srom_1(43363) <= 508383;
srom_1(43364) <= 330037;
srom_1(43365) <= 189480;
srom_1(43366) <= 87372;
srom_1(43367) <= 24191;
srom_1(43368) <= 234;
srom_1(43369) <= 15612;
srom_1(43370) <= 70255;
srom_1(43371) <= 163905;
srom_1(43372) <= 296124;
srom_1(43373) <= 466291;
srom_1(43374) <= 673608;
srom_1(43375) <= 917104;
srom_1(43376) <= 1195636;
srom_1(43377) <= 1507899;
srom_1(43378) <= 1852427;
srom_1(43379) <= 2227606;
srom_1(43380) <= 2631676;
srom_1(43381) <= 3062742;
srom_1(43382) <= 3518783;
srom_1(43383) <= 3997660;
srom_1(43384) <= 4497128;
srom_1(43385) <= 5014845;
srom_1(43386) <= 5548382;
srom_1(43387) <= 6095238;
srom_1(43388) <= 6652848;
srom_1(43389) <= 7218598;
srom_1(43390) <= 7789834;
srom_1(43391) <= 8363879;
srom_1(43392) <= 8938039;
srom_1(43393) <= 9509623;
srom_1(43394) <= 10075950;
srom_1(43395) <= 10634364;
srom_1(43396) <= 11182247;
srom_1(43397) <= 11717030;
srom_1(43398) <= 12236205;
srom_1(43399) <= 12737337;
srom_1(43400) <= 13218077;
srom_1(43401) <= 13676169;
srom_1(43402) <= 14109466;
srom_1(43403) <= 14515936;
srom_1(43404) <= 14893673;
srom_1(43405) <= 15240906;
srom_1(43406) <= 15556005;
srom_1(43407) <= 15837495;
srom_1(43408) <= 16084054;
srom_1(43409) <= 16294526;
srom_1(43410) <= 16467925;
srom_1(43411) <= 16603437;
srom_1(43412) <= 16700426;
srom_1(43413) <= 16758439;
srom_1(43414) <= 16777203;
srom_1(43415) <= 16756630;
srom_1(43416) <= 16696816;
srom_1(43417) <= 16598042;
srom_1(43418) <= 16460772;
srom_1(43419) <= 16285648;
srom_1(43420) <= 16073492;
srom_1(43421) <= 15825300;
srom_1(43422) <= 15542234;
srom_1(43423) <= 15225622;
srom_1(43424) <= 14876949;
srom_1(43425) <= 14497850;
srom_1(43426) <= 14090103;
srom_1(43427) <= 13655619;
srom_1(43428) <= 13196437;
srom_1(43429) <= 12714709;
srom_1(43430) <= 12212694;
srom_1(43431) <= 11692747;
srom_1(43432) <= 11157306;
srom_1(43433) <= 10608881;
srom_1(43434) <= 10050045;
srom_1(43435) <= 9483417;
srom_1(43436) <= 8911656;
srom_1(43437) <= 8337442;
srom_1(43438) <= 7763468;
srom_1(43439) <= 7192425;
srom_1(43440) <= 6626992;
srom_1(43441) <= 6069819;
srom_1(43442) <= 5523520;
srom_1(43443) <= 4990657;
srom_1(43444) <= 4473727;
srom_1(43445) <= 3975156;
srom_1(43446) <= 3497281;
srom_1(43447) <= 3042343;
srom_1(43448) <= 2612476;
srom_1(43449) <= 2209695;
srom_1(43450) <= 1835889;
srom_1(43451) <= 1492810;
srom_1(43452) <= 1182069;
srom_1(43453) <= 905122;
srom_1(43454) <= 663267;
srom_1(43455) <= 457639;
srom_1(43456) <= 289201;
srom_1(43457) <= 158745;
srom_1(43458) <= 66882;
srom_1(43459) <= 14042;
srom_1(43460) <= 473;
srom_1(43461) <= 26239;
srom_1(43462) <= 91219;
srom_1(43463) <= 195108;
srom_1(43464) <= 337419;
srom_1(43465) <= 517486;
srom_1(43466) <= 734462;
srom_1(43467) <= 987332;
srom_1(43468) <= 1274908;
srom_1(43469) <= 1595843;
srom_1(43470) <= 1948632;
srom_1(43471) <= 2331620;
srom_1(43472) <= 2743012;
srom_1(43473) <= 3180877;
srom_1(43474) <= 3643163;
srom_1(43475) <= 4127703;
srom_1(43476) <= 4632223;
srom_1(43477) <= 5154358;
srom_1(43478) <= 5691660;
srom_1(43479) <= 6241608;
srom_1(43480) <= 6801625;
srom_1(43481) <= 7369083;
srom_1(43482) <= 7941322;
srom_1(43483) <= 8515659;
srom_1(43484) <= 9089400;
srom_1(43485) <= 9659855;
srom_1(43486) <= 10224348;
srom_1(43487) <= 10780233;
srom_1(43488) <= 11324903;
srom_1(43489) <= 11855804;
srom_1(43490) <= 12370446;
srom_1(43491) <= 12866415;
srom_1(43492) <= 13341386;
srom_1(43493) <= 13793133;
srom_1(43494) <= 14219535;
srom_1(43495) <= 14618594;
srom_1(43496) <= 14988439;
srom_1(43497) <= 15327335;
srom_1(43498) <= 15633693;
srom_1(43499) <= 15906076;
srom_1(43500) <= 16143207;
srom_1(43501) <= 16343974;
srom_1(43502) <= 16507436;
srom_1(43503) <= 16632825;
srom_1(43504) <= 16719555;
srom_1(43505) <= 16767218;
srom_1(43506) <= 16775591;
srom_1(43507) <= 16744634;
srom_1(43508) <= 16674493;
srom_1(43509) <= 16565497;
srom_1(43510) <= 16418156;
srom_1(43511) <= 16233162;
srom_1(43512) <= 16011383;
srom_1(43513) <= 15753857;
srom_1(43514) <= 15461794;
srom_1(43515) <= 15136561;
srom_1(43516) <= 14779686;
srom_1(43517) <= 14392840;
srom_1(43518) <= 13977838;
srom_1(43519) <= 13536627;
srom_1(43520) <= 13071274;
srom_1(43521) <= 12583963;
srom_1(43522) <= 12076979;
srom_1(43523) <= 11552699;
srom_1(43524) <= 11013581;
srom_1(43525) <= 10462153;
srom_1(43526) <= 9901002;
srom_1(43527) <= 9332759;
srom_1(43528) <= 8760089;
srom_1(43529) <= 8185676;
srom_1(43530) <= 7612215;
srom_1(43531) <= 7042395;
srom_1(43532) <= 6478888;
srom_1(43533) <= 5924336;
srom_1(43534) <= 5381339;
srom_1(43535) <= 4852445;
srom_1(43536) <= 4340133;
srom_1(43537) <= 3846806;
srom_1(43538) <= 3374777;
srom_1(43539) <= 2926260;
srom_1(43540) <= 2503357;
srom_1(43541) <= 2108052;
srom_1(43542) <= 1742199;
srom_1(43543) <= 1407513;
srom_1(43544) <= 1105564;
srom_1(43545) <= 837768;
srom_1(43546) <= 605380;
srom_1(43547) <= 409491;
srom_1(43548) <= 251018;
srom_1(43549) <= 130705;
srom_1(43550) <= 49116;
srom_1(43551) <= 6634;
srom_1(43552) <= 3458;
srom_1(43553) <= 39603;
srom_1(43554) <= 114899;
srom_1(43555) <= 228994;
srom_1(43556) <= 381351;
srom_1(43557) <= 571258;
srom_1(43558) <= 797822;
srom_1(43559) <= 1059983;
srom_1(43560) <= 1356509;
srom_1(43561) <= 1686012;
srom_1(43562) <= 2046946;
srom_1(43563) <= 2437618;
srom_1(43564) <= 2856196;
srom_1(43565) <= 3300717;
srom_1(43566) <= 3769097;
srom_1(43567) <= 4259140;
srom_1(43568) <= 4768547;
srom_1(43569) <= 5294930;
srom_1(43570) <= 5835820;
srom_1(43571) <= 6388681;
srom_1(43572) <= 6950921;
srom_1(43573) <= 7519902;
srom_1(43574) <= 8092957;
srom_1(43575) <= 8667398;
srom_1(43576) <= 9240532;
srom_1(43577) <= 9809671;
srom_1(43578) <= 10372146;
srom_1(43579) <= 10925320;
srom_1(43580) <= 11466598;
srom_1(43581) <= 11993442;
srom_1(43582) <= 12503382;
srom_1(43583) <= 12994027;
srom_1(43584) <= 13463075;
srom_1(43585) <= 13908327;
srom_1(43586) <= 14327695;
srom_1(43587) <= 14719213;
srom_1(43588) <= 15081044;
srom_1(43589) <= 15411493;
srom_1(43590) <= 15709008;
srom_1(43591) <= 15972196;
srom_1(43592) <= 16199821;
srom_1(43593) <= 16390818;
srom_1(43594) <= 16544289;
srom_1(43595) <= 16659515;
srom_1(43596) <= 16735956;
srom_1(43597) <= 16773254;
srom_1(43598) <= 16771233;
srom_1(43599) <= 16729903;
srom_1(43600) <= 16649457;
srom_1(43601) <= 16530274;
srom_1(43602) <= 16372912;
srom_1(43603) <= 16178109;
srom_1(43604) <= 15946778;
srom_1(43605) <= 15680004;
srom_1(43606) <= 15379038;
srom_1(43607) <= 15045292;
srom_1(43608) <= 14680330;
srom_1(43609) <= 14285864;
srom_1(43610) <= 13863744;
srom_1(43611) <= 13415949;
srom_1(43612) <= 12944579;
srom_1(43613) <= 12451845;
srom_1(43614) <= 11940057;
srom_1(43615) <= 11411614;
srom_1(43616) <= 10868996;
srom_1(43617) <= 10314747;
srom_1(43618) <= 9751465;
srom_1(43619) <= 9181792;
srom_1(43620) <= 8608400;
srom_1(43621) <= 8033976;
srom_1(43622) <= 7461216;
srom_1(43623) <= 6892805;
srom_1(43624) <= 6331408;
srom_1(43625) <= 5779658;
srom_1(43626) <= 5240143;
srom_1(43627) <= 4715391;
srom_1(43628) <= 4207865;
srom_1(43629) <= 3719943;
srom_1(43630) <= 3253915;
srom_1(43631) <= 2811964;
srom_1(43632) <= 2396165;
srom_1(43633) <= 2008466;
srom_1(43634) <= 1650686;
srom_1(43635) <= 1324502;
srom_1(43636) <= 1031444;
srom_1(43637) <= 772887;
srom_1(43638) <= 550042;
srom_1(43639) <= 363955;
srom_1(43640) <= 215498;
srom_1(43641) <= 105368;
srom_1(43642) <= 34081;
srom_1(43643) <= 1971;
srom_1(43644) <= 9189;
srom_1(43645) <= 55701;
srom_1(43646) <= 141288;
srom_1(43647) <= 265550;
srom_1(43648) <= 427904;
srom_1(43649) <= 627589;
srom_1(43650) <= 863667;
srom_1(43651) <= 1135033;
srom_1(43652) <= 1440413;
srom_1(43653) <= 1778375;
srom_1(43654) <= 2147336;
srom_1(43655) <= 2545563;
srom_1(43656) <= 2971191;
srom_1(43657) <= 3422223;
srom_1(43658) <= 3896543;
srom_1(43659) <= 4391929;
srom_1(43660) <= 4906057;
srom_1(43661) <= 5436515;
srom_1(43662) <= 5980817;
srom_1(43663) <= 6536409;
srom_1(43664) <= 7100688;
srom_1(43665) <= 7671005;
srom_1(43666) <= 8244688;
srom_1(43667) <= 8819046;
srom_1(43668) <= 9391385;
srom_1(43669) <= 9959022;
srom_1(43670) <= 10519295;
srom_1(43671) <= 11069576;
srom_1(43672) <= 11607285;
srom_1(43673) <= 12129900;
srom_1(43674) <= 12634972;
srom_1(43675) <= 13120131;
srom_1(43676) <= 13583102;
srom_1(43677) <= 14021714;
srom_1(43678) <= 14433911;
srom_1(43679) <= 14817759;
srom_1(43680) <= 15171458;
srom_1(43681) <= 15493351;
srom_1(43682) <= 15781927;
srom_1(43683) <= 16035833;
srom_1(43684) <= 16253879;
srom_1(43685) <= 16435041;
srom_1(43686) <= 16578472;
srom_1(43687) <= 16683497;
srom_1(43688) <= 16749624;
srom_1(43689) <= 16776544;
srom_1(43690) <= 16764130;
srom_1(43691) <= 16712440;
srom_1(43692) <= 16621717;
srom_1(43693) <= 16492386;
srom_1(43694) <= 16325054;
srom_1(43695) <= 16120505;
srom_1(43696) <= 15879698;
srom_1(43697) <= 15603763;
srom_1(43698) <= 15293994;
srom_1(43699) <= 14951843;
srom_1(43700) <= 14578914;
srom_1(43701) <= 14176957;
srom_1(43702) <= 13747857;
srom_1(43703) <= 13293625;
srom_1(43704) <= 12816392;
srom_1(43705) <= 12318396;
srom_1(43706) <= 11801971;
srom_1(43707) <= 11269540;
srom_1(43708) <= 10723600;
srom_1(43709) <= 10166709;
srom_1(43710) <= 9601481;
srom_1(43711) <= 9030565;
srom_1(43712) <= 8456638;
srom_1(43713) <= 7882393;
srom_1(43714) <= 7310521;
srom_1(43715) <= 6743705;
srom_1(43716) <= 6184603;
srom_1(43717) <= 5635836;
srom_1(43718) <= 5099977;
srom_1(43719) <= 4579540;
srom_1(43720) <= 4076965;
srom_1(43721) <= 3594609;
srom_1(43722) <= 3134733;
srom_1(43723) <= 2699495;
srom_1(43724) <= 2290935;
srom_1(43725) <= 1910969;
srom_1(43726) <= 1561378;
srom_1(43727) <= 1243803;
srom_1(43728) <= 959733;
srom_1(43729) <= 710499;
srom_1(43730) <= 497270;
srom_1(43731) <= 321047;
srom_1(43732) <= 182655;
srom_1(43733) <= 82743;
srom_1(43734) <= 21781;
srom_1(43735) <= 53;
srom_1(43736) <= 17663;
srom_1(43737) <= 74526;
srom_1(43738) <= 170378;
srom_1(43739) <= 304767;
srom_1(43740) <= 477064;
srom_1(43741) <= 686461;
srom_1(43742) <= 931976;
srom_1(43743) <= 1212458;
srom_1(43744) <= 1526591;
srom_1(43745) <= 1872903;
srom_1(43746) <= 2249769;
srom_1(43747) <= 2655422;
srom_1(43748) <= 3087960;
srom_1(43749) <= 3545354;
srom_1(43750) <= 4025460;
srom_1(43751) <= 4526027;
srom_1(43752) <= 5044706;
srom_1(43753) <= 5579066;
srom_1(43754) <= 6126601;
srom_1(43755) <= 6684744;
srom_1(43756) <= 7250876;
srom_1(43757) <= 7822344;
srom_1(43758) <= 8396466;
srom_1(43759) <= 8970553;
srom_1(43760) <= 9541910;
srom_1(43761) <= 10107859;
srom_1(43762) <= 10665745;
srom_1(43763) <= 11212954;
srom_1(43764) <= 11746918;
srom_1(43765) <= 12265134;
srom_1(43766) <= 12765171;
srom_1(43767) <= 13244686;
srom_1(43768) <= 13701428;
srom_1(43769) <= 14133257;
srom_1(43770) <= 14538147;
srom_1(43771) <= 14914200;
srom_1(43772) <= 15259652;
srom_1(43773) <= 15572883;
srom_1(43774) <= 15852425;
srom_1(43775) <= 16096967;
srom_1(43776) <= 16305361;
srom_1(43777) <= 16476631;
srom_1(43778) <= 16609973;
srom_1(43779) <= 16704763;
srom_1(43780) <= 16760555;
srom_1(43781) <= 16777088;
srom_1(43782) <= 16754285;
srom_1(43783) <= 16692253;
srom_1(43784) <= 16591281;
srom_1(43785) <= 16451845;
srom_1(43786) <= 16274597;
srom_1(43787) <= 16060369;
srom_1(43788) <= 15810166;
srom_1(43789) <= 15525160;
srom_1(43790) <= 15206689;
srom_1(43791) <= 14856245;
srom_1(43792) <= 14475472;
srom_1(43793) <= 14066156;
srom_1(43794) <= 13630216;
srom_1(43795) <= 13169696;
srom_1(43796) <= 12686756;
srom_1(43797) <= 12183660;
srom_1(43798) <= 11662769;
srom_1(43799) <= 11126523;
srom_1(43800) <= 10577439;
srom_1(43801) <= 10018090;
srom_1(43802) <= 9451100;
srom_1(43803) <= 8879128;
srom_1(43804) <= 8304855;
srom_1(43805) <= 7730975;
srom_1(43806) <= 7160179;
srom_1(43807) <= 6595144;
srom_1(43808) <= 6038519;
srom_1(43809) <= 5492914;
srom_1(43810) <= 4960888;
srom_1(43811) <= 4444936;
srom_1(43812) <= 3947477;
srom_1(43813) <= 3470844;
srom_1(43814) <= 3017272;
srom_1(43815) <= 2588888;
srom_1(43816) <= 2187701;
srom_1(43817) <= 1815592;
srom_1(43818) <= 1474306;
srom_1(43819) <= 1165444;
srom_1(43820) <= 890454;
srom_1(43821) <= 650625;
srom_1(43822) <= 447082;
srom_1(43823) <= 280780;
srom_1(43824) <= 152498;
srom_1(43825) <= 62838;
srom_1(43826) <= 12220;
srom_1(43827) <= 882;
srom_1(43828) <= 28877;
srom_1(43829) <= 96074;
srom_1(43830) <= 202157;
srom_1(43831) <= 346630;
srom_1(43832) <= 528814;
srom_1(43833) <= 747855;
srom_1(43834) <= 1002726;
srom_1(43835) <= 1292232;
srom_1(43836) <= 1615016;
srom_1(43837) <= 1969563;
srom_1(43838) <= 2354212;
srom_1(43839) <= 2767157;
srom_1(43840) <= 3206464;
srom_1(43841) <= 3670071;
srom_1(43842) <= 4155806;
srom_1(43843) <= 4661389;
srom_1(43844) <= 5184451;
srom_1(43845) <= 5722538;
srom_1(43846) <= 6273127;
srom_1(43847) <= 6833636;
srom_1(43848) <= 7401437;
srom_1(43849) <= 7973867;
srom_1(43850) <= 8548242;
srom_1(43851) <= 9121869;
srom_1(43852) <= 9692057;
srom_1(43853) <= 10256132;
srom_1(43854) <= 10811451;
srom_1(43855) <= 11355407;
srom_1(43856) <= 11885452;
srom_1(43857) <= 12399098;
srom_1(43858) <= 12893938;
srom_1(43859) <= 13367651;
srom_1(43860) <= 13818015;
srom_1(43861) <= 14242919;
srom_1(43862) <= 14640370;
srom_1(43863) <= 15008504;
srom_1(43864) <= 15345596;
srom_1(43865) <= 15650064;
srom_1(43866) <= 15920480;
srom_1(43867) <= 16155577;
srom_1(43868) <= 16354251;
srom_1(43869) <= 16515572;
srom_1(43870) <= 16638783;
srom_1(43871) <= 16723306;
srom_1(43872) <= 16768745;
srom_1(43873) <= 16774886;
srom_1(43874) <= 16741702;
srom_1(43875) <= 16669346;
srom_1(43876) <= 16558160;
srom_1(43877) <= 16408664;
srom_1(43878) <= 16221558;
srom_1(43879) <= 15997722;
srom_1(43880) <= 15738204;
srom_1(43881) <= 15444221;
srom_1(43882) <= 15117151;
srom_1(43883) <= 14758530;
srom_1(43884) <= 14370037;
srom_1(43885) <= 13953496;
srom_1(43886) <= 13510858;
srom_1(43887) <= 13044201;
srom_1(43888) <= 12555712;
srom_1(43889) <= 12047682;
srom_1(43890) <= 11522494;
srom_1(43891) <= 10982610;
srom_1(43892) <= 10430561;
srom_1(43893) <= 9868937;
srom_1(43894) <= 9300371;
srom_1(43895) <= 8727530;
srom_1(43896) <= 8153099;
srom_1(43897) <= 7579773;
srom_1(43898) <= 7010240;
srom_1(43899) <= 6447170;
srom_1(43900) <= 5893204;
srom_1(43901) <= 5350940;
srom_1(43902) <= 4822921;
srom_1(43903) <= 4311623;
srom_1(43904) <= 3819442;
srom_1(43905) <= 3348689;
srom_1(43906) <= 2901569;
srom_1(43907) <= 2480180;
srom_1(43908) <= 2086497;
srom_1(43909) <= 1722367;
srom_1(43910) <= 1389498;
srom_1(43911) <= 1089449;
srom_1(43912) <= 823629;
srom_1(43913) <= 593284;
srom_1(43914) <= 399494;
srom_1(43915) <= 243167;
srom_1(43916) <= 125037;
srom_1(43917) <= 45658;
srom_1(43918) <= 5402;
srom_1(43919) <= 4457;
srom_1(43920) <= 42829;
srom_1(43921) <= 120337;
srom_1(43922) <= 236617;
srom_1(43923) <= 391125;
srom_1(43924) <= 583137;
srom_1(43925) <= 811750;
srom_1(43926) <= 1075894;
srom_1(43927) <= 1374330;
srom_1(43928) <= 1705658;
srom_1(43929) <= 2068325;
srom_1(43930) <= 2460630;
srom_1(43931) <= 2880733;
srom_1(43932) <= 3326665;
srom_1(43933) <= 3796333;
srom_1(43934) <= 4287537;
srom_1(43935) <= 4797972;
srom_1(43936) <= 5325244;
srom_1(43937) <= 5866882;
srom_1(43938) <= 6420344;
srom_1(43939) <= 6983037;
srom_1(43940) <= 7552321;
srom_1(43941) <= 8125527;
srom_1(43942) <= 8699966;
srom_1(43943) <= 9272945;
srom_1(43944) <= 9841777;
srom_1(43945) <= 10403795;
srom_1(43946) <= 10956363;
srom_1(43947) <= 11496889;
srom_1(43948) <= 12022840;
srom_1(43949) <= 12531749;
srom_1(43950) <= 13021229;
srom_1(43951) <= 13488986;
srom_1(43952) <= 13932824;
srom_1(43953) <= 14350664;
srom_1(43954) <= 14740546;
srom_1(43955) <= 15100642;
srom_1(43956) <= 15429262;
srom_1(43957) <= 15724866;
srom_1(43958) <= 15986069;
srom_1(43959) <= 16211644;
srom_1(43960) <= 16400534;
srom_1(43961) <= 16551853;
srom_1(43962) <= 16664892;
srom_1(43963) <= 16739121;
srom_1(43964) <= 16774191;
srom_1(43965) <= 16769939;
srom_1(43966) <= 16726383;
srom_1(43967) <= 16643729;
srom_1(43968) <= 16522364;
srom_1(43969) <= 16362857;
srom_1(43970) <= 16165956;
srom_1(43971) <= 15932584;
srom_1(43972) <= 15663835;
srom_1(43973) <= 15360971;
srom_1(43974) <= 15025411;
srom_1(43975) <= 14658729;
srom_1(43976) <= 14262644;
srom_1(43977) <= 13839013;
srom_1(43978) <= 13389824;
srom_1(43979) <= 12917182;
srom_1(43980) <= 12423304;
srom_1(43981) <= 11910507;
srom_1(43982) <= 11381193;
srom_1(43983) <= 10837847;
srom_1(43984) <= 10283015;
srom_1(43985) <= 9719300;
srom_1(43986) <= 9149344;
srom_1(43987) <= 8575821;
srom_1(43988) <= 8001421;
srom_1(43989) <= 7428835;
srom_1(43990) <= 6860751;
srom_1(43991) <= 6299831;
srom_1(43992) <= 5748707;
srom_1(43993) <= 5209961;
srom_1(43994) <= 4686122;
srom_1(43995) <= 4179644;
srom_1(43996) <= 3692904;
srom_1(43997) <= 3228184;
srom_1(43998) <= 2787662;
srom_1(43999) <= 2373406;
srom_1(44000) <= 1987356;
srom_1(44001) <= 1631325;
srom_1(44002) <= 1306981;
srom_1(44003) <= 1015844;
srom_1(44004) <= 759281;
srom_1(44005) <= 538495;
srom_1(44006) <= 354521;
srom_1(44007) <= 208221;
srom_1(44008) <= 100282;
srom_1(44009) <= 31209;
srom_1(44010) <= 1328;
srom_1(44011) <= 10777;
srom_1(44012) <= 59513;
srom_1(44013) <= 147306;
srom_1(44014) <= 273746;
srom_1(44015) <= 438240;
srom_1(44016) <= 640015;
srom_1(44017) <= 878126;
srom_1(44018) <= 1151456;
srom_1(44019) <= 1458724;
srom_1(44020) <= 1798489;
srom_1(44021) <= 2169156;
srom_1(44022) <= 2568989;
srom_1(44023) <= 2996112;
srom_1(44024) <= 3448523;
srom_1(44025) <= 3924099;
srom_1(44026) <= 4420611;
srom_1(44027) <= 4935730;
srom_1(44028) <= 5467040;
srom_1(44029) <= 6012051;
srom_1(44030) <= 6568207;
srom_1(44031) <= 7132899;
srom_1(44032) <= 7703479;
srom_1(44033) <= 8277272;
srom_1(44034) <= 8851587;
srom_1(44035) <= 9423732;
srom_1(44036) <= 9991022;
srom_1(44037) <= 10550798;
srom_1(44038) <= 11100434;
srom_1(44039) <= 11637354;
srom_1(44040) <= 12159039;
srom_1(44041) <= 12663044;
srom_1(44042) <= 13147004;
srom_1(44043) <= 13608651;
srom_1(44044) <= 14045819;
srom_1(44045) <= 14456458;
srom_1(44046) <= 14838643;
srom_1(44047) <= 15190581;
srom_1(44048) <= 15510623;
srom_1(44049) <= 15797268;
srom_1(44050) <= 16049170;
srom_1(44051) <= 16265149;
srom_1(44052) <= 16444193;
srom_1(44053) <= 16585461;
srom_1(44054) <= 16688292;
srom_1(44055) <= 16752202;
srom_1(44056) <= 16776892;
srom_1(44057) <= 16762247;
srom_1(44058) <= 16708335;
srom_1(44059) <= 16615409;
srom_1(44060) <= 16483905;
srom_1(44061) <= 16314439;
srom_1(44062) <= 16107806;
srom_1(44063) <= 15864976;
srom_1(44064) <= 15587085;
srom_1(44065) <= 15275439;
srom_1(44066) <= 14931498;
srom_1(44067) <= 14556875;
srom_1(44068) <= 14153327;
srom_1(44069) <= 13722747;
srom_1(44070) <= 13267152;
srom_1(44071) <= 12788681;
srom_1(44072) <= 12289576;
srom_1(44073) <= 11772178;
srom_1(44074) <= 11238913;
srom_1(44075) <= 10692282;
srom_1(44076) <= 10134849;
srom_1(44077) <= 9569226;
srom_1(44078) <= 8998068;
srom_1(44079) <= 8424051;
srom_1(44080) <= 7849869;
srom_1(44081) <= 7278212;
srom_1(44082) <= 6711763;
srom_1(44083) <= 6153177;
srom_1(44084) <= 5605073;
srom_1(44085) <= 5070023;
srom_1(44086) <= 4550534;
srom_1(44087) <= 4049044;
srom_1(44088) <= 3567903;
srom_1(44089) <= 3109368;
srom_1(44090) <= 2675590;
srom_1(44091) <= 2268601;
srom_1(44092) <= 1890312;
srom_1(44093) <= 1542495;
srom_1(44094) <= 1226782;
srom_1(44095) <= 944653;
srom_1(44096) <= 697432;
srom_1(44097) <= 486277;
srom_1(44098) <= 312178;
srom_1(44099) <= 175953;
srom_1(44100) <= 78240;
srom_1(44101) <= 19497;
srom_1(44102) <= 0;
srom_1(44103) <= 19840;
srom_1(44104) <= 78923;
srom_1(44105) <= 176974;
srom_1(44106) <= 313532;
srom_1(44107) <= 487957;
srom_1(44108) <= 699430;
srom_1(44109) <= 946961;
srom_1(44110) <= 1229388;
srom_1(44111) <= 1545387;
srom_1(44112) <= 1893477;
srom_1(44113) <= 2272024;
srom_1(44114) <= 2679254;
srom_1(44115) <= 3113257;
srom_1(44116) <= 3571998;
srom_1(44117) <= 4053326;
srom_1(44118) <= 4554983;
srom_1(44119) <= 5074618;
srom_1(44120) <= 5609793;
srom_1(44121) <= 6157999;
srom_1(44122) <= 6716665;
srom_1(44123) <= 7283171;
srom_1(44124) <= 7854861;
srom_1(44125) <= 8429054;
srom_1(44126) <= 9003057;
srom_1(44127) <= 9574179;
srom_1(44128) <= 10139742;
srom_1(44129) <= 10697092;
srom_1(44130) <= 11243618;
srom_1(44131) <= 11776755;
srom_1(44132) <= 12294004;
srom_1(44133) <= 12792939;
srom_1(44134) <= 13271221;
srom_1(44135) <= 13726607;
srom_1(44136) <= 14156961;
srom_1(44137) <= 14560265;
srom_1(44138) <= 14934628;
srom_1(44139) <= 15278294;
srom_1(44140) <= 15589653;
srom_1(44141) <= 15867243;
srom_1(44142) <= 16109763;
srom_1(44143) <= 16316077;
srom_1(44144) <= 16485215;
srom_1(44145) <= 16616386;
srom_1(44146) <= 16708974;
srom_1(44147) <= 16762545;
srom_1(44148) <= 16776847;
srom_1(44149) <= 16751814;
srom_1(44150) <= 16687564;
srom_1(44151) <= 16584396;
srom_1(44152) <= 16442796;
srom_1(44153) <= 16263427;
srom_1(44154) <= 16047130;
srom_1(44155) <= 15794920;
srom_1(44156) <= 15507979;
srom_1(44157) <= 15187652;
srom_1(44158) <= 14835443;
srom_1(44159) <= 14453002;
srom_1(44160) <= 14042124;
srom_1(44161) <= 13604733;
srom_1(44162) <= 13142883;
srom_1(44163) <= 12658738;
srom_1(44164) <= 12154570;
srom_1(44165) <= 11632741;
srom_1(44166) <= 11095699;
srom_1(44167) <= 10545963;
srom_1(44168) <= 9986111;
srom_1(44169) <= 9418767;
srom_1(44170) <= 8846592;
srom_1(44171) <= 8272270;
srom_1(44172) <= 7698493;
srom_1(44173) <= 7127952;
srom_1(44174) <= 6563323;
srom_1(44175) <= 6007254;
srom_1(44176) <= 5462351;
srom_1(44177) <= 4931171;
srom_1(44178) <= 4416203;
srom_1(44179) <= 3919864;
srom_1(44180) <= 3444480;
srom_1(44181) <= 2992281;
srom_1(44182) <= 2565387;
srom_1(44183) <= 2165800;
srom_1(44184) <= 1795394;
srom_1(44185) <= 1455906;
srom_1(44186) <= 1148928;
srom_1(44187) <= 875899;
srom_1(44188) <= 638100;
srom_1(44189) <= 436645;
srom_1(44190) <= 272480;
srom_1(44191) <= 146374;
srom_1(44192) <= 58919;
srom_1(44193) <= 10525;
srom_1(44194) <= 1418;
srom_1(44195) <= 31642;
srom_1(44196) <= 101055;
srom_1(44197) <= 209330;
srom_1(44198) <= 355961;
srom_1(44199) <= 540260;
srom_1(44200) <= 761363;
srom_1(44201) <= 1018232;
srom_1(44202) <= 1309663;
srom_1(44203) <= 1634291;
srom_1(44204) <= 1990591;
srom_1(44205) <= 2376894;
srom_1(44206) <= 2791388;
srom_1(44207) <= 3232129;
srom_1(44208) <= 3697051;
srom_1(44209) <= 4183973;
srom_1(44210) <= 4690611;
srom_1(44211) <= 5214592;
srom_1(44212) <= 5753456;
srom_1(44213) <= 6304677;
srom_1(44214) <= 6865671;
srom_1(44215) <= 7433806;
srom_1(44216) <= 8006418;
srom_1(44217) <= 8580823;
srom_1(44218) <= 9154326;
srom_1(44219) <= 9724239;
srom_1(44220) <= 10287888;
srom_1(44221) <= 10842631;
srom_1(44222) <= 11385867;
srom_1(44223) <= 11915047;
srom_1(44224) <= 12427690;
srom_1(44225) <= 12921393;
srom_1(44226) <= 13393840;
srom_1(44227) <= 13842815;
srom_1(44228) <= 14266214;
srom_1(44229) <= 14662051;
srom_1(44230) <= 15028470;
srom_1(44231) <= 15363752;
srom_1(44232) <= 15666325;
srom_1(44233) <= 15934770;
srom_1(44234) <= 16167829;
srom_1(44235) <= 16364408;
srom_1(44236) <= 16523586;
srom_1(44237) <= 16644617;
srom_1(44238) <= 16726932;
srom_1(44239) <= 16770146;
srom_1(44240) <= 16774056;
srom_1(44241) <= 16738643;
srom_1(44242) <= 16664075;
srom_1(44243) <= 16550700;
srom_1(44244) <= 16399050;
srom_1(44245) <= 16209836;
srom_1(44246) <= 15983946;
srom_1(44247) <= 15722439;
srom_1(44248) <= 15426541;
srom_1(44249) <= 15097640;
srom_1(44250) <= 14737277;
srom_1(44251) <= 14347144;
srom_1(44252) <= 13929069;
srom_1(44253) <= 13485013;
srom_1(44254) <= 13017058;
srom_1(44255) <= 12527398;
srom_1(44256) <= 12018331;
srom_1(44257) <= 11492242;
srom_1(44258) <= 10951599;
srom_1(44259) <= 10398938;
srom_1(44260) <= 9836850;
srom_1(44261) <= 9267970;
srom_1(44262) <= 8694966;
srom_1(44263) <= 8120526;
srom_1(44264) <= 7547343;
srom_1(44265) <= 6978105;
srom_1(44266) <= 6415482;
srom_1(44267) <= 5862111;
srom_1(44268) <= 5320587;
srom_1(44269) <= 4793451;
srom_1(44270) <= 4283173;
srom_1(44271) <= 3792148;
srom_1(44272) <= 3322676;
srom_1(44273) <= 2876961;
srom_1(44274) <= 2457091;
srom_1(44275) <= 2065037;
srom_1(44276) <= 1702636;
srom_1(44277) <= 1371587;
srom_1(44278) <= 1073444;
srom_1(44279) <= 809604;
srom_1(44280) <= 581305;
srom_1(44281) <= 389617;
srom_1(44282) <= 235439;
srom_1(44283) <= 119494;
srom_1(44284) <= 42325;
srom_1(44285) <= 4296;
srom_1(44286) <= 5583;
srom_1(44287) <= 46181;
srom_1(44288) <= 125899;
srom_1(44289) <= 244364;
srom_1(44290) <= 401021;
srom_1(44291) <= 595133;
srom_1(44292) <= 825792;
srom_1(44293) <= 1091916;
srom_1(44294) <= 1392257;
srom_1(44295) <= 1725405;
srom_1(44296) <= 2089800;
srom_1(44297) <= 2483732;
srom_1(44298) <= 2905354;
srom_1(44299) <= 3352689;
srom_1(44300) <= 3823639;
srom_1(44301) <= 4315996;
srom_1(44302) <= 4827450;
srom_1(44303) <= 5355604;
srom_1(44304) <= 5897981;
srom_1(44305) <= 6452037;
srom_1(44306) <= 7015175;
srom_1(44307) <= 7584753;
srom_1(44308) <= 8158100;
srom_1(44309) <= 8732529;
srom_1(44310) <= 9305344;
srom_1(44311) <= 9873861;
srom_1(44312) <= 10435413;
srom_1(44313) <= 10987367;
srom_1(44314) <= 11527134;
srom_1(44315) <= 12052184;
srom_1(44316) <= 12560054;
srom_1(44317) <= 13048362;
srom_1(44318) <= 13514819;
srom_1(44319) <= 13957238;
srom_1(44320) <= 14373544;
srom_1(44321) <= 14761784;
srom_1(44322) <= 15120138;
srom_1(44323) <= 15446925;
srom_1(44324) <= 15740614;
srom_1(44325) <= 15999827;
srom_1(44326) <= 16223348;
srom_1(44327) <= 16410129;
srom_1(44328) <= 16559294;
srom_1(44329) <= 16670145;
srom_1(44330) <= 16742160;
srom_1(44331) <= 16775003;
srom_1(44332) <= 16768519;
srom_1(44333) <= 16722739;
srom_1(44334) <= 16637877;
srom_1(44335) <= 16514331;
srom_1(44336) <= 16352681;
srom_1(44337) <= 16153685;
srom_1(44338) <= 15918276;
srom_1(44339) <= 15647557;
srom_1(44340) <= 15342799;
srom_1(44341) <= 15005430;
srom_1(44342) <= 14637033;
srom_1(44343) <= 14239335;
srom_1(44344) <= 13814200;
srom_1(44345) <= 13363623;
srom_1(44346) <= 12889717;
srom_1(44347) <= 12394703;
srom_1(44348) <= 11880903;
srom_1(44349) <= 11350727;
srom_1(44350) <= 10806661;
srom_1(44351) <= 10251255;
srom_1(44352) <= 9687114;
srom_1(44353) <= 9116885;
srom_1(44354) <= 8543240;
srom_1(44355) <= 7968870;
srom_1(44356) <= 7396469;
srom_1(44357) <= 6828720;
srom_1(44358) <= 6268286;
srom_1(44359) <= 5717794;
srom_1(44360) <= 5179828;
srom_1(44361) <= 4656908;
srom_1(44362) <= 4151487;
srom_1(44363) <= 3665936;
srom_1(44364) <= 3202531;
srom_1(44365) <= 2763445;
srom_1(44366) <= 2350737;
srom_1(44367) <= 1966344;
srom_1(44368) <= 1612066;
srom_1(44369) <= 1289566;
srom_1(44370) <= 1000355;
srom_1(44371) <= 745791;
srom_1(44372) <= 527067;
srom_1(44373) <= 345208;
srom_1(44374) <= 201067;
srom_1(44375) <= 95321;
srom_1(44376) <= 28464;
srom_1(44377) <= 811;
srom_1(44378) <= 12492;
srom_1(44379) <= 63450;
srom_1(44380) <= 153449;
srom_1(44381) <= 282065;
srom_1(44382) <= 448695;
srom_1(44383) <= 652558;
srom_1(44384) <= 892698;
srom_1(44385) <= 1167989;
srom_1(44386) <= 1477140;
srom_1(44387) <= 1818701;
srom_1(44388) <= 2191071;
srom_1(44389) <= 2592503;
srom_1(44390) <= 3021115;
srom_1(44391) <= 3474898;
srom_1(44392) <= 3951722;
srom_1(44393) <= 4449352;
srom_1(44394) <= 4965455;
srom_1(44395) <= 5497610;
srom_1(44396) <= 6043322;
srom_1(44397) <= 6600032;
srom_1(44398) <= 7165129;
srom_1(44399) <= 7735963;
srom_1(44400) <= 8309858;
srom_1(44401) <= 8884122;
srom_1(44402) <= 9456062;
srom_1(44403) <= 10022997;
srom_1(44404) <= 10582268;
srom_1(44405) <= 11131252;
srom_1(44406) <= 11667374;
srom_1(44407) <= 12188121;
srom_1(44408) <= 12691051;
srom_1(44409) <= 13173806;
srom_1(44410) <= 13634121;
srom_1(44411) <= 14069838;
srom_1(44412) <= 14478913;
srom_1(44413) <= 14859430;
srom_1(44414) <= 15209602;
srom_1(44415) <= 15527788;
srom_1(44416) <= 15812496;
srom_1(44417) <= 16062391;
srom_1(44418) <= 16276301;
srom_1(44419) <= 16453223;
srom_1(44420) <= 16592327;
srom_1(44421) <= 16692961;
srom_1(44422) <= 16754653;
srom_1(44423) <= 16777114;
srom_1(44424) <= 16760238;
srom_1(44425) <= 16704105;
srom_1(44426) <= 16608978;
srom_1(44427) <= 16475302;
srom_1(44428) <= 16303705;
srom_1(44429) <= 16094992;
srom_1(44430) <= 15850140;
srom_1(44431) <= 15570299;
srom_1(44432) <= 15256781;
srom_1(44433) <= 14911055;
srom_1(44434) <= 14534743;
srom_1(44435) <= 14129610;
srom_1(44436) <= 13697555;
srom_1(44437) <= 13240605;
srom_1(44438) <= 12760902;
srom_1(44439) <= 12260696;
srom_1(44440) <= 11742333;
srom_1(44441) <= 11208243;
srom_1(44442) <= 10660930;
srom_1(44443) <= 10102962;
srom_1(44444) <= 9536954;
srom_1(44445) <= 8965562;
srom_1(44446) <= 8391464;
srom_1(44447) <= 7817352;
srom_1(44448) <= 7245920;
srom_1(44449) <= 6679845;
srom_1(44450) <= 6121784;
srom_1(44451) <= 5574353;
srom_1(44452) <= 5040119;
srom_1(44453) <= 4521586;
srom_1(44454) <= 4021188;
srom_1(44455) <= 3541270;
srom_1(44456) <= 3084083;
srom_1(44457) <= 2651771;
srom_1(44458) <= 2246360;
srom_1(44459) <= 1869753;
srom_1(44460) <= 1523715;
srom_1(44461) <= 1209868;
srom_1(44462) <= 929686;
srom_1(44463) <= 684480;
srom_1(44464) <= 475402;
srom_1(44465) <= 303432;
srom_1(44466) <= 169376;
srom_1(44467) <= 73862;
srom_1(44468) <= 17340;
srom_1(44469) <= 73;
srom_1(44470) <= 22143;
srom_1(44471) <= 83446;
srom_1(44472) <= 183695;
srom_1(44473) <= 322419;
srom_1(44474) <= 498969;
srom_1(44475) <= 712515;
srom_1(44476) <= 962058;
srom_1(44477) <= 1246426;
srom_1(44478) <= 1564287;
srom_1(44479) <= 1914149;
srom_1(44480) <= 2294371;
srom_1(44481) <= 2703172;
srom_1(44482) <= 3138634;
srom_1(44483) <= 3598715;
srom_1(44484) <= 4081257;
srom_1(44485) <= 4583998;
srom_1(44486) <= 5104580;
srom_1(44487) <= 5640562;
srom_1(44488) <= 6189430;
srom_1(44489) <= 6748611;
srom_1(44490) <= 7315483;
srom_1(44491) <= 7887387;
srom_1(44492) <= 8461641;
srom_1(44493) <= 9035553;
srom_1(44494) <= 9606431;
srom_1(44495) <= 10171598;
srom_1(44496) <= 10728404;
srom_1(44497) <= 11274238;
srom_1(44498) <= 11806541;
srom_1(44499) <= 12322815;
srom_1(44500) <= 12820641;
srom_1(44501) <= 13297683;
srom_1(44502) <= 13751705;
srom_1(44503) <= 14180577;
srom_1(44504) <= 14582289;
srom_1(44505) <= 14954957;
srom_1(44506) <= 15296833;
srom_1(44507) <= 15606314;
srom_1(44508) <= 15881948;
srom_1(44509) <= 16122444;
srom_1(44510) <= 16326673;
srom_1(44511) <= 16493677;
srom_1(44512) <= 16622674;
srom_1(44513) <= 16713059;
srom_1(44514) <= 16764408;
srom_1(44515) <= 16776479;
srom_1(44516) <= 16749217;
srom_1(44517) <= 16682749;
srom_1(44518) <= 16577388;
srom_1(44519) <= 16433626;
srom_1(44520) <= 16252138;
srom_1(44521) <= 16033775;
srom_1(44522) <= 15779562;
srom_1(44523) <= 15490690;
srom_1(44524) <= 15168514;
srom_1(44525) <= 14814544;
srom_1(44526) <= 14430441;
srom_1(44527) <= 14018006;
srom_1(44528) <= 13579172;
srom_1(44529) <= 13115999;
srom_1(44530) <= 12630657;
srom_1(44531) <= 12125422;
srom_1(44532) <= 11602664;
srom_1(44533) <= 11064835;
srom_1(44534) <= 10514455;
srom_1(44535) <= 9954107;
srom_1(44536) <= 9386418;
srom_1(44537) <= 8814049;
srom_1(44538) <= 8239686;
srom_1(44539) <= 7666021;
srom_1(44540) <= 7095744;
srom_1(44541) <= 6531530;
srom_1(44542) <= 5976025;
srom_1(44543) <= 5431833;
srom_1(44544) <= 4901506;
srom_1(44545) <= 4387531;
srom_1(44546) <= 3892319;
srom_1(44547) <= 3418192;
srom_1(44548) <= 2967372;
srom_1(44549) <= 2541975;
srom_1(44550) <= 2143994;
srom_1(44551) <= 1775296;
srom_1(44552) <= 1437611;
srom_1(44553) <= 1132521;
srom_1(44554) <= 861458;
srom_1(44555) <= 625692;
srom_1(44556) <= 426328;
srom_1(44557) <= 264303;
srom_1(44558) <= 140375;
srom_1(44559) <= 55127;
srom_1(44560) <= 8956;
srom_1(44561) <= 2081;
srom_1(44562) <= 34533;
srom_1(44563) <= 106160;
srom_1(44564) <= 216627;
srom_1(44565) <= 365414;
srom_1(44566) <= 551825;
srom_1(44567) <= 774986;
srom_1(44568) <= 1033849;
srom_1(44569) <= 1327201;
srom_1(44570) <= 1653667;
srom_1(44571) <= 2011715;
srom_1(44572) <= 2399667;
srom_1(44573) <= 2815703;
srom_1(44574) <= 3257872;
srom_1(44575) <= 3724101;
srom_1(44576) <= 4212203;
srom_1(44577) <= 4719890;
srom_1(44578) <= 5244781;
srom_1(44579) <= 5784414;
srom_1(44580) <= 6336259;
srom_1(44581) <= 6897728;
srom_1(44582) <= 7466189;
srom_1(44583) <= 8038975;
srom_1(44584) <= 8613401;
srom_1(44585) <= 9186772;
srom_1(44586) <= 9756401;
srom_1(44587) <= 10319615;
srom_1(44588) <= 10873775;
srom_1(44589) <= 11416281;
srom_1(44590) <= 11944588;
srom_1(44591) <= 12456221;
srom_1(44592) <= 12948779;
srom_1(44593) <= 13419953;
srom_1(44594) <= 13867533;
srom_1(44595) <= 14289421;
srom_1(44596) <= 14683638;
srom_1(44597) <= 15048335;
srom_1(44598) <= 15381802;
srom_1(44599) <= 15682476;
srom_1(44600) <= 15948947;
srom_1(44601) <= 16179964;
srom_1(44602) <= 16374445;
srom_1(44603) <= 16531478;
srom_1(44604) <= 16650326;
srom_1(44605) <= 16730432;
srom_1(44606) <= 16771420;
srom_1(44607) <= 16773098;
srom_1(44608) <= 16735459;
srom_1(44609) <= 16658678;
srom_1(44610) <= 16543116;
srom_1(44611) <= 16389315;
srom_1(44612) <= 16197996;
srom_1(44613) <= 15970056;
srom_1(44614) <= 15706564;
srom_1(44615) <= 15408755;
srom_1(44616) <= 15078027;
srom_1(44617) <= 14715929;
srom_1(44618) <= 14324161;
srom_1(44619) <= 13904559;
srom_1(44620) <= 13459090;
srom_1(44621) <= 12989844;
srom_1(44622) <= 12499022;
srom_1(44623) <= 11988924;
srom_1(44624) <= 11461943;
srom_1(44625) <= 10920551;
srom_1(44626) <= 10367285;
srom_1(44627) <= 9804740;
srom_1(44628) <= 9235555;
srom_1(44629) <= 8662398;
srom_1(44630) <= 8087957;
srom_1(44631) <= 7514926;
srom_1(44632) <= 6945992;
srom_1(44633) <= 6383823;
srom_1(44634) <= 5831055;
srom_1(44635) <= 5290280;
srom_1(44636) <= 4764035;
srom_1(44637) <= 4254786;
srom_1(44638) <= 3764922;
srom_1(44639) <= 3296740;
srom_1(44640) <= 2852436;
srom_1(44641) <= 2434093;
srom_1(44642) <= 2043672;
srom_1(44643) <= 1683005;
srom_1(44644) <= 1353783;
srom_1(44645) <= 1057550;
srom_1(44646) <= 795694;
srom_1(44647) <= 569444;
srom_1(44648) <= 379861;
srom_1(44649) <= 227834;
srom_1(44650) <= 114075;
srom_1(44651) <= 39119;
srom_1(44652) <= 3316;
srom_1(44653) <= 6835;
srom_1(44654) <= 49658;
srom_1(44655) <= 131586;
srom_1(44656) <= 252234;
srom_1(44657) <= 411036;
srom_1(44658) <= 607248;
srom_1(44659) <= 839949;
srom_1(44660) <= 1108048;
srom_1(44661) <= 1410289;
srom_1(44662) <= 1745253;
srom_1(44663) <= 2111370;
srom_1(44664) <= 2506923;
srom_1(44665) <= 2930058;
srom_1(44666) <= 3378789;
srom_1(44667) <= 3851013;
srom_1(44668) <= 4344516;
srom_1(44669) <= 4856983;
srom_1(44670) <= 5386010;
srom_1(44671) <= 5929118;
srom_1(44672) <= 6483759;
srom_1(44673) <= 7047333;
srom_1(44674) <= 7617197;
srom_1(44675) <= 8190677;
srom_1(44676) <= 8765087;
srom_1(44677) <= 9337730;
srom_1(44678) <= 9905923;
srom_1(44679) <= 10467000;
srom_1(44680) <= 11018332;
srom_1(44681) <= 11557331;
srom_1(44682) <= 12081472;
srom_1(44683) <= 12588295;
srom_1(44684) <= 13075424;
srom_1(44685) <= 13540576;
srom_1(44686) <= 13981568;
srom_1(44687) <= 14396333;
srom_1(44688) <= 14782925;
srom_1(44689) <= 15139532;
srom_1(44690) <= 15464482;
srom_1(44691) <= 15756251;
srom_1(44692) <= 16013470;
srom_1(44693) <= 16234933;
srom_1(44694) <= 16419603;
srom_1(44695) <= 16566612;
srom_1(44696) <= 16675272;
srom_1(44697) <= 16745073;
srom_1(44698) <= 16775688;
srom_1(44699) <= 16766972;
srom_1(44700) <= 16718968;
srom_1(44701) <= 16631900;
srom_1(44702) <= 16506176;
srom_1(44703) <= 16342386;
srom_1(44704) <= 16141298;
srom_1(44705) <= 15903854;
srom_1(44706) <= 15631170;
srom_1(44707) <= 15324522;
srom_1(44708) <= 14985350;
srom_1(44709) <= 14615243;
srom_1(44710) <= 14215937;
srom_1(44711) <= 13789305;
srom_1(44712) <= 13337348;
srom_1(44713) <= 12862184;
srom_1(44714) <= 12366041;
srom_1(44715) <= 11851248;
srom_1(44716) <= 11320216;
srom_1(44717) <= 10775438;
srom_1(44718) <= 10219466;
srom_1(44719) <= 9654910;
srom_1(44720) <= 9084415;
srom_1(44721) <= 8510657;
srom_1(44722) <= 7936327;
srom_1(44723) <= 7364117;
srom_1(44724) <= 6796712;
srom_1(44725) <= 6236772;
srom_1(44726) <= 5686923;
srom_1(44727) <= 5149742;
srom_1(44728) <= 4627750;
srom_1(44729) <= 4123394;
srom_1(44730) <= 3639039;
srom_1(44731) <= 3176956;
srom_1(44732) <= 2739312;
srom_1(44733) <= 2328160;
srom_1(44734) <= 1945427;
srom_1(44735) <= 1592909;
srom_1(44736) <= 1272258;
srom_1(44737) <= 984978;
srom_1(44738) <= 732416;
srom_1(44739) <= 515757;
srom_1(44740) <= 336016;
srom_1(44741) <= 194037;
srom_1(44742) <= 90484;
srom_1(44743) <= 25845;
srom_1(44744) <= 421;
srom_1(44745) <= 14333;
srom_1(44746) <= 67514;
srom_1(44747) <= 159715;
srom_1(44748) <= 290505;
srom_1(44749) <= 459270;
srom_1(44750) <= 665218;
srom_1(44751) <= 907383;
srom_1(44752) <= 1184631;
srom_1(44753) <= 1495660;
srom_1(44754) <= 1839013;
srom_1(44755) <= 2213080;
srom_1(44756) <= 2616105;
srom_1(44757) <= 3046200;
srom_1(44758) <= 3501347;
srom_1(44759) <= 3979412;
srom_1(44760) <= 4478153;
srom_1(44761) <= 4995232;
srom_1(44762) <= 5528223;
srom_1(44763) <= 6074628;
srom_1(44764) <= 6631884;
srom_1(44765) <= 7197377;
srom_1(44766) <= 7768457;
srom_1(44767) <= 8342445;
srom_1(44768) <= 8916649;
srom_1(44769) <= 9488377;
srom_1(44770) <= 10054948;
srom_1(44771) <= 10613705;
srom_1(44772) <= 11162028;
srom_1(44773) <= 11697345;
srom_1(44774) <= 12217146;
srom_1(44775) <= 12718994;
srom_1(44776) <= 13200535;
srom_1(44777) <= 13659512;
srom_1(44778) <= 14093771;
srom_1(44779) <= 14501277;
srom_1(44780) <= 14880119;
srom_1(44781) <= 15228519;
srom_1(44782) <= 15544845;
srom_1(44783) <= 15827613;
srom_1(44784) <= 16075497;
srom_1(44785) <= 16287334;
srom_1(44786) <= 16462132;
srom_1(44787) <= 16599069;
srom_1(44788) <= 16697506;
srom_1(44789) <= 16756979;
srom_1(44790) <= 16777209;
srom_1(44791) <= 16758103;
srom_1(44792) <= 16699750;
srom_1(44793) <= 16602422;
srom_1(44794) <= 16466577;
srom_1(44795) <= 16292852;
srom_1(44796) <= 16082061;
srom_1(44797) <= 15835193;
srom_1(44798) <= 15553405;
srom_1(44799) <= 15238019;
srom_1(44800) <= 14890513;
srom_1(44801) <= 14512518;
srom_1(44802) <= 14105806;
srom_1(44803) <= 13672284;
srom_1(44804) <= 13213985;
srom_1(44805) <= 12733058;
srom_1(44806) <= 12231759;
srom_1(44807) <= 11712437;
srom_1(44808) <= 11177530;
srom_1(44809) <= 10629543;
srom_1(44810) <= 10071049;
srom_1(44811) <= 9504664;
srom_1(44812) <= 8933047;
srom_1(44813) <= 8358876;
srom_1(44814) <= 7784844;
srom_1(44815) <= 7213644;
srom_1(44816) <= 6647954;
srom_1(44817) <= 6090426;
srom_1(44818) <= 5543675;
srom_1(44819) <= 5010265;
srom_1(44820) <= 4492697;
srom_1(44821) <= 3993398;
srom_1(44822) <= 3514710;
srom_1(44823) <= 3058878;
srom_1(44824) <= 2628038;
srom_1(44825) <= 2224212;
srom_1(44826) <= 1849292;
srom_1(44827) <= 1505038;
srom_1(44828) <= 1193063;
srom_1(44829) <= 914831;
srom_1(44830) <= 671645;
srom_1(44831) <= 464647;
srom_1(44832) <= 294807;
srom_1(44833) <= 162922;
srom_1(44834) <= 69610;
srom_1(44835) <= 15309;
srom_1(44836) <= 272;
srom_1(44837) <= 24572;
srom_1(44838) <= 88093;
srom_1(44839) <= 190539;
srom_1(44840) <= 331428;
srom_1(44841) <= 510100;
srom_1(44842) <= 725716;
srom_1(44843) <= 977267;
srom_1(44844) <= 1263572;
srom_1(44845) <= 1583289;
srom_1(44846) <= 1934918;
srom_1(44847) <= 2316811;
srom_1(44848) <= 2727177;
srom_1(44849) <= 3164091;
srom_1(44850) <= 3625504;
srom_1(44851) <= 4109253;
srom_1(44852) <= 4613070;
srom_1(44853) <= 5134592;
srom_1(44854) <= 5671372;
srom_1(44855) <= 6220895;
srom_1(44856) <= 6780583;
srom_1(44857) <= 7347811;
srom_1(44858) <= 7919920;
srom_1(44859) <= 8494227;
srom_1(44860) <= 9068039;
srom_1(44861) <= 9638664;
srom_1(44862) <= 10203428;
srom_1(44863) <= 10759681;
srom_1(44864) <= 11304816;
srom_1(44865) <= 11836275;
srom_1(44866) <= 12351567;
srom_1(44867) <= 12848275;
srom_1(44868) <= 13324071;
srom_1(44869) <= 13776722;
srom_1(44870) <= 14204107;
srom_1(44871) <= 14604221;
srom_1(44872) <= 14975187;
srom_1(44873) <= 15315267;
srom_1(44874) <= 15622866;
srom_1(44875) <= 15896540;
srom_1(44876) <= 16135007;
srom_1(44877) <= 16337149;
srom_1(44878) <= 16502017;
srom_1(44879) <= 16628839;
srom_1(44880) <= 16717019;
srom_1(44881) <= 16766145;
srom_1(44882) <= 16775985;
srom_1(44883) <= 16746494;
srom_1(44884) <= 16677810;
srom_1(44885) <= 16570255;
srom_1(44886) <= 16424334;
srom_1(44887) <= 16240730;
srom_1(44888) <= 16020305;
srom_1(44889) <= 15764093;
srom_1(44890) <= 15473294;
srom_1(44891) <= 15149272;
srom_1(44892) <= 14793548;
srom_1(44893) <= 14407789;
srom_1(44894) <= 13993803;
srom_1(44895) <= 13553533;
srom_1(44896) <= 13089043;
srom_1(44897) <= 12602511;
srom_1(44898) <= 12096218;
srom_1(44899) <= 11572539;
srom_1(44900) <= 11033930;
srom_1(44901) <= 10482915;
srom_1(44902) <= 9922080;
srom_1(44903) <= 9354054;
srom_1(44904) <= 8781500;
srom_1(44905) <= 8207104;
srom_1(44906) <= 7633560;
srom_1(44907) <= 7063556;
srom_1(44908) <= 6499765;
srom_1(44909) <= 5944832;
srom_1(44910) <= 5401359;
srom_1(44911) <= 4871893;
srom_1(44912) <= 4358919;
srom_1(44913) <= 3864842;
srom_1(44914) <= 3391978;
srom_1(44915) <= 2942545;
srom_1(44916) <= 2518650;
srom_1(44917) <= 2122282;
srom_1(44918) <= 1755298;
srom_1(44919) <= 1419421;
srom_1(44920) <= 1116224;
srom_1(44921) <= 847130;
srom_1(44922) <= 613401;
srom_1(44923) <= 416132;
srom_1(44924) <= 256249;
srom_1(44925) <= 134501;
srom_1(44926) <= 51460;
srom_1(44927) <= 7514;
srom_1(44928) <= 2870;
srom_1(44929) <= 37550;
srom_1(44930) <= 111391;
srom_1(44931) <= 224046;
srom_1(44932) <= 374988;
srom_1(44933) <= 563509;
srom_1(44934) <= 788724;
srom_1(44935) <= 1049577;
srom_1(44936) <= 1344846;
srom_1(44937) <= 1673145;
srom_1(44938) <= 2032936;
srom_1(44939) <= 2422530;
srom_1(44940) <= 2840102;
srom_1(44941) <= 3283692;
srom_1(44942) <= 3751221;
srom_1(44943) <= 4240496;
srom_1(44944) <= 4749223;
srom_1(44945) <= 5275017;
srom_1(44946) <= 5815411;
srom_1(44947) <= 6367872;
srom_1(44948) <= 6929808;
srom_1(44949) <= 7498586;
srom_1(44950) <= 8071537;
srom_1(44951) <= 8645975;
srom_1(44952) <= 9219206;
srom_1(44953) <= 9788542;
srom_1(44954) <= 10351313;
srom_1(44955) <= 10904881;
srom_1(44956) <= 11446649;
srom_1(44957) <= 11974076;
srom_1(44958) <= 12484691;
srom_1(44959) <= 12976097;
srom_1(44960) <= 13445991;
srom_1(44961) <= 13892169;
srom_1(44962) <= 14312539;
srom_1(44963) <= 14705129;
srom_1(44964) <= 15068099;
srom_1(44965) <= 15399747;
srom_1(44966) <= 15698517;
srom_1(44967) <= 15963009;
srom_1(44968) <= 16191981;
srom_1(44969) <= 16384361;
srom_1(44970) <= 16539246;
srom_1(44971) <= 16655910;
srom_1(44972) <= 16733806;
srom_1(44973) <= 16772568;
srom_1(44974) <= 16772014;
srom_1(44975) <= 16732149;
srom_1(44976) <= 16653157;
srom_1(44977) <= 16535410;
srom_1(44978) <= 16379460;
srom_1(44979) <= 16186038;
srom_1(44980) <= 15956051;
srom_1(44981) <= 15690578;
srom_1(44982) <= 15390864;
srom_1(44983) <= 15058313;
srom_1(44984) <= 14694486;
srom_1(44985) <= 14301088;
srom_1(44986) <= 13879965;
srom_1(44987) <= 13433091;
srom_1(44988) <= 12962562;
srom_1(44989) <= 12470583;
srom_1(44990) <= 11959463;
srom_1(44991) <= 11431598;
srom_1(44992) <= 10889464;
srom_1(44993) <= 10335602;
srom_1(44994) <= 9772610;
srom_1(44995) <= 9203127;
srom_1(44996) <= 8629826;
srom_1(44997) <= 8055393;
srom_1(44998) <= 7482522;
srom_1(44999) <= 6913901;
srom_1(45000) <= 6352195;
srom_1(45001) <= 5800038;
srom_1(45002) <= 5260020;
srom_1(45003) <= 4734673;
srom_1(45004) <= 4226461;
srom_1(45005) <= 3737766;
srom_1(45006) <= 3270881;
srom_1(45007) <= 2827995;
srom_1(45008) <= 2411184;
srom_1(45009) <= 2022403;
srom_1(45010) <= 1663476;
srom_1(45011) <= 1336085;
srom_1(45012) <= 1041766;
srom_1(45013) <= 781898;
srom_1(45014) <= 557701;
srom_1(45015) <= 370226;
srom_1(45016) <= 220352;
srom_1(45017) <= 108782;
srom_1(45018) <= 36038;
srom_1(45019) <= 2463;
srom_1(45020) <= 8213;
srom_1(45021) <= 53262;
srom_1(45022) <= 137398;
srom_1(45023) <= 260227;
srom_1(45024) <= 421172;
srom_1(45025) <= 619480;
srom_1(45026) <= 854219;
srom_1(45027) <= 1124290;
srom_1(45028) <= 1428426;
srom_1(45029) <= 1765201;
srom_1(45030) <= 2133035;
srom_1(45031) <= 2530203;
srom_1(45032) <= 2954844;
srom_1(45033) <= 3404965;
srom_1(45034) <= 3878456;
srom_1(45035) <= 4373097;
srom_1(45036) <= 4886568;
srom_1(45037) <= 5416462;
srom_1(45038) <= 5960292;
srom_1(45039) <= 6515510;
srom_1(45040) <= 7079512;
srom_1(45041) <= 7649652;
srom_1(45042) <= 8223258;
srom_1(45043) <= 8797639;
srom_1(45044) <= 9370101;
srom_1(45045) <= 9937962;
srom_1(45046) <= 10498556;
srom_1(45047) <= 11049257;
srom_1(45048) <= 11587481;
srom_1(45049) <= 12110704;
srom_1(45050) <= 12616473;
srom_1(45051) <= 13102416;
srom_1(45052) <= 13566255;
srom_1(45053) <= 14005813;
srom_1(45054) <= 14419031;
srom_1(45055) <= 14803970;
srom_1(45056) <= 15158825;
srom_1(45057) <= 15481932;
srom_1(45058) <= 15771776;
srom_1(45059) <= 16026998;
srom_1(45060) <= 16246401;
srom_1(45061) <= 16428956;
srom_1(45062) <= 16573807;
srom_1(45063) <= 16680275;
srom_1(45064) <= 16747860;
srom_1(45065) <= 16776246;
srom_1(45066) <= 16765299;
srom_1(45067) <= 16715071;
srom_1(45068) <= 16625798;
srom_1(45069) <= 16497898;
srom_1(45070) <= 16331970;
srom_1(45071) <= 16128793;
srom_1(45072) <= 15889320;
srom_1(45073) <= 15614673;
srom_1(45074) <= 15306141;
srom_1(45075) <= 14965170;
srom_1(45076) <= 14593359;
srom_1(45077) <= 14192452;
srom_1(45078) <= 13764329;
srom_1(45079) <= 13310997;
srom_1(45080) <= 12834583;
srom_1(45081) <= 12337320;
srom_1(45082) <= 11821540;
srom_1(45083) <= 11289661;
srom_1(45084) <= 10744179;
srom_1(45085) <= 10187651;
srom_1(45086) <= 9622686;
srom_1(45087) <= 9051934;
srom_1(45088) <= 8478072;
srom_1(45089) <= 7903790;
srom_1(45090) <= 7331781;
srom_1(45091) <= 6764729;
srom_1(45092) <= 6205291;
srom_1(45093) <= 5656092;
srom_1(45094) <= 5119706;
srom_1(45095) <= 4598649;
srom_1(45096) <= 4095365;
srom_1(45097) <= 3612213;
srom_1(45098) <= 3151460;
srom_1(45099) <= 2715265;
srom_1(45100) <= 2305674;
srom_1(45101) <= 1924609;
srom_1(45102) <= 1573855;
srom_1(45103) <= 1255058;
srom_1(45104) <= 969713;
srom_1(45105) <= 719157;
srom_1(45106) <= 504566;
srom_1(45107) <= 326946;
srom_1(45108) <= 187130;
srom_1(45109) <= 85774;
srom_1(45110) <= 23352;
srom_1(45111) <= 158;
srom_1(45112) <= 16300;
srom_1(45113) <= 71703;
srom_1(45114) <= 166106;
srom_1(45115) <= 299068;
srom_1(45116) <= 469964;
srom_1(45117) <= 677994;
srom_1(45118) <= 922181;
srom_1(45119) <= 1201381;
srom_1(45120) <= 1514285;
srom_1(45121) <= 1859424;
srom_1(45122) <= 2235181;
srom_1(45123) <= 2639794;
srom_1(45124) <= 3071364;
srom_1(45125) <= 3527869;
srom_1(45126) <= 4007168;
srom_1(45127) <= 4507013;
srom_1(45128) <= 5025060;
srom_1(45129) <= 5558879;
srom_1(45130) <= 6105969;
srom_1(45131) <= 6663762;
srom_1(45132) <= 7229644;
srom_1(45133) <= 7800960;
srom_1(45134) <= 8375032;
srom_1(45135) <= 8949168;
srom_1(45136) <= 9520675;
srom_1(45137) <= 10086874;
srom_1(45138) <= 10645109;
srom_1(45139) <= 11192762;
srom_1(45140) <= 11727266;
srom_1(45141) <= 12246113;
srom_1(45142) <= 12746871;
srom_1(45143) <= 13227192;
srom_1(45144) <= 13684823;
srom_1(45145) <= 14117619;
srom_1(45146) <= 14523549;
srom_1(45147) <= 14900710;
srom_1(45148) <= 15247334;
srom_1(45149) <= 15561794;
srom_1(45150) <= 15842618;
srom_1(45151) <= 16088486;
srom_1(45152) <= 16298248;
srom_1(45153) <= 16470918;
srom_1(45154) <= 16605688;
srom_1(45155) <= 16701925;
srom_1(45156) <= 16759178;
srom_1(45157) <= 16777178;
srom_1(45158) <= 16755842;
srom_1(45159) <= 16695268;
srom_1(45160) <= 16595742;
srom_1(45161) <= 16457730;
srom_1(45162) <= 16281879;
srom_1(45163) <= 16069014;
srom_1(45164) <= 15820132;
srom_1(45165) <= 15536402;
srom_1(45166) <= 15219153;
srom_1(45167) <= 14869874;
srom_1(45168) <= 14490201;
srom_1(45169) <= 14081916;
srom_1(45170) <= 13646933;
srom_1(45171) <= 13187292;
srom_1(45172) <= 12705149;
srom_1(45173) <= 12202763;
srom_1(45174) <= 11682492;
srom_1(45175) <= 11146774;
srom_1(45176) <= 10598123;
srom_1(45177) <= 10039110;
srom_1(45178) <= 9472358;
srom_1(45179) <= 8900524;
srom_1(45180) <= 8326288;
srom_1(45181) <= 7752346;
srom_1(45182) <= 7181387;
srom_1(45183) <= 6616088;
srom_1(45184) <= 6059102;
srom_1(45185) <= 5513040;
srom_1(45186) <= 4980462;
srom_1(45187) <= 4463866;
srom_1(45188) <= 3965675;
srom_1(45189) <= 3488224;
srom_1(45190) <= 3033753;
srom_1(45191) <= 2604393;
srom_1(45192) <= 2202156;
srom_1(45193) <= 1828931;
srom_1(45194) <= 1486465;
srom_1(45195) <= 1176367;
srom_1(45196) <= 900088;
srom_1(45197) <= 658927;
srom_1(45198) <= 454012;
srom_1(45199) <= 286305;
srom_1(45200) <= 156593;
srom_1(45201) <= 65483;
srom_1(45202) <= 13404;
srom_1(45203) <= 599;
srom_1(45204) <= 27128;
srom_1(45205) <= 92866;
srom_1(45206) <= 197507;
srom_1(45207) <= 340558;
srom_1(45208) <= 521349;
srom_1(45209) <= 739033;
srom_1(45210) <= 992588;
srom_1(45211) <= 1280826;
srom_1(45212) <= 1602394;
srom_1(45213) <= 1955785;
srom_1(45214) <= 2339342;
srom_1(45215) <= 2751266;
srom_1(45216) <= 3189626;
srom_1(45217) <= 3652365;
srom_1(45218) <= 4137314;
srom_1(45219) <= 4642199;
srom_1(45220) <= 5164652;
srom_1(45221) <= 5702223;
srom_1(45222) <= 6252392;
srom_1(45223) <= 6812578;
srom_1(45224) <= 7380155;
srom_1(45225) <= 7952461;
srom_1(45226) <= 8526812;
srom_1(45227) <= 9100514;
srom_1(45228) <= 9670879;
srom_1(45229) <= 10235230;
srom_1(45230) <= 10790922;
srom_1(45231) <= 11335349;
srom_1(45232) <= 11865957;
srom_1(45233) <= 12380259;
srom_1(45234) <= 12875843;
srom_1(45235) <= 13350384;
srom_1(45236) <= 13801658;
srom_1(45237) <= 14227549;
srom_1(45238) <= 14626058;
srom_1(45239) <= 14995318;
srom_1(45240) <= 15333597;
srom_1(45241) <= 15639308;
srom_1(45242) <= 15911019;
srom_1(45243) <= 16147454;
srom_1(45244) <= 16347505;
srom_1(45245) <= 16510234;
srom_1(45246) <= 16634878;
srom_1(45247) <= 16720853;
srom_1(45248) <= 16767755;
srom_1(45249) <= 16775364;
srom_1(45250) <= 16743645;
srom_1(45251) <= 16672746;
srom_1(45252) <= 16563000;
srom_1(45253) <= 16414921;
srom_1(45254) <= 16229204;
srom_1(45255) <= 16006720;
srom_1(45256) <= 15748512;
srom_1(45257) <= 15455791;
srom_1(45258) <= 15129929;
srom_1(45259) <= 14772455;
srom_1(45260) <= 14385045;
srom_1(45261) <= 13969516;
srom_1(45262) <= 13527816;
srom_1(45263) <= 13062016;
srom_1(45264) <= 12574301;
srom_1(45265) <= 12066958;
srom_1(45266) <= 11542366;
srom_1(45267) <= 11002985;
srom_1(45268) <= 10451344;
srom_1(45269) <= 9890030;
srom_1(45270) <= 9321675;
srom_1(45271) <= 8748945;
srom_1(45272) <= 8174526;
srom_1(45273) <= 7601110;
srom_1(45274) <= 7031387;
srom_1(45275) <= 6468028;
srom_1(45276) <= 5913676;
srom_1(45277) <= 5370930;
srom_1(45278) <= 4842334;
srom_1(45279) <= 4330368;
srom_1(45280) <= 3837433;
srom_1(45281) <= 3365839;
srom_1(45282) <= 2917800;
srom_1(45283) <= 2495414;
srom_1(45284) <= 2100664;
srom_1(45285) <= 1735400;
srom_1(45286) <= 1401335;
srom_1(45287) <= 1100036;
srom_1(45288) <= 832916;
srom_1(45289) <= 601227;
srom_1(45290) <= 406055;
srom_1(45291) <= 248317;
srom_1(45292) <= 128751;
srom_1(45293) <= 47918;
srom_1(45294) <= 6198;
srom_1(45295) <= 3786;
srom_1(45296) <= 40693;
srom_1(45297) <= 116746;
srom_1(45298) <= 231589;
srom_1(45299) <= 384683;
srom_1(45300) <= 575310;
srom_1(45301) <= 802576;
srom_1(45302) <= 1065416;
srom_1(45303) <= 1362597;
srom_1(45304) <= 1692725;
srom_1(45305) <= 2054252;
srom_1(45306) <= 2445484;
srom_1(45307) <= 2864585;
srom_1(45308) <= 3309589;
srom_1(45309) <= 3778411;
srom_1(45310) <= 4268852;
srom_1(45311) <= 4778612;
srom_1(45312) <= 5305300;
srom_1(45313) <= 5846447;
srom_1(45314) <= 6399515;
srom_1(45315) <= 6961911;
srom_1(45316) <= 7530996;
srom_1(45317) <= 8104104;
srom_1(45318) <= 8678545;
srom_1(45319) <= 9251627;
srom_1(45320) <= 9820662;
srom_1(45321) <= 10382982;
srom_1(45322) <= 10935949;
srom_1(45323) <= 11476971;
srom_1(45324) <= 12003510;
srom_1(45325) <= 12513098;
srom_1(45326) <= 13003345;
srom_1(45327) <= 13471952;
srom_1(45328) <= 13916721;
srom_1(45329) <= 14335567;
srom_1(45330) <= 14726525;
srom_1(45331) <= 15087763;
srom_1(45332) <= 15417586;
srom_1(45333) <= 15714448;
srom_1(45334) <= 15976957;
srom_1(45335) <= 16203881;
srom_1(45336) <= 16394157;
srom_1(45337) <= 16546892;
srom_1(45338) <= 16661369;
srom_1(45339) <= 16737053;
srom_1(45340) <= 16773589;
srom_1(45341) <= 16770804;
srom_1(45342) <= 16728712;
srom_1(45343) <= 16647511;
srom_1(45344) <= 16527581;
srom_1(45345) <= 16369484;
srom_1(45346) <= 16173962;
srom_1(45347) <= 15941932;
srom_1(45348) <= 15674482;
srom_1(45349) <= 15372866;
srom_1(45350) <= 15038498;
srom_1(45351) <= 14672947;
srom_1(45352) <= 14277926;
srom_1(45353) <= 13855289;
srom_1(45354) <= 13407016;
srom_1(45355) <= 12935210;
srom_1(45356) <= 12442083;
srom_1(45357) <= 11929949;
srom_1(45358) <= 11401207;
srom_1(45359) <= 10858339;
srom_1(45360) <= 10303889;
srom_1(45361) <= 9740458;
srom_1(45362) <= 9170687;
srom_1(45363) <= 8597249;
srom_1(45364) <= 8022833;
srom_1(45365) <= 7450132;
srom_1(45366) <= 6881832;
srom_1(45367) <= 6320597;
srom_1(45368) <= 5769060;
srom_1(45369) <= 5229807;
srom_1(45370) <= 4705367;
srom_1(45371) <= 4198199;
srom_1(45372) <= 3710681;
srom_1(45373) <= 3245099;
srom_1(45374) <= 2803637;
srom_1(45375) <= 2388365;
srom_1(45376) <= 2001230;
srom_1(45377) <= 1644048;
srom_1(45378) <= 1318493;
srom_1(45379) <= 1026092;
srom_1(45380) <= 768217;
srom_1(45381) <= 546077;
srom_1(45382) <= 360712;
srom_1(45383) <= 212994;
srom_1(45384) <= 103613;
srom_1(45385) <= 33084;
srom_1(45386) <= 1737;
srom_1(45387) <= 9718;
srom_1(45388) <= 56991;
srom_1(45389) <= 143334;
srom_1(45390) <= 268342;
srom_1(45391) <= 431428;
srom_1(45392) <= 631829;
srom_1(45393) <= 868603;
srom_1(45394) <= 1140642;
srom_1(45395) <= 1446668;
srom_1(45396) <= 1785248;
srom_1(45397) <= 2154794;
srom_1(45398) <= 2553571;
srom_1(45399) <= 2979711;
srom_1(45400) <= 3431216;
srom_1(45401) <= 3905967;
srom_1(45402) <= 4401739;
srom_1(45403) <= 4916207;
srom_1(45404) <= 5446958;
srom_1(45405) <= 5991503;
srom_1(45406) <= 6547289;
srom_1(45407) <= 7111710;
srom_1(45408) <= 7682119;
srom_1(45409) <= 8255840;
srom_1(45410) <= 8830184;
srom_1(45411) <= 9402458;
srom_1(45412) <= 9969977;
srom_1(45413) <= 10530081;
srom_1(45414) <= 11080142;
srom_1(45415) <= 11617582;
srom_1(45416) <= 12139880;
srom_1(45417) <= 12644587;
srom_1(45418) <= 13129337;
srom_1(45419) <= 13591855;
srom_1(45420) <= 14029974;
srom_1(45421) <= 14441638;
srom_1(45422) <= 14824918;
srom_1(45423) <= 15178015;
srom_1(45424) <= 15499275;
srom_1(45425) <= 15787190;
srom_1(45426) <= 16040411;
srom_1(45427) <= 16257750;
srom_1(45428) <= 16438187;
srom_1(45429) <= 16580878;
srom_1(45430) <= 16685152;
srom_1(45431) <= 16750521;
srom_1(45432) <= 16776678;
srom_1(45433) <= 16763500;
srom_1(45434) <= 16711049;
srom_1(45435) <= 16619572;
srom_1(45436) <= 16489497;
srom_1(45437) <= 16321434;
srom_1(45438) <= 16116172;
srom_1(45439) <= 15874672;
srom_1(45440) <= 15598067;
srom_1(45441) <= 15287655;
srom_1(45442) <= 14944890;
srom_1(45443) <= 14571382;
srom_1(45444) <= 14168879;
srom_1(45445) <= 13739272;
srom_1(45446) <= 13284573;
srom_1(45447) <= 12806915;
srom_1(45448) <= 12308538;
srom_1(45449) <= 11791780;
srom_1(45450) <= 11259062;
srom_1(45451) <= 10712885;
srom_1(45452) <= 10155807;
srom_1(45453) <= 9590443;
srom_1(45454) <= 9019443;
srom_1(45455) <= 8445485;
srom_1(45456) <= 7871260;
srom_1(45457) <= 7299461;
srom_1(45458) <= 6732770;
srom_1(45459) <= 6173843;
srom_1(45460) <= 5625302;
srom_1(45461) <= 5089719;
srom_1(45462) <= 4569606;
srom_1(45463) <= 4067401;
srom_1(45464) <= 3585460;
srom_1(45465) <= 3126043;
srom_1(45466) <= 2691303;
srom_1(45467) <= 2283280;
srom_1(45468) <= 1903887;
srom_1(45469) <= 1554904;
srom_1(45470) <= 1237965;
srom_1(45471) <= 954559;
srom_1(45472) <= 706013;
srom_1(45473) <= 493494;
srom_1(45474) <= 317998;
srom_1(45475) <= 180347;
srom_1(45476) <= 81188;
srom_1(45477) <= 20985;
srom_1(45478) <= 21;
srom_1(45479) <= 18394;
srom_1(45480) <= 76017;
srom_1(45481) <= 172621;
srom_1(45482) <= 307753;
srom_1(45483) <= 480779;
srom_1(45484) <= 690887;
srom_1(45485) <= 937092;
srom_1(45486) <= 1218240;
srom_1(45487) <= 1533013;
srom_1(45488) <= 1879933;
srom_1(45489) <= 2257375;
srom_1(45490) <= 2663569;
srom_1(45491) <= 3096609;
srom_1(45492) <= 3554465;
srom_1(45493) <= 4034990;
srom_1(45494) <= 4535931;
srom_1(45495) <= 5054938;
srom_1(45496) <= 5589578;
srom_1(45497) <= 6137344;
srom_1(45498) <= 6695666;
srom_1(45499) <= 7261928;
srom_1(45500) <= 7833472;
srom_1(45501) <= 8407620;
srom_1(45502) <= 8981679;
srom_1(45503) <= 9552956;
srom_1(45504) <= 10118774;
srom_1(45505) <= 10676478;
srom_1(45506) <= 11223454;
srom_1(45507) <= 11757136;
srom_1(45508) <= 12275022;
srom_1(45509) <= 12774683;
srom_1(45510) <= 13253776;
srom_1(45511) <= 13710055;
srom_1(45512) <= 14141380;
srom_1(45513) <= 14545728;
srom_1(45514) <= 14921203;
srom_1(45515) <= 15266044;
srom_1(45516) <= 15578635;
srom_1(45517) <= 15857510;
srom_1(45518) <= 16101360;
srom_1(45519) <= 16309042;
srom_1(45520) <= 16479583;
srom_1(45521) <= 16612182;
srom_1(45522) <= 16706218;
srom_1(45523) <= 16761250;
srom_1(45524) <= 16777020;
srom_1(45525) <= 16753454;
srom_1(45526) <= 16690662;
srom_1(45527) <= 16588939;
srom_1(45528) <= 16448761;
srom_1(45529) <= 16270787;
srom_1(45530) <= 16055851;
srom_1(45531) <= 15804960;
srom_1(45532) <= 15519291;
srom_1(45533) <= 15200185;
srom_1(45534) <= 14849136;
srom_1(45535) <= 14467792;
srom_1(45536) <= 14057940;
srom_1(45537) <= 13621503;
srom_1(45538) <= 13160527;
srom_1(45539) <= 12677174;
srom_1(45540) <= 12173710;
srom_1(45541) <= 11652497;
srom_1(45542) <= 11115978;
srom_1(45543) <= 10566669;
srom_1(45544) <= 10007147;
srom_1(45545) <= 9440035;
srom_1(45546) <= 8867993;
srom_1(45547) <= 8293702;
srom_1(45548) <= 7719857;
srom_1(45549) <= 7149147;
srom_1(45550) <= 6584250;
srom_1(45551) <= 6027814;
srom_1(45552) <= 5482448;
srom_1(45553) <= 4950711;
srom_1(45554) <= 4435095;
srom_1(45555) <= 3938018;
srom_1(45556) <= 3461812;
srom_1(45557) <= 3008709;
srom_1(45558) <= 2580834;
srom_1(45559) <= 2180194;
srom_1(45560) <= 1808668;
srom_1(45561) <= 1467997;
srom_1(45562) <= 1159779;
srom_1(45563) <= 885459;
srom_1(45564) <= 646325;
srom_1(45565) <= 443496;
srom_1(45566) <= 277925;
srom_1(45567) <= 150388;
srom_1(45568) <= 61482;
srom_1(45569) <= 11626;
srom_1(45570) <= 1051;
srom_1(45571) <= 29809;
srom_1(45572) <= 97765;
srom_1(45573) <= 204598;
srom_1(45574) <= 349810;
srom_1(45575) <= 532718;
srom_1(45576) <= 752465;
srom_1(45577) <= 1008021;
srom_1(45578) <= 1298186;
srom_1(45579) <= 1621601;
srom_1(45580) <= 1976749;
srom_1(45581) <= 2361965;
srom_1(45582) <= 2775441;
srom_1(45583) <= 3215239;
srom_1(45584) <= 3679297;
srom_1(45585) <= 4165439;
srom_1(45586) <= 4671385;
srom_1(45587) <= 5194761;
srom_1(45588) <= 5733115;
srom_1(45589) <= 6283922;
srom_1(45590) <= 6844598;
srom_1(45591) <= 7412514;
srom_1(45592) <= 7985008;
srom_1(45593) <= 8559394;
srom_1(45594) <= 9132979;
srom_1(45595) <= 9703074;
srom_1(45596) <= 10267005;
srom_1(45597) <= 10822127;
srom_1(45598) <= 11365838;
srom_1(45599) <= 11895587;
srom_1(45600) <= 12408891;
srom_1(45601) <= 12903342;
srom_1(45602) <= 13376623;
srom_1(45603) <= 13826512;
srom_1(45604) <= 14250902;
srom_1(45605) <= 14647801;
srom_1(45606) <= 15015349;
srom_1(45607) <= 15351822;
srom_1(45608) <= 15655642;
srom_1(45609) <= 15925384;
srom_1(45610) <= 16159783;
srom_1(45611) <= 16357741;
srom_1(45612) <= 16518329;
srom_1(45613) <= 16640794;
srom_1(45614) <= 16724561;
srom_1(45615) <= 16769239;
srom_1(45616) <= 16774616;
srom_1(45617) <= 16740669;
srom_1(45618) <= 16667556;
srom_1(45619) <= 16555620;
srom_1(45620) <= 16405387;
srom_1(45621) <= 16217560;
srom_1(45622) <= 15993020;
srom_1(45623) <= 15732820;
srom_1(45624) <= 15438181;
srom_1(45625) <= 15110484;
srom_1(45626) <= 14751266;
srom_1(45627) <= 14362212;
srom_1(45628) <= 13945145;
srom_1(45629) <= 13502021;
srom_1(45630) <= 13034919;
srom_1(45631) <= 12546028;
srom_1(45632) <= 12037643;
srom_1(45633) <= 11512145;
srom_1(45634) <= 10972000;
srom_1(45635) <= 10419741;
srom_1(45636) <= 9857957;
srom_1(45637) <= 9289283;
srom_1(45638) <= 8716385;
srom_1(45639) <= 8141950;
srom_1(45640) <= 7568672;
srom_1(45641) <= 6999239;
srom_1(45642) <= 6436321;
srom_1(45643) <= 5882558;
srom_1(45644) <= 5340546;
srom_1(45645) <= 4812828;
srom_1(45646) <= 4301878;
srom_1(45647) <= 3810093;
srom_1(45648) <= 3339777;
srom_1(45649) <= 2893137;
srom_1(45650) <= 2472267;
srom_1(45651) <= 2079141;
srom_1(45652) <= 1715602;
srom_1(45653) <= 1383356;
srom_1(45654) <= 1083959;
srom_1(45655) <= 818816;
srom_1(45656) <= 589171;
srom_1(45657) <= 396100;
srom_1(45658) <= 240508;
srom_1(45659) <= 123126;
srom_1(45660) <= 44503;
srom_1(45661) <= 5009;
srom_1(45662) <= 4828;
srom_1(45663) <= 43962;
srom_1(45664) <= 122226;
srom_1(45665) <= 239255;
srom_1(45666) <= 394499;
srom_1(45667) <= 587229;
srom_1(45668) <= 816543;
srom_1(45669) <= 1081366;
srom_1(45670) <= 1380454;
srom_1(45671) <= 1712406;
srom_1(45672) <= 2075665;
srom_1(45673) <= 2468527;
srom_1(45674) <= 2889151;
srom_1(45675) <= 3335563;
srom_1(45676) <= 3805671;
srom_1(45677) <= 4297270;
srom_1(45678) <= 4808055;
srom_1(45679) <= 5335630;
srom_1(45680) <= 5877522;
srom_1(45681) <= 6431189;
srom_1(45682) <= 6994034;
srom_1(45683) <= 7563420;
srom_1(45684) <= 8136675;
srom_1(45685) <= 8711112;
srom_1(45686) <= 9284036;
srom_1(45687) <= 9852761;
srom_1(45688) <= 10414620;
srom_1(45689) <= 10966979;
srom_1(45690) <= 11507246;
srom_1(45691) <= 12032890;
srom_1(45692) <= 12541444;
srom_1(45693) <= 13030524;
srom_1(45694) <= 13497836;
srom_1(45695) <= 13941190;
srom_1(45696) <= 14358505;
srom_1(45697) <= 14747826;
srom_1(45698) <= 15107326;
srom_1(45699) <= 15435320;
srom_1(45700) <= 15730269;
srom_1(45701) <= 15990790;
srom_1(45702) <= 16215663;
srom_1(45703) <= 16403831;
srom_1(45704) <= 16554414;
srom_1(45705) <= 16666704;
srom_1(45706) <= 16740175;
srom_1(45707) <= 16774483;
srom_1(45708) <= 16769467;
srom_1(45709) <= 16725150;
srom_1(45710) <= 16641740;
srom_1(45711) <= 16519628;
srom_1(45712) <= 16359388;
srom_1(45713) <= 16161769;
srom_1(45714) <= 15927699;
srom_1(45715) <= 15658276;
srom_1(45716) <= 15354763;
srom_1(45717) <= 15018584;
srom_1(45718) <= 14651314;
srom_1(45719) <= 14254676;
srom_1(45720) <= 13830530;
srom_1(45721) <= 13380865;
srom_1(45722) <= 12907789;
srom_1(45723) <= 12413522;
srom_1(45724) <= 11900380;
srom_1(45725) <= 11370771;
srom_1(45726) <= 10827177;
srom_1(45727) <= 10272148;
srom_1(45728) <= 9708286;
srom_1(45729) <= 9138236;
srom_1(45730) <= 8564670;
srom_1(45731) <= 7990279;
srom_1(45732) <= 7417756;
srom_1(45733) <= 6849785;
srom_1(45734) <= 6289031;
srom_1(45735) <= 5738122;
srom_1(45736) <= 5199642;
srom_1(45737) <= 4676116;
srom_1(45738) <= 4170000;
srom_1(45739) <= 3683666;
srom_1(45740) <= 3219395;
srom_1(45741) <= 2779364;
srom_1(45742) <= 2365637;
srom_1(45743) <= 1980154;
srom_1(45744) <= 1624722;
srom_1(45745) <= 1301008;
srom_1(45746) <= 1010530;
srom_1(45747) <= 754651;
srom_1(45748) <= 534570;
srom_1(45749) <= 351320;
srom_1(45750) <= 205759;
srom_1(45751) <= 98570;
srom_1(45752) <= 30256;
srom_1(45753) <= 1137;
srom_1(45754) <= 11350;
srom_1(45755) <= 60846;
srom_1(45756) <= 149395;
srom_1(45757) <= 276580;
srom_1(45758) <= 441805;
srom_1(45759) <= 644295;
srom_1(45760) <= 883101;
srom_1(45761) <= 1157103;
srom_1(45762) <= 1465016;
srom_1(45763) <= 1805396;
srom_1(45764) <= 2176647;
srom_1(45765) <= 2577028;
srom_1(45766) <= 3004661;
srom_1(45767) <= 3457542;
srom_1(45768) <= 3933546;
srom_1(45769) <= 4430441;
srom_1(45770) <= 4945898;
srom_1(45771) <= 5477498;
srom_1(45772) <= 6022750;
srom_1(45773) <= 6579096;
srom_1(45774) <= 7143928;
srom_1(45775) <= 7714596;
srom_1(45776) <= 8288425;
srom_1(45777) <= 8862724;
srom_1(45778) <= 9434799;
srom_1(45779) <= 10001969;
srom_1(45780) <= 10561572;
srom_1(45781) <= 11110987;
srom_1(45782) <= 11647634;
srom_1(45783) <= 12169000;
srom_1(45784) <= 12672637;
srom_1(45785) <= 13156186;
srom_1(45786) <= 13617377;
srom_1(45787) <= 14054049;
srom_1(45788) <= 14464154;
srom_1(45789) <= 14845768;
srom_1(45790) <= 15197103;
srom_1(45791) <= 15516510;
srom_1(45792) <= 15802492;
srom_1(45793) <= 16053708;
srom_1(45794) <= 16268980;
srom_1(45795) <= 16447297;
srom_1(45796) <= 16587825;
srom_1(45797) <= 16689904;
srom_1(45798) <= 16753055;
srom_1(45799) <= 16776983;
srom_1(45800) <= 16761574;
srom_1(45801) <= 16706902;
srom_1(45802) <= 16613222;
srom_1(45803) <= 16480974;
srom_1(45804) <= 16310779;
srom_1(45805) <= 16103433;
srom_1(45806) <= 15859911;
srom_1(45807) <= 15581352;
srom_1(45808) <= 15269065;
srom_1(45809) <= 14924512;
srom_1(45810) <= 14549311;
srom_1(45811) <= 14145219;
srom_1(45812) <= 13714133;
srom_1(45813) <= 13258074;
srom_1(45814) <= 12779181;
srom_1(45815) <= 12279698;
srom_1(45816) <= 11761968;
srom_1(45817) <= 11228420;
srom_1(45818) <= 10681555;
srom_1(45819) <= 10123938;
srom_1(45820) <= 9558183;
srom_1(45821) <= 8986943;
srom_1(45822) <= 8412898;
srom_1(45823) <= 7838738;
srom_1(45824) <= 7267158;
srom_1(45825) <= 6700836;
srom_1(45826) <= 6142428;
srom_1(45827) <= 5594554;
srom_1(45828) <= 5059782;
srom_1(45829) <= 4540620;
srom_1(45830) <= 4039502;
srom_1(45831) <= 3558779;
srom_1(45832) <= 3100705;
srom_1(45833) <= 2667427;
srom_1(45834) <= 2260978;
srom_1(45835) <= 1883264;
srom_1(45836) <= 1536055;
srom_1(45837) <= 1220981;
srom_1(45838) <= 939518;
srom_1(45839) <= 692986;
srom_1(45840) <= 482541;
srom_1(45841) <= 309171;
srom_1(45842) <= 173688;
srom_1(45843) <= 76728;
srom_1(45844) <= 18745;
srom_1(45845) <= 11;
srom_1(45846) <= 20614;
srom_1(45847) <= 80457;
srom_1(45848) <= 179260;
srom_1(45849) <= 316560;
srom_1(45850) <= 491712;
srom_1(45851) <= 703896;
srom_1(45852) <= 952115;
srom_1(45853) <= 1235207;
srom_1(45854) <= 1551844;
srom_1(45855) <= 1900541;
srom_1(45856) <= 2279662;
srom_1(45857) <= 2687431;
srom_1(45858) <= 3121934;
srom_1(45859) <= 3581134;
srom_1(45860) <= 4062879;
srom_1(45861) <= 4564908;
srom_1(45862) <= 5084867;
srom_1(45863) <= 5620320;
srom_1(45864) <= 6168753;
srom_1(45865) <= 6727596;
srom_1(45866) <= 7294229;
srom_1(45867) <= 7865993;
srom_1(45868) <= 8440208;
srom_1(45869) <= 9014181;
srom_1(45870) <= 9585220;
srom_1(45871) <= 10150648;
srom_1(45872) <= 10707813;
srom_1(45873) <= 11254103;
srom_1(45874) <= 11786955;
srom_1(45875) <= 12303872;
srom_1(45876) <= 12802428;
srom_1(45877) <= 13280286;
srom_1(45878) <= 13735206;
srom_1(45879) <= 14165054;
srom_1(45880) <= 14567814;
srom_1(45881) <= 14941597;
srom_1(45882) <= 15284651;
srom_1(45883) <= 15595367;
srom_1(45884) <= 15872289;
srom_1(45885) <= 16114117;
srom_1(45886) <= 16319717;
srom_1(45887) <= 16488125;
srom_1(45888) <= 16618552;
srom_1(45889) <= 16710386;
srom_1(45890) <= 16763197;
srom_1(45891) <= 16776736;
srom_1(45892) <= 16750940;
srom_1(45893) <= 16685930;
srom_1(45894) <= 16582011;
srom_1(45895) <= 16439671;
srom_1(45896) <= 16259576;
srom_1(45897) <= 16042572;
srom_1(45898) <= 15789676;
srom_1(45899) <= 15502073;
srom_1(45900) <= 15181113;
srom_1(45901) <= 14828301;
srom_1(45902) <= 14445291;
srom_1(45903) <= 14033878;
srom_1(45904) <= 13595994;
srom_1(45905) <= 13133690;
srom_1(45906) <= 12649134;
srom_1(45907) <= 12144600;
srom_1(45908) <= 11622452;
srom_1(45909) <= 11085140;
srom_1(45910) <= 10535183;
srom_1(45911) <= 9975160;
srom_1(45912) <= 9407697;
srom_1(45913) <= 8835455;
srom_1(45914) <= 8261117;
srom_1(45915) <= 7687378;
srom_1(45916) <= 7116926;
srom_1(45917) <= 6552438;
srom_1(45918) <= 5996561;
srom_1(45919) <= 5451901;
srom_1(45920) <= 4921012;
srom_1(45921) <= 4406383;
srom_1(45922) <= 3910429;
srom_1(45923) <= 3435474;
srom_1(45924) <= 2983746;
srom_1(45925) <= 2557364;
srom_1(45926) <= 2158326;
srom_1(45927) <= 1788504;
srom_1(45928) <= 1449633;
srom_1(45929) <= 1143300;
srom_1(45930) <= 870943;
srom_1(45931) <= 633840;
srom_1(45932) <= 433101;
srom_1(45933) <= 269668;
srom_1(45934) <= 144307;
srom_1(45935) <= 57607;
srom_1(45936) <= 9974;
srom_1(45937) <= 1631;
srom_1(45938) <= 32617;
srom_1(45939) <= 102788;
srom_1(45940) <= 211814;
srom_1(45941) <= 359183;
srom_1(45942) <= 544205;
srom_1(45943) <= 766012;
srom_1(45944) <= 1023565;
srom_1(45945) <= 1315654;
srom_1(45946) <= 1640911;
srom_1(45947) <= 1997810;
srom_1(45948) <= 2384678;
srom_1(45949) <= 2799700;
srom_1(45950) <= 3240931;
srom_1(45951) <= 3706301;
srom_1(45952) <= 4193628;
srom_1(45953) <= 4700626;
srom_1(45954) <= 5224919;
srom_1(45955) <= 5764047;
srom_1(45956) <= 6315483;
srom_1(45957) <= 6876640;
srom_1(45958) <= 7444888;
srom_1(45959) <= 8017561;
srom_1(45960) <= 8591974;
srom_1(45961) <= 9165433;
srom_1(45962) <= 9735249;
srom_1(45963) <= 10298751;
srom_1(45964) <= 10853295;
srom_1(45965) <= 11396281;
srom_1(45966) <= 11925164;
srom_1(45967) <= 12437462;
srom_1(45968) <= 12930774;
srom_1(45969) <= 13402786;
srom_1(45970) <= 13851285;
srom_1(45971) <= 14274167;
srom_1(45972) <= 14669450;
srom_1(45973) <= 15035280;
srom_1(45974) <= 15369942;
srom_1(45975) <= 15671865;
srom_1(45976) <= 15939635;
srom_1(45977) <= 16171996;
srom_1(45978) <= 16367857;
srom_1(45979) <= 16526301;
srom_1(45980) <= 16646585;
srom_1(45981) <= 16728144;
srom_1(45982) <= 16770596;
srom_1(45983) <= 16773742;
srom_1(45984) <= 16737568;
srom_1(45985) <= 16662242;
srom_1(45986) <= 16548118;
srom_1(45987) <= 16395732;
srom_1(45988) <= 16205797;
srom_1(45989) <= 15979205;
srom_1(45990) <= 15717018;
srom_1(45991) <= 15420465;
srom_1(45992) <= 15090938;
srom_1(45993) <= 14729981;
srom_1(45994) <= 14339288;
srom_1(45995) <= 13920689;
srom_1(45996) <= 13476149;
srom_1(45997) <= 13007751;
srom_1(45998) <= 12517693;
srom_1(45999) <= 12008272;
srom_1(46000) <= 11481877;
srom_1(46001) <= 10940977;
srom_1(46002) <= 10388108;
srom_1(46003) <= 9825862;
srom_1(46004) <= 9256877;
srom_1(46005) <= 8683820;
srom_1(46006) <= 8109378;
srom_1(46007) <= 7536246;
srom_1(46008) <= 6967112;
srom_1(46009) <= 6404643;
srom_1(46010) <= 5851477;
srom_1(46011) <= 5310209;
srom_1(46012) <= 4783376;
srom_1(46013) <= 4273450;
srom_1(46014) <= 3782821;
srom_1(46015) <= 3313791;
srom_1(46016) <= 2868557;
srom_1(46017) <= 2449210;
srom_1(46018) <= 2057714;
srom_1(46019) <= 1695905;
srom_1(46020) <= 1365482;
srom_1(46021) <= 1067992;
srom_1(46022) <= 804831;
srom_1(46023) <= 577232;
srom_1(46024) <= 386264;
srom_1(46025) <= 232822;
srom_1(46026) <= 117625;
srom_1(46027) <= 41214;
srom_1(46028) <= 3946;
srom_1(46029) <= 5997;
srom_1(46030) <= 47357;
srom_1(46031) <= 127832;
srom_1(46032) <= 247044;
srom_1(46033) <= 404435;
srom_1(46034) <= 599266;
srom_1(46035) <= 830625;
srom_1(46036) <= 1097425;
srom_1(46037) <= 1398416;
srom_1(46038) <= 1732187;
srom_1(46039) <= 2097172;
srom_1(46040) <= 2491660;
srom_1(46041) <= 2913800;
srom_1(46042) <= 3361614;
srom_1(46043) <= 3833000;
srom_1(46044) <= 4325750;
srom_1(46045) <= 4837552;
srom_1(46046) <= 5366006;
srom_1(46047) <= 5908634;
srom_1(46048) <= 6462891;
srom_1(46049) <= 7026179;
srom_1(46050) <= 7595856;
srom_1(46051) <= 8169250;
srom_1(46052) <= 8743673;
srom_1(46053) <= 9316431;
srom_1(46054) <= 9884837;
srom_1(46055) <= 10446228;
srom_1(46056) <= 10997970;
srom_1(46057) <= 11537475;
srom_1(46058) <= 12062214;
srom_1(46059) <= 12569727;
srom_1(46060) <= 13057633;
srom_1(46061) <= 13523644;
srom_1(46062) <= 13965575;
srom_1(46063) <= 14381354;
srom_1(46064) <= 14769030;
srom_1(46065) <= 15126787;
srom_1(46066) <= 15452946;
srom_1(46067) <= 15745978;
srom_1(46068) <= 16004509;
srom_1(46069) <= 16227326;
srom_1(46070) <= 16413385;
srom_1(46071) <= 16561813;
srom_1(46072) <= 16671914;
srom_1(46073) <= 16743171;
srom_1(46074) <= 16775251;
srom_1(46075) <= 16768004;
srom_1(46076) <= 16721462;
srom_1(46077) <= 16635845;
srom_1(46078) <= 16511554;
srom_1(46079) <= 16349171;
srom_1(46080) <= 16149458;
srom_1(46081) <= 15913353;
srom_1(46082) <= 15641961;
srom_1(46083) <= 15336555;
srom_1(46084) <= 14998569;
srom_1(46085) <= 14629586;
srom_1(46086) <= 14231337;
srom_1(46087) <= 13805689;
srom_1(46088) <= 13354639;
srom_1(46089) <= 12880301;
srom_1(46090) <= 12384900;
srom_1(46091) <= 11870759;
srom_1(46092) <= 11340289;
srom_1(46093) <= 10795978;
srom_1(46094) <= 10240378;
srom_1(46095) <= 9676094;
srom_1(46096) <= 9105773;
srom_1(46097) <= 8532088;
srom_1(46098) <= 7957731;
srom_1(46099) <= 7385394;
srom_1(46100) <= 6817762;
srom_1(46101) <= 6257496;
srom_1(46102) <= 5707224;
srom_1(46103) <= 5169525;
srom_1(46104) <= 4646922;
srom_1(46105) <= 4141865;
srom_1(46106) <= 3656722;
srom_1(46107) <= 3193768;
srom_1(46108) <= 2755176;
srom_1(46109) <= 2343000;
srom_1(46110) <= 1959174;
srom_1(46111) <= 1605498;
srom_1(46112) <= 1283630;
srom_1(46113) <= 995080;
srom_1(46114) <= 741200;
srom_1(46115) <= 523182;
srom_1(46116) <= 342048;
srom_1(46117) <= 198647;
srom_1(46118) <= 93651;
srom_1(46119) <= 27553;
srom_1(46120) <= 663;
srom_1(46121) <= 13107;
srom_1(46122) <= 64827;
srom_1(46123) <= 155580;
srom_1(46124) <= 284940;
srom_1(46125) <= 452301;
srom_1(46126) <= 656878;
srom_1(46127) <= 897712;
srom_1(46128) <= 1173673;
srom_1(46129) <= 1483467;
srom_1(46130) <= 1825642;
srom_1(46131) <= 2198593;
srom_1(46132) <= 2600572;
srom_1(46133) <= 3029692;
srom_1(46134) <= 3483942;
srom_1(46135) <= 3961192;
srom_1(46136) <= 4459203;
srom_1(46137) <= 4975641;
srom_1(46138) <= 5508083;
srom_1(46139) <= 6054033;
srom_1(46140) <= 6610930;
srom_1(46141) <= 7176164;
srom_1(46142) <= 7747084;
srom_1(46143) <= 8321011;
srom_1(46144) <= 8895256;
srom_1(46145) <= 9467125;
srom_1(46146) <= 10033936;
srom_1(46147) <= 10593031;
srom_1(46148) <= 11141790;
srom_1(46149) <= 11677638;
srom_1(46150) <= 12198062;
srom_1(46151) <= 12700623;
srom_1(46152) <= 13182963;
srom_1(46153) <= 13642820;
srom_1(46154) <= 14078039;
srom_1(46155) <= 14486578;
srom_1(46156) <= 14866522;
srom_1(46157) <= 15216088;
srom_1(46158) <= 15533638;
srom_1(46159) <= 15817683;
srom_1(46160) <= 16066890;
srom_1(46161) <= 16280091;
srom_1(46162) <= 16456286;
srom_1(46163) <= 16594649;
srom_1(46164) <= 16694531;
srom_1(46165) <= 16755464;
srom_1(46166) <= 16777161;
srom_1(46167) <= 16759522;
srom_1(46168) <= 16702629;
srom_1(46169) <= 16606748;
srom_1(46170) <= 16472330;
srom_1(46171) <= 16300004;
srom_1(46172) <= 16090579;
srom_1(46173) <= 15845037;
srom_1(46174) <= 15564529;
srom_1(46175) <= 15250371;
srom_1(46176) <= 14904035;
srom_1(46177) <= 14527147;
srom_1(46178) <= 14121473;
srom_1(46179) <= 13688915;
srom_1(46180) <= 13231502;
srom_1(46181) <= 12751380;
srom_1(46182) <= 12250799;
srom_1(46183) <= 11732106;
srom_1(46184) <= 11197735;
srom_1(46185) <= 10650191;
srom_1(46186) <= 10092042;
srom_1(46187) <= 9525904;
srom_1(46188) <= 8954434;
srom_1(46189) <= 8380310;
srom_1(46190) <= 7806225;
srom_1(46191) <= 7234871;
srom_1(46192) <= 6668927;
srom_1(46193) <= 6111047;
srom_1(46194) <= 5563848;
srom_1(46195) <= 5029895;
srom_1(46196) <= 4511692;
srom_1(46197) <= 4011669;
srom_1(46198) <= 3532171;
srom_1(46199) <= 3075447;
srom_1(46200) <= 2643638;
srom_1(46201) <= 2238769;
srom_1(46202) <= 1862739;
srom_1(46203) <= 1517311;
srom_1(46204) <= 1204104;
srom_1(46205) <= 924589;
srom_1(46206) <= 680074;
srom_1(46207) <= 471708;
srom_1(46208) <= 300466;
srom_1(46209) <= 167153;
srom_1(46210) <= 72393;
srom_1(46211) <= 16630;
srom_1(46212) <= 127;
srom_1(46213) <= 22960;
srom_1(46214) <= 85022;
srom_1(46215) <= 186023;
srom_1(46216) <= 325489;
srom_1(46217) <= 502765;
srom_1(46218) <= 717021;
srom_1(46219) <= 967251;
srom_1(46220) <= 1252283;
srom_1(46221) <= 1570779;
srom_1(46222) <= 1921246;
srom_1(46223) <= 2302041;
srom_1(46224) <= 2711379;
srom_1(46225) <= 3147338;
srom_1(46226) <= 3607876;
srom_1(46227) <= 4090832;
srom_1(46228) <= 4593942;
srom_1(46229) <= 5114846;
srom_1(46230) <= 5651103;
srom_1(46231) <= 6200196;
srom_1(46232) <= 6759551;
srom_1(46233) <= 7326546;
srom_1(46234) <= 7898521;
srom_1(46235) <= 8472794;
srom_1(46236) <= 9046673;
srom_1(46237) <= 9617465;
srom_1(46238) <= 10182496;
srom_1(46239) <= 10739113;
srom_1(46240) <= 11284709;
srom_1(46241) <= 11816724;
srom_1(46242) <= 12332663;
srom_1(46243) <= 12830107;
srom_1(46244) <= 13306723;
srom_1(46245) <= 13760277;
srom_1(46246) <= 14188641;
srom_1(46247) <= 14589806;
srom_1(46248) <= 14961892;
srom_1(46249) <= 15303154;
srom_1(46250) <= 15611991;
srom_1(46251) <= 15886955;
srom_1(46252) <= 16126757;
srom_1(46253) <= 16330272;
srom_1(46254) <= 16496545;
srom_1(46255) <= 16624798;
srom_1(46256) <= 16714429;
srom_1(46257) <= 16765016;
srom_1(46258) <= 16776324;
srom_1(46259) <= 16748299;
srom_1(46260) <= 16681073;
srom_1(46261) <= 16574960;
srom_1(46262) <= 16430459;
srom_1(46263) <= 16248247;
srom_1(46264) <= 16029178;
srom_1(46265) <= 15774280;
srom_1(46266) <= 15484748;
srom_1(46267) <= 15161939;
srom_1(46268) <= 14807369;
srom_1(46269) <= 14422698;
srom_1(46270) <= 14009732;
srom_1(46271) <= 13570406;
srom_1(46272) <= 13106781;
srom_1(46273) <= 12621030;
srom_1(46274) <= 12115433;
srom_1(46275) <= 11592359;
srom_1(46276) <= 11054261;
srom_1(46277) <= 10503664;
srom_1(46278) <= 9943148;
srom_1(46279) <= 9375342;
srom_1(46280) <= 8802910;
srom_1(46281) <= 8228534;
srom_1(46282) <= 7654909;
srom_1(46283) <= 7084725;
srom_1(46284) <= 6520655;
srom_1(46285) <= 5965344;
srom_1(46286) <= 5421397;
srom_1(46287) <= 4891364;
srom_1(46288) <= 4377731;
srom_1(46289) <= 3882907;
srom_1(46290) <= 3409211;
srom_1(46291) <= 2958865;
srom_1(46292) <= 2533981;
srom_1(46293) <= 2136552;
srom_1(46294) <= 1768440;
srom_1(46295) <= 1431373;
srom_1(46296) <= 1126931;
srom_1(46297) <= 856541;
srom_1(46298) <= 621472;
srom_1(46299) <= 422825;
srom_1(46300) <= 261532;
srom_1(46301) <= 138351;
srom_1(46302) <= 53857;
srom_1(46303) <= 8448;
srom_1(46304) <= 2337;
srom_1(46305) <= 35551;
srom_1(46306) <= 107936;
srom_1(46307) <= 219152;
srom_1(46308) <= 368677;
srom_1(46309) <= 555811;
srom_1(46310) <= 779675;
srom_1(46311) <= 1039220;
srom_1(46312) <= 1333229;
srom_1(46313) <= 1660323;
srom_1(46314) <= 2018968;
srom_1(46315) <= 2407482;
srom_1(46316) <= 2824044;
srom_1(46317) <= 3266700;
srom_1(46318) <= 3733375;
srom_1(46319) <= 4221880;
srom_1(46320) <= 4729923;
srom_1(46321) <= 5255124;
srom_1(46322) <= 5795019;
srom_1(46323) <= 6347075;
srom_1(46324) <= 6908706;
srom_1(46325) <= 7477276;
srom_1(46326) <= 8050119;
srom_1(46327) <= 8624550;
srom_1(46328) <= 9197875;
srom_1(46329) <= 9767404;
srom_1(46330) <= 10330468;
srom_1(46331) <= 10884426;
srom_1(46332) <= 11426680;
srom_1(46333) <= 11954687;
srom_1(46334) <= 12465972;
srom_1(46335) <= 12958137;
srom_1(46336) <= 13428873;
srom_1(46337) <= 13875974;
srom_1(46338) <= 14297343;
srom_1(46339) <= 14691004;
srom_1(46340) <= 15055111;
srom_1(46341) <= 15387956;
srom_1(46342) <= 15687979;
srom_1(46343) <= 15953772;
srom_1(46344) <= 16184090;
srom_1(46345) <= 16377853;
srom_1(46346) <= 16534150;
srom_1(46347) <= 16652251;
srom_1(46348) <= 16731601;
srom_1(46349) <= 16771827;
srom_1(46350) <= 16772742;
srom_1(46351) <= 16734340;
srom_1(46352) <= 16656803;
srom_1(46353) <= 16540493;
srom_1(46354) <= 16385956;
srom_1(46355) <= 16193916;
srom_1(46356) <= 15965275;
srom_1(46357) <= 15701105;
srom_1(46358) <= 15402643;
srom_1(46359) <= 15071291;
srom_1(46360) <= 14708601;
srom_1(46361) <= 14316274;
srom_1(46362) <= 13896150;
srom_1(46363) <= 13450200;
srom_1(46364) <= 12980514;
srom_1(46365) <= 12489295;
srom_1(46366) <= 11978847;
srom_1(46367) <= 11451563;
srom_1(46368) <= 10909915;
srom_1(46369) <= 10356444;
srom_1(46370) <= 9793745;
srom_1(46371) <= 9224457;
srom_1(46372) <= 8651250;
srom_1(46373) <= 8076811;
srom_1(46374) <= 7503834;
srom_1(46375) <= 6935006;
srom_1(46376) <= 6372994;
srom_1(46377) <= 5820435;
srom_1(46378) <= 5279918;
srom_1(46379) <= 4753979;
srom_1(46380) <= 4245084;
srom_1(46381) <= 3755620;
srom_1(46382) <= 3287881;
srom_1(46383) <= 2844061;
srom_1(46384) <= 2426242;
srom_1(46385) <= 2036382;
srom_1(46386) <= 1676309;
srom_1(46387) <= 1347714;
srom_1(46388) <= 1052135;
srom_1(46389) <= 790959;
srom_1(46390) <= 565412;
srom_1(46391) <= 376550;
srom_1(46392) <= 225259;
srom_1(46393) <= 112250;
srom_1(46394) <= 38050;
srom_1(46395) <= 3010;
srom_1(46396) <= 7292;
srom_1(46397) <= 50878;
srom_1(46398) <= 133561;
srom_1(46399) <= 254956;
srom_1(46400) <= 414492;
srom_1(46401) <= 611421;
srom_1(46402) <= 844820;
srom_1(46403) <= 1113595;
srom_1(46404) <= 1416485;
srom_1(46405) <= 1752069;
srom_1(46406) <= 2118774;
srom_1(46407) <= 2514881;
srom_1(46408) <= 2938532;
srom_1(46409) <= 3387740;
srom_1(46410) <= 3860398;
srom_1(46411) <= 4354291;
srom_1(46412) <= 4867103;
srom_1(46413) <= 5396428;
srom_1(46414) <= 5939784;
srom_1(46415) <= 6494623;
srom_1(46416) <= 7058345;
srom_1(46417) <= 7628304;
srom_1(46418) <= 8201828;
srom_1(46419) <= 8776229;
srom_1(46420) <= 9348811;
srom_1(46421) <= 9916891;
srom_1(46422) <= 10477805;
srom_1(46423) <= 11028921;
srom_1(46424) <= 11567656;
srom_1(46425) <= 12091483;
srom_1(46426) <= 12597947;
srom_1(46427) <= 13084671;
srom_1(46428) <= 13549374;
srom_1(46429) <= 13989876;
srom_1(46430) <= 14404112;
srom_1(46431) <= 14790139;
srom_1(46432) <= 15146147;
srom_1(46433) <= 15470467;
srom_1(46434) <= 15761577;
srom_1(46435) <= 16018113;
srom_1(46436) <= 16238872;
srom_1(46437) <= 16422818;
srom_1(46438) <= 16569089;
srom_1(46439) <= 16676998;
srom_1(46440) <= 16746041;
srom_1(46441) <= 16775893;
srom_1(46442) <= 16766414;
srom_1(46443) <= 16717648;
srom_1(46444) <= 16629825;
srom_1(46445) <= 16503356;
srom_1(46446) <= 16338834;
srom_1(46447) <= 16137031;
srom_1(46448) <= 15898892;
srom_1(46449) <= 15625536;
srom_1(46450) <= 15318243;
srom_1(46451) <= 14978454;
srom_1(46452) <= 14607764;
srom_1(46453) <= 14207909;
srom_1(46454) <= 13780766;
srom_1(46455) <= 13328337;
srom_1(46456) <= 12852744;
srom_1(46457) <= 12356218;
srom_1(46458) <= 11841085;
srom_1(46459) <= 11309763;
srom_1(46460) <= 10764743;
srom_1(46461) <= 10208580;
srom_1(46462) <= 9643883;
srom_1(46463) <= 9073299;
srom_1(46464) <= 8499504;
srom_1(46465) <= 7925190;
srom_1(46466) <= 7353048;
srom_1(46467) <= 6785763;
srom_1(46468) <= 6225994;
srom_1(46469) <= 5676366;
srom_1(46470) <= 5139456;
srom_1(46471) <= 4617784;
srom_1(46472) <= 4113793;
srom_1(46473) <= 3629849;
srom_1(46474) <= 3168221;
srom_1(46475) <= 2731072;
srom_1(46476) <= 2320454;
srom_1(46477) <= 1938291;
srom_1(46478) <= 1586376;
srom_1(46479) <= 1266359;
srom_1(46480) <= 979741;
srom_1(46481) <= 727865;
srom_1(46482) <= 511913;
srom_1(46483) <= 332898;
srom_1(46484) <= 191659;
srom_1(46485) <= 88858;
srom_1(46486) <= 24977;
srom_1(46487) <= 317;
srom_1(46488) <= 14992;
srom_1(46489) <= 68933;
srom_1(46490) <= 161889;
srom_1(46491) <= 293422;
srom_1(46492) <= 462917;
srom_1(46493) <= 669578;
srom_1(46494) <= 912436;
srom_1(46495) <= 1190352;
srom_1(46496) <= 1502023;
srom_1(46497) <= 1845988;
srom_1(46498) <= 2220634;
srom_1(46499) <= 2624203;
srom_1(46500) <= 3054804;
srom_1(46501) <= 3510416;
srom_1(46502) <= 3988904;
srom_1(46503) <= 4488024;
srom_1(46504) <= 5005435;
srom_1(46505) <= 5538711;
srom_1(46506) <= 6085351;
srom_1(46507) <= 6642791;
srom_1(46508) <= 7208419;
srom_1(46509) <= 7779581;
srom_1(46510) <= 8353598;
srom_1(46511) <= 8927780;
srom_1(46512) <= 9499434;
srom_1(46513) <= 10065878;
srom_1(46514) <= 10624457;
srom_1(46515) <= 11172552;
srom_1(46516) <= 11707591;
srom_1(46517) <= 12227067;
srom_1(46518) <= 12728543;
srom_1(46519) <= 13209667;
srom_1(46520) <= 13668184;
srom_1(46521) <= 14101943;
srom_1(46522) <= 14508910;
srom_1(46523) <= 14887177;
srom_1(46524) <= 15234970;
srom_1(46525) <= 15550658;
srom_1(46526) <= 15832761;
srom_1(46527) <= 16079956;
srom_1(46528) <= 16291083;
srom_1(46529) <= 16465153;
srom_1(46530) <= 16601349;
srom_1(46531) <= 16699032;
srom_1(46532) <= 16757746;
srom_1(46533) <= 16777213;
srom_1(46534) <= 16757343;
srom_1(46535) <= 16698230;
srom_1(46536) <= 16600150;
srom_1(46537) <= 16463563;
srom_1(46538) <= 16289110;
srom_1(46539) <= 16077608;
srom_1(46540) <= 15830051;
srom_1(46541) <= 15547597;
srom_1(46542) <= 15231573;
srom_1(46543) <= 14883460;
srom_1(46544) <= 14504890;
srom_1(46545) <= 14097639;
srom_1(46546) <= 13663616;
srom_1(46547) <= 13204857;
srom_1(46548) <= 12723513;
srom_1(46549) <= 12221841;
srom_1(46550) <= 11702194;
srom_1(46551) <= 11167008;
srom_1(46552) <= 10618793;
srom_1(46553) <= 10060120;
srom_1(46554) <= 9493609;
srom_1(46555) <= 8921916;
srom_1(46556) <= 8347722;
srom_1(46557) <= 7773720;
srom_1(46558) <= 7202601;
srom_1(46559) <= 6637044;
srom_1(46560) <= 6079701;
srom_1(46561) <= 5533185;
srom_1(46562) <= 5000059;
srom_1(46563) <= 4482823;
srom_1(46564) <= 3983902;
srom_1(46565) <= 3505637;
srom_1(46566) <= 3050269;
srom_1(46567) <= 2619935;
srom_1(46568) <= 2216652;
srom_1(46569) <= 1842312;
srom_1(46570) <= 1498670;
srom_1(46571) <= 1187336;
srom_1(46572) <= 909772;
srom_1(46573) <= 667279;
srom_1(46574) <= 460994;
srom_1(46575) <= 291884;
srom_1(46576) <= 160742;
srom_1(46577) <= 68184;
srom_1(46578) <= 14643;
srom_1(46579) <= 370;
srom_1(46580) <= 25433;
srom_1(46581) <= 89713;
srom_1(46582) <= 192910;
srom_1(46583) <= 334539;
srom_1(46584) <= 513937;
srom_1(46585) <= 730261;
srom_1(46586) <= 982498;
srom_1(46587) <= 1269465;
srom_1(46588) <= 1589816;
srom_1(46589) <= 1942049;
srom_1(46590) <= 2324512;
srom_1(46591) <= 2735412;
srom_1(46592) <= 3172822;
srom_1(46593) <= 3634690;
srom_1(46594) <= 4118850;
srom_1(46595) <= 4623034;
srom_1(46596) <= 5144875;
srom_1(46597) <= 5681927;
srom_1(46598) <= 6231672;
srom_1(46599) <= 6791531;
srom_1(46600) <= 7358880;
srom_1(46601) <= 7931057;
srom_1(46602) <= 8505380;
srom_1(46603) <= 9079155;
srom_1(46604) <= 9649692;
srom_1(46605) <= 10214316;
srom_1(46606) <= 10770378;
srom_1(46607) <= 11315271;
srom_1(46608) <= 11846440;
srom_1(46609) <= 12361394;
srom_1(46610) <= 12857718;
srom_1(46611) <= 13333085;
srom_1(46612) <= 13785266;
srom_1(46613) <= 14212140;
srom_1(46614) <= 14611705;
srom_1(46615) <= 14982089;
srom_1(46616) <= 15321553;
srom_1(46617) <= 15628506;
srom_1(46618) <= 15901508;
srom_1(46619) <= 16139280;
srom_1(46620) <= 16340707;
srom_1(46621) <= 16504843;
srom_1(46622) <= 16630920;
srom_1(46623) <= 16718345;
srom_1(46624) <= 16766710;
srom_1(46625) <= 16775787;
srom_1(46626) <= 16745533;
srom_1(46627) <= 16676091;
srom_1(46628) <= 16567786;
srom_1(46629) <= 16421126;
srom_1(46630) <= 16236799;
srom_1(46631) <= 16015668;
srom_1(46632) <= 15758772;
srom_1(46633) <= 15467315;
srom_1(46634) <= 15142663;
srom_1(46635) <= 14786340;
srom_1(46636) <= 14400015;
srom_1(46637) <= 13985500;
srom_1(46638) <= 13544740;
srom_1(46639) <= 13079800;
srom_1(46640) <= 12592863;
srom_1(46641) <= 12086210;
srom_1(46642) <= 11562217;
srom_1(46643) <= 11023343;
srom_1(46644) <= 10472113;
srom_1(46645) <= 9911113;
srom_1(46646) <= 9342973;
srom_1(46647) <= 8770359;
srom_1(46648) <= 8195954;
srom_1(46649) <= 7622452;
srom_1(46650) <= 7052543;
srom_1(46651) <= 6488899;
srom_1(46652) <= 5934164;
srom_1(46653) <= 5390939;
srom_1(46654) <= 4861770;
srom_1(46655) <= 4349140;
srom_1(46656) <= 3855453;
srom_1(46657) <= 3383023;
srom_1(46658) <= 2934066;
srom_1(46659) <= 2510687;
srom_1(46660) <= 2114872;
srom_1(46661) <= 1748476;
srom_1(46662) <= 1413219;
srom_1(46663) <= 1110671;
srom_1(46664) <= 842252;
srom_1(46665) <= 609221;
srom_1(46666) <= 412669;
srom_1(46667) <= 253520;
srom_1(46668) <= 132519;
srom_1(46669) <= 50233;
srom_1(46670) <= 7049;
srom_1(46671) <= 3169;
srom_1(46672) <= 38611;
srom_1(46673) <= 113210;
srom_1(46674) <= 226614;
srom_1(46675) <= 378293;
srom_1(46676) <= 567535;
srom_1(46677) <= 793452;
srom_1(46678) <= 1054986;
srom_1(46679) <= 1350910;
srom_1(46680) <= 1679836;
srom_1(46681) <= 2040221;
srom_1(46682) <= 2430376;
srom_1(46683) <= 2848472;
srom_1(46684) <= 3292547;
srom_1(46685) <= 3760519;
srom_1(46686) <= 4250195;
srom_1(46687) <= 4759276;
srom_1(46688) <= 5285377;
srom_1(46689) <= 5826029;
srom_1(46690) <= 6378699;
srom_1(46691) <= 6940794;
srom_1(46692) <= 7509678;
srom_1(46693) <= 8082683;
srom_1(46694) <= 8657123;
srom_1(46695) <= 9230304;
srom_1(46696) <= 9799538;
srom_1(46697) <= 10362156;
srom_1(46698) <= 10915519;
srom_1(46699) <= 11457032;
srom_1(46700) <= 11984157;
srom_1(46701) <= 12494421;
srom_1(46702) <= 12985431;
srom_1(46703) <= 13454885;
srom_1(46704) <= 13900581;
srom_1(46705) <= 14320430;
srom_1(46706) <= 14712463;
srom_1(46707) <= 15074841;
srom_1(46708) <= 15405865;
srom_1(46709) <= 15703982;
srom_1(46710) <= 15967796;
srom_1(46711) <= 16196068;
srom_1(46712) <= 16387727;
srom_1(46713) <= 16541877;
srom_1(46714) <= 16657793;
srom_1(46715) <= 16734931;
srom_1(46716) <= 16772931;
srom_1(46717) <= 16771614;
srom_1(46718) <= 16730987;
srom_1(46719) <= 16651239;
srom_1(46720) <= 16532744;
srom_1(46721) <= 16376059;
srom_1(46722) <= 16181918;
srom_1(46723) <= 15951232;
srom_1(46724) <= 15685081;
srom_1(46725) <= 15384716;
srom_1(46726) <= 15051542;
srom_1(46727) <= 14687125;
srom_1(46728) <= 14293171;
srom_1(46729) <= 13871528;
srom_1(46730) <= 13424175;
srom_1(46731) <= 12953208;
srom_1(46732) <= 12460836;
srom_1(46733) <= 11949367;
srom_1(46734) <= 11421202;
srom_1(46735) <= 10878815;
srom_1(46736) <= 10324751;
srom_1(46737) <= 9761607;
srom_1(46738) <= 9192026;
srom_1(46739) <= 8618676;
srom_1(46740) <= 8044248;
srom_1(46741) <= 7471435;
srom_1(46742) <= 6902922;
srom_1(46743) <= 6341376;
srom_1(46744) <= 5789431;
srom_1(46745) <= 5249674;
srom_1(46746) <= 4724636;
srom_1(46747) <= 4216781;
srom_1(46748) <= 3728488;
srom_1(46749) <= 3262048;
srom_1(46750) <= 2819648;
srom_1(46751) <= 2403363;
srom_1(46752) <= 2015145;
srom_1(46753) <= 1656815;
srom_1(46754) <= 1330052;
srom_1(46755) <= 1036389;
srom_1(46756) <= 777203;
srom_1(46757) <= 553709;
srom_1(46758) <= 366956;
srom_1(46759) <= 217820;
srom_1(46760) <= 106999;
srom_1(46761) <= 35013;
srom_1(46762) <= 2200;
srom_1(46763) <= 8714;
srom_1(46764) <= 54524;
srom_1(46765) <= 139416;
srom_1(46766) <= 262990;
srom_1(46767) <= 424669;
srom_1(46768) <= 623693;
srom_1(46769) <= 859130;
srom_1(46770) <= 1129874;
srom_1(46771) <= 1434658;
srom_1(46772) <= 1772051;
srom_1(46773) <= 2140471;
srom_1(46774) <= 2538191;
srom_1(46775) <= 2963346;
srom_1(46776) <= 3413941;
srom_1(46777) <= 3887865;
srom_1(46778) <= 4382893;
srom_1(46779) <= 4896707;
srom_1(46780) <= 5426894;
srom_1(46781) <= 5970971;
srom_1(46782) <= 6526384;
srom_1(46783) <= 7090530;
srom_1(46784) <= 7660763;
srom_1(46785) <= 8234409;
srom_1(46786) <= 8808779;
srom_1(46787) <= 9381178;
srom_1(46788) <= 9948922;
srom_1(46789) <= 10509350;
srom_1(46790) <= 11059832;
srom_1(46791) <= 11597789;
srom_1(46792) <= 12120696;
srom_1(46793) <= 12626103;
srom_1(46794) <= 13111638;
srom_1(46795) <= 13575026;
srom_1(46796) <= 14014092;
srom_1(46797) <= 14426779;
srom_1(46798) <= 14811150;
srom_1(46799) <= 15165404;
srom_1(46800) <= 15487880;
srom_1(46801) <= 15777064;
srom_1(46802) <= 16031602;
srom_1(46803) <= 16250299;
srom_1(46804) <= 16432129;
srom_1(46805) <= 16576241;
srom_1(46806) <= 16681958;
srom_1(46807) <= 16748785;
srom_1(46808) <= 16776408;
srom_1(46809) <= 16764698;
srom_1(46810) <= 16713709;
srom_1(46811) <= 16623681;
srom_1(46812) <= 16495036;
srom_1(46813) <= 16328377;
srom_1(46814) <= 16124486;
srom_1(46815) <= 15884319;
srom_1(46816) <= 15609002;
srom_1(46817) <= 15299825;
srom_1(46818) <= 14958240;
srom_1(46819) <= 14585847;
srom_1(46820) <= 14184394;
srom_1(46821) <= 13755762;
srom_1(46822) <= 13301962;
srom_1(46823) <= 12825121;
srom_1(46824) <= 12327475;
srom_1(46825) <= 11811360;
srom_1(46826) <= 11279193;
srom_1(46827) <= 10733472;
srom_1(46828) <= 10176755;
srom_1(46829) <= 9611652;
srom_1(46830) <= 9040815;
srom_1(46831) <= 8466918;
srom_1(46832) <= 7892655;
srom_1(46833) <= 7320717;
srom_1(46834) <= 6753787;
srom_1(46835) <= 6194524;
srom_1(46836) <= 5645549;
srom_1(46837) <= 5109437;
srom_1(46838) <= 4588702;
srom_1(46839) <= 4085787;
srom_1(46840) <= 3603048;
srom_1(46841) <= 3142751;
srom_1(46842) <= 2707054;
srom_1(46843) <= 2297999;
srom_1(46844) <= 1917506;
srom_1(46845) <= 1567357;
srom_1(46846) <= 1249196;
srom_1(46847) <= 964513;
srom_1(46848) <= 714645;
srom_1(46849) <= 500763;
srom_1(46850) <= 323870;
srom_1(46851) <= 184795;
srom_1(46852) <= 84190;
srom_1(46853) <= 22528;
srom_1(46854) <= 97;
srom_1(46855) <= 17002;
srom_1(46856) <= 73165;
srom_1(46857) <= 168322;
srom_1(46858) <= 302027;
srom_1(46859) <= 473652;
srom_1(46860) <= 682394;
srom_1(46861) <= 927272;
srom_1(46862) <= 1207139;
srom_1(46863) <= 1520683;
srom_1(46864) <= 1866433;
srom_1(46865) <= 2242767;
srom_1(46866) <= 2647921;
srom_1(46867) <= 3079996;
srom_1(46868) <= 3536964;
srom_1(46869) <= 4016683;
srom_1(46870) <= 4516904;
srom_1(46871) <= 5035280;
srom_1(46872) <= 5569382;
srom_1(46873) <= 6116703;
srom_1(46874) <= 6674679;
srom_1(46875) <= 7240691;
srom_1(46876) <= 7812087;
srom_1(46877) <= 8386186;
srom_1(46878) <= 8960297;
srom_1(46879) <= 9531726;
srom_1(46880) <= 10097795;
srom_1(46881) <= 10655849;
srom_1(46882) <= 11203272;
srom_1(46883) <= 11737495;
srom_1(46884) <= 12256014;
srom_1(46885) <= 12756398;
srom_1(46886) <= 13236299;
srom_1(46887) <= 13693468;
srom_1(46888) <= 14125761;
srom_1(46889) <= 14531150;
srom_1(46890) <= 14907735;
srom_1(46891) <= 15253749;
srom_1(46892) <= 15567571;
srom_1(46893) <= 15847727;
srom_1(46894) <= 16092906;
srom_1(46895) <= 16301956;
srom_1(46896) <= 16473897;
srom_1(46897) <= 16607925;
srom_1(46898) <= 16703408;
srom_1(46899) <= 16759901;
srom_1(46900) <= 16777138;
srom_1(46901) <= 16755039;
srom_1(46902) <= 16693706;
srom_1(46903) <= 16593428;
srom_1(46904) <= 16454674;
srom_1(46905) <= 16278096;
srom_1(46906) <= 16064522;
srom_1(46907) <= 15814952;
srom_1(46908) <= 15530558;
srom_1(46909) <= 15212672;
srom_1(46910) <= 14862787;
srom_1(46911) <= 14482541;
srom_1(46912) <= 14073720;
srom_1(46913) <= 13638238;
srom_1(46914) <= 13178140;
srom_1(46915) <= 12695581;
srom_1(46916) <= 12192826;
srom_1(46917) <= 11672231;
srom_1(46918) <= 11136238;
srom_1(46919) <= 10587361;
srom_1(46920) <= 10028173;
srom_1(46921) <= 9461297;
srom_1(46922) <= 8889390;
srom_1(46923) <= 8315135;
srom_1(46924) <= 7741225;
srom_1(46925) <= 7170350;
srom_1(46926) <= 6605188;
srom_1(46927) <= 6048389;
srom_1(46928) <= 5502565;
srom_1(46929) <= 4970273;
srom_1(46930) <= 4454012;
srom_1(46931) <= 3956201;
srom_1(46932) <= 3479176;
srom_1(46933) <= 3025172;
srom_1(46934) <= 2596320;
srom_1(46935) <= 2194629;
srom_1(46936) <= 1821984;
srom_1(46937) <= 1480132;
srom_1(46938) <= 1170677;
srom_1(46939) <= 895069;
srom_1(46940) <= 654600;
srom_1(46941) <= 450399;
srom_1(46942) <= 283423;
srom_1(46943) <= 154455;
srom_1(46944) <= 64100;
srom_1(46945) <= 12781;
srom_1(46946) <= 739;
srom_1(46947) <= 28031;
srom_1(46948) <= 94529;
srom_1(46949) <= 199920;
srom_1(46950) <= 343711;
srom_1(46951) <= 525227;
srom_1(46952) <= 743617;
srom_1(46953) <= 997858;
srom_1(46954) <= 1286756;
srom_1(46955) <= 1608957;
srom_1(46956) <= 1962950;
srom_1(46957) <= 2347075;
srom_1(46958) <= 2759531;
srom_1(46959) <= 3198384;
srom_1(46960) <= 3661575;
srom_1(46961) <= 4146933;
srom_1(46962) <= 4652182;
srom_1(46963) <= 5174952;
srom_1(46964) <= 5712792;
srom_1(46965) <= 6263180;
srom_1(46966) <= 6823535;
srom_1(46967) <= 7391229;
srom_1(46968) <= 7963600;
srom_1(46969) <= 8537964;
srom_1(46970) <= 9111627;
srom_1(46971) <= 9681900;
srom_1(46972) <= 10246109;
srom_1(46973) <= 10801607;
srom_1(46974) <= 11345789;
srom_1(46975) <= 11876104;
srom_1(46976) <= 12390066;
srom_1(46977) <= 12885263;
srom_1(46978) <= 13359373;
srom_1(46979) <= 13810174;
srom_1(46980) <= 14235552;
srom_1(46981) <= 14633511;
srom_1(46982) <= 15002185;
srom_1(46983) <= 15339846;
srom_1(46984) <= 15644911;
srom_1(46985) <= 15915948;
srom_1(46986) <= 16151687;
srom_1(46987) <= 16351022;
srom_1(46988) <= 16513019;
srom_1(46989) <= 16636917;
srom_1(46990) <= 16722136;
srom_1(46991) <= 16768277;
srom_1(46992) <= 16775122;
srom_1(46993) <= 16742640;
srom_1(46994) <= 16670984;
srom_1(46995) <= 16560488;
srom_1(46996) <= 16411671;
srom_1(46997) <= 16225232;
srom_1(46998) <= 16002044;
srom_1(46999) <= 15743154;
srom_1(47000) <= 15449776;
srom_1(47001) <= 15123285;
srom_1(47002) <= 14765214;
srom_1(47003) <= 14377240;
srom_1(47004) <= 13961184;
srom_1(47005) <= 13518996;
srom_1(47006) <= 13052749;
srom_1(47007) <= 12564631;
srom_1(47008) <= 12056931;
srom_1(47009) <= 11532028;
srom_1(47010) <= 10992384;
srom_1(47011) <= 10440531;
srom_1(47012) <= 9879055;
srom_1(47013) <= 9310590;
srom_1(47014) <= 8737802;
srom_1(47015) <= 8163376;
srom_1(47016) <= 7590006;
srom_1(47017) <= 7020381;
srom_1(47018) <= 6457173;
srom_1(47019) <= 5903021;
srom_1(47020) <= 5360525;
srom_1(47021) <= 4832229;
srom_1(47022) <= 4320610;
srom_1(47023) <= 3828067;
srom_1(47024) <= 3356911;
srom_1(47025) <= 2909349;
srom_1(47026) <= 2487482;
srom_1(47027) <= 2093287;
srom_1(47028) <= 1728613;
srom_1(47029) <= 1395170;
srom_1(47030) <= 1094521;
srom_1(47031) <= 828077;
srom_1(47032) <= 597087;
srom_1(47033) <= 402634;
srom_1(47034) <= 245630;
srom_1(47035) <= 126812;
srom_1(47036) <= 46735;
srom_1(47037) <= 5777;
srom_1(47038) <= 4128;
srom_1(47039) <= 41798;
srom_1(47040) <= 118608;
srom_1(47041) <= 234199;
srom_1(47042) <= 388029;
srom_1(47043) <= 579376;
srom_1(47044) <= 807344;
srom_1(47045) <= 1070863;
srom_1(47046) <= 1368697;
srom_1(47047) <= 1699450;
srom_1(47048) <= 2061570;
srom_1(47049) <= 2453361;
srom_1(47050) <= 2872983;
srom_1(47051) <= 3318471;
srom_1(47052) <= 3787734;
srom_1(47053) <= 4278572;
srom_1(47054) <= 4788683;
srom_1(47055) <= 5315676;
srom_1(47056) <= 5857079;
srom_1(47057) <= 6410353;
srom_1(47058) <= 6972903;
srom_1(47059) <= 7542093;
srom_1(47060) <= 8115251;
srom_1(47061) <= 8689692;
srom_1(47062) <= 9262721;
srom_1(47063) <= 9831651;
srom_1(47064) <= 10393814;
srom_1(47065) <= 10946574;
srom_1(47066) <= 11487339;
srom_1(47067) <= 12013572;
srom_1(47068) <= 12522807;
srom_1(47069) <= 13012655;
srom_1(47070) <= 13480820;
srom_1(47071) <= 13925105;
srom_1(47072) <= 14343428;
srom_1(47073) <= 14733827;
srom_1(47074) <= 15094470;
srom_1(47075) <= 15423668;
srom_1(47076) <= 15719876;
srom_1(47077) <= 15981705;
srom_1(47078) <= 16207927;
srom_1(47079) <= 16397482;
srom_1(47080) <= 16549480;
srom_1(47081) <= 16663209;
srom_1(47082) <= 16738136;
srom_1(47083) <= 16773909;
srom_1(47084) <= 16770361;
srom_1(47085) <= 16727507;
srom_1(47086) <= 16645550;
srom_1(47087) <= 16524873;
srom_1(47088) <= 16366042;
srom_1(47089) <= 16169802;
srom_1(47090) <= 15937074;
srom_1(47091) <= 15668948;
srom_1(47092) <= 15366682;
srom_1(47093) <= 15031694;
srom_1(47094) <= 14665553;
srom_1(47095) <= 14269979;
srom_1(47096) <= 13846824;
srom_1(47097) <= 13398074;
srom_1(47098) <= 12925832;
srom_1(47099) <= 12432315;
srom_1(47100) <= 11919834;
srom_1(47101) <= 11390795;
srom_1(47102) <= 10847677;
srom_1(47103) <= 10293028;
srom_1(47104) <= 9729449;
srom_1(47105) <= 9159582;
srom_1(47106) <= 8586099;
srom_1(47107) <= 8011690;
srom_1(47108) <= 7439049;
srom_1(47109) <= 6870861;
srom_1(47110) <= 6309789;
srom_1(47111) <= 5758467;
srom_1(47112) <= 5219477;
srom_1(47113) <= 4695349;
srom_1(47114) <= 4188540;
srom_1(47115) <= 3701426;
srom_1(47116) <= 3236293;
srom_1(47117) <= 2795320;
srom_1(47118) <= 2380576;
srom_1(47119) <= 1994005;
srom_1(47120) <= 1637422;
srom_1(47121) <= 1312496;
srom_1(47122) <= 1020754;
srom_1(47123) <= 763561;
srom_1(47124) <= 542125;
srom_1(47125) <= 357484;
srom_1(47126) <= 210503;
srom_1(47127) <= 101873;
srom_1(47128) <= 32102;
srom_1(47129) <= 1517;
srom_1(47130) <= 10262;
srom_1(47131) <= 58296;
srom_1(47132) <= 145394;
srom_1(47133) <= 271148;
srom_1(47134) <= 434966;
srom_1(47135) <= 636082;
srom_1(47136) <= 873553;
srom_1(47137) <= 1146264;
srom_1(47138) <= 1452936;
srom_1(47139) <= 1792133;
srom_1(47140) <= 2162263;
srom_1(47141) <= 2561590;
srom_1(47142) <= 2988242;
srom_1(47143) <= 3440218;
srom_1(47144) <= 3915399;
srom_1(47145) <= 4411556;
srom_1(47146) <= 4926363;
srom_1(47147) <= 5457406;
srom_1(47148) <= 6002194;
srom_1(47149) <= 6558173;
srom_1(47150) <= 7122735;
srom_1(47151) <= 7693233;
srom_1(47152) <= 8266993;
srom_1(47153) <= 8841322;
srom_1(47154) <= 9413529;
srom_1(47155) <= 9980929;
srom_1(47156) <= 10540863;
srom_1(47157) <= 11090704;
srom_1(47158) <= 11627873;
srom_1(47159) <= 12149853;
srom_1(47160) <= 12654195;
srom_1(47161) <= 13138534;
srom_1(47162) <= 13600599;
srom_1(47163) <= 14038224;
srom_1(47164) <= 14449355;
srom_1(47165) <= 14832065;
srom_1(47166) <= 15184560;
srom_1(47167) <= 15505186;
srom_1(47168) <= 15792440;
srom_1(47169) <= 16044975;
srom_1(47170) <= 16261607;
srom_1(47171) <= 16441319;
srom_1(47172) <= 16583270;
srom_1(47173) <= 16686793;
srom_1(47174) <= 16751402;
srom_1(47175) <= 16776796;
srom_1(47176) <= 16762855;
srom_1(47177) <= 16709644;
srom_1(47178) <= 16617413;
srom_1(47179) <= 16486594;
srom_1(47180) <= 16317801;
srom_1(47181) <= 16111825;
srom_1(47182) <= 15869632;
srom_1(47183) <= 15592358;
srom_1(47184) <= 15281304;
srom_1(47185) <= 14937927;
srom_1(47186) <= 14563838;
srom_1(47187) <= 14160791;
srom_1(47188) <= 13730677;
srom_1(47189) <= 13275512;
srom_1(47190) <= 12797430;
srom_1(47191) <= 12298674;
srom_1(47192) <= 11781582;
srom_1(47193) <= 11248580;
srom_1(47194) <= 10702166;
srom_1(47195) <= 10144902;
srom_1(47196) <= 9579404;
srom_1(47197) <= 9008321;
srom_1(47198) <= 8434332;
srom_1(47199) <= 7860128;
srom_1(47200) <= 7288403;
srom_1(47201) <= 6721837;
srom_1(47202) <= 6163087;
srom_1(47203) <= 5614773;
srom_1(47204) <= 5079467;
srom_1(47205) <= 4559678;
srom_1(47206) <= 4057845;
srom_1(47207) <= 3576320;
srom_1(47208) <= 3117361;
srom_1(47209) <= 2683122;
srom_1(47210) <= 2275637;
srom_1(47211) <= 1896818;
srom_1(47212) <= 1548441;
srom_1(47213) <= 1232140;
srom_1(47214) <= 949398;
srom_1(47215) <= 701541;
srom_1(47216) <= 489732;
srom_1(47217) <= 314963;
srom_1(47218) <= 178054;
srom_1(47219) <= 79647;
srom_1(47220) <= 20204;
srom_1(47221) <= 3;
srom_1(47222) <= 19139;
srom_1(47223) <= 77523;
srom_1(47224) <= 174880;
srom_1(47225) <= 310754;
srom_1(47226) <= 484507;
srom_1(47227) <= 695326;
srom_1(47228) <= 942222;
srom_1(47229) <= 1224035;
srom_1(47230) <= 1539446;
srom_1(47231) <= 1886976;
srom_1(47232) <= 2264993;
srom_1(47233) <= 2671726;
srom_1(47234) <= 3105268;
srom_1(47235) <= 3563585;
srom_1(47236) <= 4044528;
srom_1(47237) <= 4545842;
srom_1(47238) <= 5065176;
srom_1(47239) <= 5600095;
srom_1(47240) <= 6148090;
srom_1(47241) <= 6706592;
srom_1(47242) <= 7272981;
srom_1(47243) <= 7844602;
srom_1(47244) <= 8418774;
srom_1(47245) <= 8992804;
srom_1(47246) <= 9564001;
srom_1(47247) <= 10129686;
srom_1(47248) <= 10687207;
srom_1(47249) <= 11233949;
srom_1(47250) <= 11767348;
srom_1(47251) <= 12284903;
srom_1(47252) <= 12784187;
srom_1(47253) <= 13262858;
srom_1(47254) <= 13718672;
srom_1(47255) <= 14149492;
srom_1(47256) <= 14553297;
srom_1(47257) <= 14928194;
srom_1(47258) <= 15272424;
srom_1(47259) <= 15584374;
srom_1(47260) <= 15862581;
srom_1(47261) <= 16105739;
srom_1(47262) <= 16312709;
srom_1(47263) <= 16482520;
srom_1(47264) <= 16614376;
srom_1(47265) <= 16707659;
srom_1(47266) <= 16761931;
srom_1(47267) <= 16776937;
srom_1(47268) <= 16752608;
srom_1(47269) <= 16689056;
srom_1(47270) <= 16586582;
srom_1(47271) <= 16445664;
srom_1(47272) <= 16266964;
srom_1(47273) <= 16051319;
srom_1(47274) <= 15799741;
srom_1(47275) <= 15513410;
srom_1(47276) <= 15193669;
srom_1(47277) <= 14842016;
srom_1(47278) <= 14460101;
srom_1(47279) <= 14049714;
srom_1(47280) <= 13612781;
srom_1(47281) <= 13151349;
srom_1(47282) <= 12667584;
srom_1(47283) <= 12163753;
srom_1(47284) <= 11642219;
srom_1(47285) <= 11105428;
srom_1(47286) <= 10555896;
srom_1(47287) <= 9996202;
srom_1(47288) <= 9428969;
srom_1(47289) <= 8856857;
srom_1(47290) <= 8282549;
srom_1(47291) <= 7708739;
srom_1(47292) <= 7138117;
srom_1(47293) <= 6573359;
srom_1(47294) <= 6017113;
srom_1(47295) <= 5471988;
srom_1(47296) <= 4940540;
srom_1(47297) <= 4425261;
srom_1(47298) <= 3928568;
srom_1(47299) <= 3452789;
srom_1(47300) <= 3000156;
srom_1(47301) <= 2572791;
srom_1(47302) <= 2172699;
srom_1(47303) <= 1801755;
srom_1(47304) <= 1461700;
srom_1(47305) <= 1154126;
srom_1(47306) <= 880478;
srom_1(47307) <= 642038;
srom_1(47308) <= 439925;
srom_1(47309) <= 275085;
srom_1(47310) <= 148293;
srom_1(47311) <= 60142;
srom_1(47312) <= 11046;
srom_1(47313) <= 1236;
srom_1(47314) <= 30756;
srom_1(47315) <= 99470;
srom_1(47316) <= 207054;
srom_1(47317) <= 353004;
srom_1(47318) <= 536636;
srom_1(47319) <= 757089;
srom_1(47320) <= 1013328;
srom_1(47321) <= 1304153;
srom_1(47322) <= 1628199;
srom_1(47323) <= 1983947;
srom_1(47324) <= 2369729;
srom_1(47325) <= 2783735;
srom_1(47326) <= 3224024;
srom_1(47327) <= 3688532;
srom_1(47328) <= 4175080;
srom_1(47329) <= 4681387;
srom_1(47330) <= 5205078;
srom_1(47331) <= 5743698;
srom_1(47332) <= 6294720;
srom_1(47333) <= 6855562;
srom_1(47334) <= 7423593;
srom_1(47335) <= 7996149;
srom_1(47336) <= 8570545;
srom_1(47337) <= 9144088;
srom_1(47338) <= 9714089;
srom_1(47339) <= 10277873;
srom_1(47340) <= 10832799;
srom_1(47341) <= 11376263;
srom_1(47342) <= 11905716;
srom_1(47343) <= 12418677;
srom_1(47344) <= 12912739;
srom_1(47345) <= 13385586;
srom_1(47346) <= 13835000;
srom_1(47347) <= 14258875;
srom_1(47348) <= 14655222;
srom_1(47349) <= 15022182;
srom_1(47350) <= 15358035;
srom_1(47351) <= 15661207;
srom_1(47352) <= 15930274;
srom_1(47353) <= 16163976;
srom_1(47354) <= 16361217;
srom_1(47355) <= 16521071;
srom_1(47356) <= 16642790;
srom_1(47357) <= 16725802;
srom_1(47358) <= 16769718;
srom_1(47359) <= 16774331;
srom_1(47360) <= 16739622;
srom_1(47361) <= 16665751;
srom_1(47362) <= 16553067;
srom_1(47363) <= 16402096;
srom_1(47364) <= 16213547;
srom_1(47365) <= 15988304;
srom_1(47366) <= 15727424;
srom_1(47367) <= 15432130;
srom_1(47368) <= 15103806;
srom_1(47369) <= 14743992;
srom_1(47370) <= 14354376;
srom_1(47371) <= 13936784;
srom_1(47372) <= 13493174;
srom_1(47373) <= 13025628;
srom_1(47374) <= 12536337;
srom_1(47375) <= 12027596;
srom_1(47376) <= 11501791;
srom_1(47377) <= 10961386;
srom_1(47378) <= 10408917;
srom_1(47379) <= 9846975;
srom_1(47380) <= 9278193;
srom_1(47381) <= 8705240;
srom_1(47382) <= 8130802;
srom_1(47383) <= 7557572;
srom_1(47384) <= 6988240;
srom_1(47385) <= 6425475;
srom_1(47386) <= 5871915;
srom_1(47387) <= 5330158;
srom_1(47388) <= 4802742;
srom_1(47389) <= 4292141;
srom_1(47390) <= 3800751;
srom_1(47391) <= 3330874;
srom_1(47392) <= 2884715;
srom_1(47393) <= 2464365;
srom_1(47394) <= 2071797;
srom_1(47395) <= 1708849;
srom_1(47396) <= 1377226;
srom_1(47397) <= 1078481;
srom_1(47398) <= 814016;
srom_1(47399) <= 585071;
srom_1(47400) <= 392720;
srom_1(47401) <= 237864;
srom_1(47402) <= 121229;
srom_1(47403) <= 43363;
srom_1(47404) <= 4631;
srom_1(47405) <= 5214;
srom_1(47406) <= 45110;
srom_1(47407) <= 124131;
srom_1(47408) <= 241907;
srom_1(47409) <= 397886;
srom_1(47410) <= 591336;
srom_1(47411) <= 821350;
srom_1(47412) <= 1086850;
srom_1(47413) <= 1386590;
srom_1(47414) <= 1719165;
srom_1(47415) <= 2083015;
srom_1(47416) <= 2476434;
srom_1(47417) <= 2897578;
srom_1(47418) <= 3344471;
srom_1(47419) <= 3815017;
srom_1(47420) <= 4307011;
srom_1(47421) <= 4818145;
srom_1(47422) <= 5346022;
srom_1(47423) <= 5888166;
srom_1(47424) <= 6442036;
srom_1(47425) <= 7005034;
srom_1(47426) <= 7574520;
srom_1(47427) <= 8147824;
srom_1(47428) <= 8722257;
srom_1(47429) <= 9295125;
srom_1(47430) <= 9863742;
srom_1(47431) <= 10425442;
srom_1(47432) <= 10977590;
srom_1(47433) <= 11517598;
srom_1(47434) <= 12042933;
srom_1(47435) <= 12551131;
srom_1(47436) <= 13039810;
srom_1(47437) <= 13506678;
srom_1(47438) <= 13949545;
srom_1(47439) <= 14366336;
srom_1(47440) <= 14755094;
srom_1(47441) <= 15113998;
srom_1(47442) <= 15441365;
srom_1(47443) <= 15735658;
srom_1(47444) <= 15995499;
srom_1(47445) <= 16219668;
srom_1(47446) <= 16407115;
srom_1(47447) <= 16556960;
srom_1(47448) <= 16668501;
srom_1(47449) <= 16741215;
srom_1(47450) <= 16774761;
srom_1(47451) <= 16768980;
srom_1(47452) <= 16723902;
srom_1(47453) <= 16639736;
srom_1(47454) <= 16516879;
srom_1(47455) <= 16355904;
srom_1(47456) <= 16157569;
srom_1(47457) <= 15922802;
srom_1(47458) <= 15652704;
srom_1(47459) <= 15348543;
srom_1(47460) <= 15011744;
srom_1(47461) <= 14643888;
srom_1(47462) <= 14246697;
srom_1(47463) <= 13822037;
srom_1(47464) <= 13371897;
srom_1(47465) <= 12898389;
srom_1(47466) <= 12403732;
srom_1(47467) <= 11890248;
srom_1(47468) <= 11360343;
srom_1(47469) <= 10816503;
srom_1(47470) <= 10261277;
srom_1(47471) <= 9697270;
srom_1(47472) <= 9127126;
srom_1(47473) <= 8553519;
srom_1(47474) <= 7979138;
srom_1(47475) <= 7406678;
srom_1(47476) <= 6838822;
srom_1(47477) <= 6278234;
srom_1(47478) <= 5727542;
srom_1(47479) <= 5189329;
srom_1(47480) <= 4666118;
srom_1(47481) <= 4160363;
srom_1(47482) <= 3674436;
srom_1(47483) <= 3210615;
srom_1(47484) <= 2771076;
srom_1(47485) <= 2357879;
srom_1(47486) <= 1972962;
srom_1(47487) <= 1618130;
srom_1(47488) <= 1295048;
srom_1(47489) <= 1005230;
srom_1(47490) <= 750035;
srom_1(47491) <= 530659;
srom_1(47492) <= 348133;
srom_1(47493) <= 203311;
srom_1(47494) <= 96872;
srom_1(47495) <= 29317;
srom_1(47496) <= 960;
srom_1(47497) <= 11937;
srom_1(47498) <= 62195;
srom_1(47499) <= 151498;
srom_1(47500) <= 279427;
srom_1(47501) <= 445384;
srom_1(47502) <= 648588;
srom_1(47503) <= 888089;
srom_1(47504) <= 1162762;
srom_1(47505) <= 1471319;
srom_1(47506) <= 1812314;
srom_1(47507) <= 2184148;
srom_1(47508) <= 2585076;
srom_1(47509) <= 3013219;
srom_1(47510) <= 3466569;
srom_1(47511) <= 3943000;
srom_1(47512) <= 4440279;
srom_1(47513) <= 4956072;
srom_1(47514) <= 5487961;
srom_1(47515) <= 6033453;
srom_1(47516) <= 6589989;
srom_1(47517) <= 7154959;
srom_1(47518) <= 7725714;
srom_1(47519) <= 8299578;
srom_1(47520) <= 8873859;
srom_1(47521) <= 9445865;
srom_1(47522) <= 10012913;
srom_1(47523) <= 10572344;
srom_1(47524) <= 11121534;
srom_1(47525) <= 11657909;
srom_1(47526) <= 12178953;
srom_1(47527) <= 12682223;
srom_1(47528) <= 13165359;
srom_1(47529) <= 13626094;
srom_1(47530) <= 14062270;
srom_1(47531) <= 14471839;
srom_1(47532) <= 14852883;
srom_1(47533) <= 15203613;
srom_1(47534) <= 15522385;
srom_1(47535) <= 15807704;
srom_1(47536) <= 16058233;
srom_1(47537) <= 16272796;
srom_1(47538) <= 16450388;
srom_1(47539) <= 16590175;
srom_1(47540) <= 16691502;
srom_1(47541) <= 16753894;
srom_1(47542) <= 16777058;
srom_1(47543) <= 16760886;
srom_1(47544) <= 16705453;
srom_1(47545) <= 16611020;
srom_1(47546) <= 16478029;
srom_1(47547) <= 16307104;
srom_1(47548) <= 16099047;
srom_1(47549) <= 15854833;
srom_1(47550) <= 15575606;
srom_1(47551) <= 15262678;
srom_1(47552) <= 14917515;
srom_1(47553) <= 14541735;
srom_1(47554) <= 14137101;
srom_1(47555) <= 13705511;
srom_1(47556) <= 13248988;
srom_1(47557) <= 12769673;
srom_1(47558) <= 12269813;
srom_1(47559) <= 11751753;
srom_1(47560) <= 11217923;
srom_1(47561) <= 10670824;
srom_1(47562) <= 10113024;
srom_1(47563) <= 9547137;
srom_1(47564) <= 8975817;
srom_1(47565) <= 8401744;
srom_1(47566) <= 7827609;
srom_1(47567) <= 7256105;
srom_1(47568) <= 6689911;
srom_1(47569) <= 6131684;
srom_1(47570) <= 5584040;
srom_1(47571) <= 5049547;
srom_1(47572) <= 4530712;
srom_1(47573) <= 4029969;
srom_1(47574) <= 3549664;
srom_1(47575) <= 3092051;
srom_1(47576) <= 2659275;
srom_1(47577) <= 2253367;
srom_1(47578) <= 1876228;
srom_1(47579) <= 1529628;
srom_1(47580) <= 1215192;
srom_1(47581) <= 934395;
srom_1(47582) <= 688553;
srom_1(47583) <= 478820;
srom_1(47584) <= 306178;
srom_1(47585) <= 171437;
srom_1(47586) <= 75230;
srom_1(47587) <= 18007;
srom_1(47588) <= 36;
srom_1(47589) <= 21403;
srom_1(47590) <= 82006;
srom_1(47591) <= 181561;
srom_1(47592) <= 319602;
srom_1(47593) <= 495482;
srom_1(47594) <= 708375;
srom_1(47595) <= 957283;
srom_1(47596) <= 1241040;
srom_1(47597) <= 1558313;
srom_1(47598) <= 1907617;
srom_1(47599) <= 2287312;
srom_1(47600) <= 2695618;
srom_1(47601) <= 3130620;
srom_1(47602) <= 3590279;
srom_1(47603) <= 4072439;
srom_1(47604) <= 4574839;
srom_1(47605) <= 5095123;
srom_1(47606) <= 5630851;
srom_1(47607) <= 6179511;
srom_1(47608) <= 6738531;
srom_1(47609) <= 7305288;
srom_1(47610) <= 7877125;
srom_1(47611) <= 8451361;
srom_1(47612) <= 9025303;
srom_1(47613) <= 9596259;
srom_1(47614) <= 10161551;
srom_1(47615) <= 10718530;
srom_1(47616) <= 11264583;
srom_1(47617) <= 11797150;
srom_1(47618) <= 12313733;
srom_1(47619) <= 12811909;
srom_1(47620) <= 13289343;
srom_1(47621) <= 13743796;
srom_1(47622) <= 14173137;
srom_1(47623) <= 14575351;
srom_1(47624) <= 14948555;
srom_1(47625) <= 15290996;
srom_1(47626) <= 15601069;
srom_1(47627) <= 15877321;
srom_1(47628) <= 16118456;
srom_1(47629) <= 16323343;
srom_1(47630) <= 16491021;
srom_1(47631) <= 16620704;
srom_1(47632) <= 16711784;
srom_1(47633) <= 16763834;
srom_1(47634) <= 16776609;
srom_1(47635) <= 16750050;
srom_1(47636) <= 16684282;
srom_1(47637) <= 16579612;
srom_1(47638) <= 16436532;
srom_1(47639) <= 16255712;
srom_1(47640) <= 16038001;
srom_1(47641) <= 15784419;
srom_1(47642) <= 15496155;
srom_1(47643) <= 15174562;
srom_1(47644) <= 14821147;
srom_1(47645) <= 14437568;
srom_1(47646) <= 14025623;
srom_1(47647) <= 13587245;
srom_1(47648) <= 13124488;
srom_1(47649) <= 12639522;
srom_1(47650) <= 12134623;
srom_1(47651) <= 11612158;
srom_1(47652) <= 11074576;
srom_1(47653) <= 10524399;
srom_1(47654) <= 9964206;
srom_1(47655) <= 9396625;
srom_1(47656) <= 8824316;
srom_1(47657) <= 8249965;
srom_1(47658) <= 7676264;
srom_1(47659) <= 7105903;
srom_1(47660) <= 6541557;
srom_1(47661) <= 5985872;
srom_1(47662) <= 5441455;
srom_1(47663) <= 4910858;
srom_1(47664) <= 4396570;
srom_1(47665) <= 3901001;
srom_1(47666) <= 3426477;
srom_1(47667) <= 2975221;
srom_1(47668) <= 2549351;
srom_1(47669) <= 2150863;
srom_1(47670) <= 1781626;
srom_1(47671) <= 1443371;
srom_1(47672) <= 1137685;
srom_1(47673) <= 866001;
srom_1(47674) <= 629593;
srom_1(47675) <= 429570;
srom_1(47676) <= 266869;
srom_1(47677) <= 142254;
srom_1(47678) <= 56309;
srom_1(47679) <= 9437;
srom_1(47680) <= 1858;
srom_1(47681) <= 33607;
srom_1(47682) <= 104536;
srom_1(47683) <= 214311;
srom_1(47684) <= 362419;
srom_1(47685) <= 548164;
srom_1(47686) <= 770676;
srom_1(47687) <= 1028910;
srom_1(47688) <= 1321657;
srom_1(47689) <= 1647544;
srom_1(47690) <= 2005041;
srom_1(47691) <= 2392473;
srom_1(47692) <= 2808023;
srom_1(47693) <= 3249742;
srom_1(47694) <= 3715560;
srom_1(47695) <= 4203290;
srom_1(47696) <= 4710647;
srom_1(47697) <= 5235252;
srom_1(47698) <= 5774643;
srom_1(47699) <= 6326293;
srom_1(47700) <= 6887613;
srom_1(47701) <= 7455972;
srom_1(47702) <= 8028704;
srom_1(47703) <= 8603124;
srom_1(47704) <= 9176538;
srom_1(47705) <= 9746257;
srom_1(47706) <= 10309610;
srom_1(47707) <= 10863954;
srom_1(47708) <= 11406691;
srom_1(47709) <= 11935275;
srom_1(47710) <= 12447227;
srom_1(47711) <= 12940147;
srom_1(47712) <= 13411723;
srom_1(47713) <= 13859744;
srom_1(47714) <= 14282110;
srom_1(47715) <= 14676838;
srom_1(47716) <= 15042079;
srom_1(47717) <= 15376119;
srom_1(47718) <= 15677393;
srom_1(47719) <= 15944487;
srom_1(47720) <= 16176148;
srom_1(47721) <= 16371292;
srom_1(47722) <= 16529002;
srom_1(47723) <= 16648538;
srom_1(47724) <= 16729341;
srom_1(47725) <= 16771032;
srom_1(47726) <= 16773414;
srom_1(47727) <= 16736477;
srom_1(47728) <= 16660394;
srom_1(47729) <= 16545522;
srom_1(47730) <= 16392399;
srom_1(47731) <= 16201744;
srom_1(47732) <= 15974450;
srom_1(47733) <= 15711584;
srom_1(47734) <= 15414378;
srom_1(47735) <= 15084225;
srom_1(47736) <= 14722674;
srom_1(47737) <= 14331421;
srom_1(47738) <= 13912300;
srom_1(47739) <= 13467276;
srom_1(47740) <= 12998437;
srom_1(47741) <= 12507980;
srom_1(47742) <= 11998207;
srom_1(47743) <= 11471507;
srom_1(47744) <= 10930350;
srom_1(47745) <= 10377274;
srom_1(47746) <= 9814872;
srom_1(47747) <= 9245782;
srom_1(47748) <= 8672673;
srom_1(47749) <= 8098231;
srom_1(47750) <= 7525151;
srom_1(47751) <= 6956120;
srom_1(47752) <= 6393807;
srom_1(47753) <= 5840848;
srom_1(47754) <= 5299836;
srom_1(47755) <= 4773309;
srom_1(47756) <= 4263734;
srom_1(47757) <= 3773503;
srom_1(47758) <= 3304914;
srom_1(47759) <= 2860164;
srom_1(47760) <= 2441338;
srom_1(47761) <= 2050402;
srom_1(47762) <= 1689187;
srom_1(47763) <= 1359388;
srom_1(47764) <= 1062552;
srom_1(47765) <= 800070;
srom_1(47766) <= 573173;
srom_1(47767) <= 382926;
srom_1(47768) <= 230220;
srom_1(47769) <= 115771;
srom_1(47770) <= 40117;
srom_1(47771) <= 3611;
srom_1(47772) <= 6426;
srom_1(47773) <= 48548;
srom_1(47774) <= 129779;
srom_1(47775) <= 249738;
srom_1(47776) <= 407863;
srom_1(47777) <= 603413;
srom_1(47778) <= 835471;
srom_1(47779) <= 1102947;
srom_1(47780) <= 1404589;
srom_1(47781) <= 1738981;
srom_1(47782) <= 2104555;
srom_1(47783) <= 2499597;
srom_1(47784) <= 2922256;
srom_1(47785) <= 3370547;
srom_1(47786) <= 3842370;
srom_1(47787) <= 4335512;
srom_1(47788) <= 4847660;
srom_1(47789) <= 5376413;
srom_1(47790) <= 5919291;
srom_1(47791) <= 6473749;
srom_1(47792) <= 7037186;
srom_1(47793) <= 7606960;
srom_1(47794) <= 8180400;
srom_1(47795) <= 8754816;
srom_1(47796) <= 9327515;
srom_1(47797) <= 9895811;
srom_1(47798) <= 10457039;
srom_1(47799) <= 11008568;
srom_1(47800) <= 11547810;
srom_1(47801) <= 12072238;
srom_1(47802) <= 12579393;
srom_1(47803) <= 13066895;
srom_1(47804) <= 13532459;
srom_1(47805) <= 13973902;
srom_1(47806) <= 14389153;
srom_1(47807) <= 14776266;
srom_1(47808) <= 15133425;
srom_1(47809) <= 15458955;
srom_1(47810) <= 15751330;
srom_1(47811) <= 16009178;
srom_1(47812) <= 16231291;
srom_1(47813) <= 16416627;
srom_1(47814) <= 16564317;
srom_1(47815) <= 16673668;
srom_1(47816) <= 16744168;
srom_1(47817) <= 16775485;
srom_1(47818) <= 16767474;
srom_1(47819) <= 16720171;
srom_1(47820) <= 16633799;
srom_1(47821) <= 16508762;
srom_1(47822) <= 16345646;
srom_1(47823) <= 16145218;
srom_1(47824) <= 15908416;
srom_1(47825) <= 15636351;
srom_1(47826) <= 15330299;
srom_1(47827) <= 14991695;
srom_1(47828) <= 14622127;
srom_1(47829) <= 14223328;
srom_1(47830) <= 13797168;
srom_1(47831) <= 13345645;
srom_1(47832) <= 12870877;
srom_1(47833) <= 12375090;
srom_1(47834) <= 11860609;
srom_1(47835) <= 11329846;
srom_1(47836) <= 10785291;
srom_1(47837) <= 10229498;
srom_1(47838) <= 9665071;
srom_1(47839) <= 9094659;
srom_1(47840) <= 8520936;
srom_1(47841) <= 7946592;
srom_1(47842) <= 7374322;
srom_1(47843) <= 6806807;
srom_1(47844) <= 6246710;
srom_1(47845) <= 5696657;
srom_1(47846) <= 5159228;
srom_1(47847) <= 4636942;
srom_1(47848) <= 4132249;
srom_1(47849) <= 3647516;
srom_1(47850) <= 3185015;
srom_1(47851) <= 2746916;
srom_1(47852) <= 2335273;
srom_1(47853) <= 1952015;
srom_1(47854) <= 1598941;
srom_1(47855) <= 1277707;
srom_1(47856) <= 989817;
srom_1(47857) <= 736623;
srom_1(47858) <= 519312;
srom_1(47859) <= 338903;
srom_1(47860) <= 196241;
srom_1(47861) <= 91997;
srom_1(47862) <= 26658;
srom_1(47863) <= 531;
srom_1(47864) <= 13738;
srom_1(47865) <= 66218;
srom_1(47866) <= 157725;
srom_1(47867) <= 287829;
srom_1(47868) <= 455921;
srom_1(47869) <= 661211;
srom_1(47870) <= 902738;
srom_1(47871) <= 1179369;
srom_1(47872) <= 1489807;
srom_1(47873) <= 1832595;
srom_1(47874) <= 2206127;
srom_1(47875) <= 2608650;
srom_1(47876) <= 3038278;
srom_1(47877) <= 3492995;
srom_1(47878) <= 3970669;
srom_1(47879) <= 4469061;
srom_1(47880) <= 4985832;
srom_1(47881) <= 5518561;
srom_1(47882) <= 6064748;
srom_1(47883) <= 6621832;
srom_1(47884) <= 7187202;
srom_1(47885) <= 7758205;
srom_1(47886) <= 8332165;
srom_1(47887) <= 8906389;
srom_1(47888) <= 9478185;
srom_1(47889) <= 10044871;
srom_1(47890) <= 10603791;
srom_1(47891) <= 11152323;
srom_1(47892) <= 11687895;
srom_1(47893) <= 12207996;
srom_1(47894) <= 12710186;
srom_1(47895) <= 13192111;
srom_1(47896) <= 13651510;
srom_1(47897) <= 14086230;
srom_1(47898) <= 14494232;
srom_1(47899) <= 14873603;
srom_1(47900) <= 15222563;
srom_1(47901) <= 15539476;
srom_1(47902) <= 15822856;
srom_1(47903) <= 16071375;
srom_1(47904) <= 16283866;
srom_1(47905) <= 16459334;
srom_1(47906) <= 16596956;
srom_1(47907) <= 16696086;
srom_1(47908) <= 16756259;
srom_1(47909) <= 16777193;
srom_1(47910) <= 16758790;
srom_1(47911) <= 16701137;
srom_1(47912) <= 16604504;
srom_1(47913) <= 16469343;
srom_1(47914) <= 16296289;
srom_1(47915) <= 16086153;
srom_1(47916) <= 15839920;
srom_1(47917) <= 15558746;
srom_1(47918) <= 15243949;
srom_1(47919) <= 14897004;
srom_1(47920) <= 14519540;
srom_1(47921) <= 14113325;
srom_1(47922) <= 13680265;
srom_1(47923) <= 13222391;
srom_1(47924) <= 12741849;
srom_1(47925) <= 12240894;
srom_1(47926) <= 11721874;
srom_1(47927) <= 11187223;
srom_1(47928) <= 10639448;
srom_1(47929) <= 10081119;
srom_1(47930) <= 9514853;
srom_1(47931) <= 8943305;
srom_1(47932) <= 8369156;
srom_1(47933) <= 7795099;
srom_1(47934) <= 7223824;
srom_1(47935) <= 6658012;
srom_1(47936) <= 6100315;
srom_1(47937) <= 5553348;
srom_1(47938) <= 5019677;
srom_1(47939) <= 4501804;
srom_1(47940) <= 4002158;
srom_1(47941) <= 3523081;
srom_1(47942) <= 3066821;
srom_1(47943) <= 2635516;
srom_1(47944) <= 2231189;
srom_1(47945) <= 1855736;
srom_1(47946) <= 1510919;
srom_1(47947) <= 1198353;
srom_1(47948) <= 919505;
srom_1(47949) <= 675682;
srom_1(47950) <= 468027;
srom_1(47951) <= 297515;
srom_1(47952) <= 164945;
srom_1(47953) <= 70938;
srom_1(47954) <= 15936;
srom_1(47955) <= 196;
srom_1(47956) <= 23792;
srom_1(47957) <= 86614;
srom_1(47958) <= 188366;
srom_1(47959) <= 328573;
srom_1(47960) <= 506575;
srom_1(47961) <= 721539;
srom_1(47962) <= 972457;
srom_1(47963) <= 1258152;
srom_1(47964) <= 1577283;
srom_1(47965) <= 1928356;
srom_1(47966) <= 2309722;
srom_1(47967) <= 2719595;
srom_1(47968) <= 3156051;
srom_1(47969) <= 3617045;
srom_1(47970) <= 4100415;
srom_1(47971) <= 4603893;
srom_1(47972) <= 5125119;
srom_1(47973) <= 5661648;
srom_1(47974) <= 6210965;
srom_1(47975) <= 6770494;
srom_1(47976) <= 7337611;
srom_1(47977) <= 7909656;
srom_1(47978) <= 8483948;
srom_1(47979) <= 9057792;
srom_1(47980) <= 9628498;
srom_1(47981) <= 10193390;
srom_1(47982) <= 10749818;
srom_1(47983) <= 11295174;
srom_1(47984) <= 11826900;
srom_1(47985) <= 12342503;
srom_1(47986) <= 12839565;
srom_1(47987) <= 13315754;
srom_1(47988) <= 13768839;
srom_1(47989) <= 14196694;
srom_1(47990) <= 14597312;
srom_1(47991) <= 14968816;
srom_1(47992) <= 15309463;
srom_1(47993) <= 15617656;
srom_1(47994) <= 15891949;
srom_1(47995) <= 16131056;
srom_1(47996) <= 16333857;
srom_1(47997) <= 16499399;
srom_1(47998) <= 16626907;
srom_1(47999) <= 16715783;
srom_1(48000) <= 16765610;
srom_1(48001) <= 16776155;
srom_1(48002) <= 16747367;
srom_1(48003) <= 16679382;
srom_1(48004) <= 16572519;
srom_1(48005) <= 16427278;
srom_1(48006) <= 16244342;
srom_1(48007) <= 16024567;
srom_1(48008) <= 15768985;
srom_1(48009) <= 15478793;
srom_1(48010) <= 15155353;
srom_1(48011) <= 14800182;
srom_1(48012) <= 14414945;
srom_1(48013) <= 14001447;
srom_1(48014) <= 13561630;
srom_1(48015) <= 13097554;
srom_1(48016) <= 12611397;
srom_1(48017) <= 12105437;
srom_1(48018) <= 11582048;
srom_1(48019) <= 11043684;
srom_1(48020) <= 10492869;
srom_1(48021) <= 9932186;
srom_1(48022) <= 9364265;
srom_1(48023) <= 8791769;
srom_1(48024) <= 8217383;
srom_1(48025) <= 7643799;
srom_1(48026) <= 7073708;
srom_1(48027) <= 6509783;
srom_1(48028) <= 5954668;
srom_1(48029) <= 5410967;
srom_1(48030) <= 4881229;
srom_1(48031) <= 4367939;
srom_1(48032) <= 3873503;
srom_1(48033) <= 3400239;
srom_1(48034) <= 2950368;
srom_1(48035) <= 2525999;
srom_1(48036) <= 2129121;
srom_1(48037) <= 1761596;
srom_1(48038) <= 1425148;
srom_1(48039) <= 1121353;
srom_1(48040) <= 851638;
srom_1(48041) <= 617265;
srom_1(48042) <= 419335;
srom_1(48043) <= 258776;
srom_1(48044) <= 136341;
srom_1(48045) <= 52603;
srom_1(48046) <= 7955;
srom_1(48047) <= 2607;
srom_1(48048) <= 36585;
srom_1(48049) <= 109727;
srom_1(48050) <= 221692;
srom_1(48051) <= 371955;
srom_1(48052) <= 559810;
srom_1(48053) <= 784377;
srom_1(48054) <= 1044604;
srom_1(48055) <= 1339268;
srom_1(48056) <= 1666990;
srom_1(48057) <= 2026231;
srom_1(48058) <= 2415308;
srom_1(48059) <= 2832396;
srom_1(48060) <= 3275538;
srom_1(48061) <= 3742658;
srom_1(48062) <= 4231564;
srom_1(48063) <= 4739964;
srom_1(48064) <= 5265473;
srom_1(48065) <= 5805628;
srom_1(48066) <= 6357896;
srom_1(48067) <= 6919686;
srom_1(48068) <= 7488364;
srom_1(48069) <= 8061264;
srom_1(48070) <= 8635699;
srom_1(48071) <= 9208976;
srom_1(48072) <= 9778405;
srom_1(48073) <= 10341317;
srom_1(48074) <= 10895072;
srom_1(48075) <= 11437074;
srom_1(48076) <= 11964780;
srom_1(48077) <= 12475716;
srom_1(48078) <= 12967486;
srom_1(48079) <= 13437785;
srom_1(48080) <= 13884406;
srom_1(48081) <= 14305255;
srom_1(48082) <= 14698360;
srom_1(48083) <= 15061875;
srom_1(48084) <= 15394098;
srom_1(48085) <= 15693469;
srom_1(48086) <= 15958585;
srom_1(48087) <= 16188203;
srom_1(48088) <= 16381246;
srom_1(48089) <= 16536809;
srom_1(48090) <= 16654162;
srom_1(48091) <= 16732755;
srom_1(48092) <= 16772219;
srom_1(48093) <= 16772370;
srom_1(48094) <= 16733206;
srom_1(48095) <= 16654912;
srom_1(48096) <= 16537854;
srom_1(48097) <= 16382582;
srom_1(48098) <= 16189823;
srom_1(48099) <= 15960482;
srom_1(48100) <= 15695633;
srom_1(48101) <= 15396519;
srom_1(48102) <= 15064543;
srom_1(48103) <= 14701261;
srom_1(48104) <= 14308377;
srom_1(48105) <= 13887732;
srom_1(48106) <= 13441301;
srom_1(48107) <= 12971176;
srom_1(48108) <= 12479561;
srom_1(48109) <= 11968763;
srom_1(48110) <= 11441176;
srom_1(48111) <= 10899275;
srom_1(48112) <= 10345600;
srom_1(48113) <= 9782748;
srom_1(48114) <= 9213358;
srom_1(48115) <= 8640101;
srom_1(48116) <= 8065665;
srom_1(48117) <= 7492743;
srom_1(48118) <= 6924022;
srom_1(48119) <= 6362169;
srom_1(48120) <= 5809819;
srom_1(48121) <= 5269561;
srom_1(48122) <= 4743930;
srom_1(48123) <= 4235390;
srom_1(48124) <= 3746325;
srom_1(48125) <= 3279030;
srom_1(48126) <= 2835696;
srom_1(48127) <= 2418401;
srom_1(48128) <= 2029102;
srom_1(48129) <= 1669626;
srom_1(48130) <= 1341657;
srom_1(48131) <= 1046733;
srom_1(48132) <= 786238;
srom_1(48133) <= 561393;
srom_1(48134) <= 373253;
srom_1(48135) <= 222699;
srom_1(48136) <= 110438;
srom_1(48137) <= 36997;
srom_1(48138) <= 2718;
srom_1(48139) <= 7765;
srom_1(48140) <= 52111;
srom_1(48141) <= 135551;
srom_1(48142) <= 257692;
srom_1(48143) <= 417961;
srom_1(48144) <= 615608;
srom_1(48145) <= 849705;
srom_1(48146) <= 1119155;
srom_1(48147) <= 1422693;
srom_1(48148) <= 1758897;
srom_1(48149) <= 2126190;
srom_1(48150) <= 2522849;
srom_1(48151) <= 2947015;
srom_1(48152) <= 3396699;
srom_1(48153) <= 3869791;
srom_1(48154) <= 4364074;
srom_1(48155) <= 4877229;
srom_1(48156) <= 5406850;
srom_1(48157) <= 5950454;
srom_1(48158) <= 6505491;
srom_1(48159) <= 7069358;
srom_1(48160) <= 7639412;
srom_1(48161) <= 8212979;
srom_1(48162) <= 8787370;
srom_1(48163) <= 9359891;
srom_1(48164) <= 9927857;
srom_1(48165) <= 10488605;
srom_1(48166) <= 11039505;
srom_1(48167) <= 11577975;
srom_1(48168) <= 12101488;
srom_1(48169) <= 12607591;
srom_1(48170) <= 13093909;
srom_1(48171) <= 13558162;
srom_1(48172) <= 13998174;
srom_1(48173) <= 14411880;
srom_1(48174) <= 14797341;
srom_1(48175) <= 15152750;
srom_1(48176) <= 15476439;
srom_1(48177) <= 15766890;
srom_1(48178) <= 16022743;
srom_1(48179) <= 16242796;
srom_1(48180) <= 16426018;
srom_1(48181) <= 16571551;
srom_1(48182) <= 16678710;
srom_1(48183) <= 16746994;
srom_1(48184) <= 16776083;
srom_1(48185) <= 16765841;
srom_1(48186) <= 16716314;
srom_1(48187) <= 16627736;
srom_1(48188) <= 16500522;
srom_1(48189) <= 16335269;
srom_1(48190) <= 16132750;
srom_1(48191) <= 15893917;
srom_1(48192) <= 15619889;
srom_1(48193) <= 15311951;
srom_1(48194) <= 14971547;
srom_1(48195) <= 14600273;
srom_1(48196) <= 14199871;
srom_1(48197) <= 13772217;
srom_1(48198) <= 13319318;
srom_1(48199) <= 12843297;
srom_1(48200) <= 12346387;
srom_1(48201) <= 11830917;
srom_1(48202) <= 11299305;
srom_1(48203) <= 10754044;
srom_1(48204) <= 10197690;
srom_1(48205) <= 9632853;
srom_1(48206) <= 9062182;
srom_1(48207) <= 8488351;
srom_1(48208) <= 7914053;
srom_1(48209) <= 7341981;
srom_1(48210) <= 6774816;
srom_1(48211) <= 6215219;
srom_1(48212) <= 5665813;
srom_1(48213) <= 5129176;
srom_1(48214) <= 4607824;
srom_1(48215) <= 4104200;
srom_1(48216) <= 3620668;
srom_1(48217) <= 3159494;
srom_1(48218) <= 2722842;
srom_1(48219) <= 2312758;
srom_1(48220) <= 1931166;
srom_1(48221) <= 1579855;
srom_1(48222) <= 1260472;
srom_1(48223) <= 974516;
srom_1(48224) <= 723327;
srom_1(48225) <= 508084;
srom_1(48226) <= 329794;
srom_1(48227) <= 189296;
srom_1(48228) <= 87246;
srom_1(48229) <= 24125;
srom_1(48230) <= 227;
srom_1(48231) <= 15666;
srom_1(48232) <= 70368;
srom_1(48233) <= 164077;
srom_1(48234) <= 296354;
srom_1(48235) <= 466578;
srom_1(48236) <= 673951;
srom_1(48237) <= 917501;
srom_1(48238) <= 1196085;
srom_1(48239) <= 1508398;
srom_1(48240) <= 1852975;
srom_1(48241) <= 2228199;
srom_1(48242) <= 2632311;
srom_1(48243) <= 3063417;
srom_1(48244) <= 3519494;
srom_1(48245) <= 3998405;
srom_1(48246) <= 4497902;
srom_1(48247) <= 5015644;
srom_1(48248) <= 5549204;
srom_1(48249) <= 6096078;
srom_1(48250) <= 6653703;
srom_1(48251) <= 7219463;
srom_1(48252) <= 7790705;
srom_1(48253) <= 8364752;
srom_1(48254) <= 8938910;
srom_1(48255) <= 9510488;
srom_1(48256) <= 10076805;
srom_1(48257) <= 10635206;
srom_1(48258) <= 11183071;
srom_1(48259) <= 11717832;
srom_1(48260) <= 12236981;
srom_1(48261) <= 12738084;
srom_1(48262) <= 13218791;
srom_1(48263) <= 13676847;
srom_1(48264) <= 14110105;
srom_1(48265) <= 14516533;
srom_1(48266) <= 14894225;
srom_1(48267) <= 15241409;
srom_1(48268) <= 15556459;
srom_1(48269) <= 15837896;
srom_1(48270) <= 16084401;
srom_1(48271) <= 16294818;
srom_1(48272) <= 16468159;
srom_1(48273) <= 16603613;
srom_1(48274) <= 16700544;
srom_1(48275) <= 16758498;
srom_1(48276) <= 16777202;
srom_1(48277) <= 16756569;
srom_1(48278) <= 16696696;
srom_1(48279) <= 16597863;
srom_1(48280) <= 16460534;
srom_1(48281) <= 16285353;
srom_1(48282) <= 16073142;
srom_1(48283) <= 15824895;
srom_1(48284) <= 15541777;
srom_1(48285) <= 15225116;
srom_1(48286) <= 14876395;
srom_1(48287) <= 14497251;
srom_1(48288) <= 14089462;
srom_1(48289) <= 13654939;
srom_1(48290) <= 13195721;
srom_1(48291) <= 12713960;
srom_1(48292) <= 12211917;
srom_1(48293) <= 11691944;
srom_1(48294) <= 11156481;
srom_1(48295) <= 10608039;
srom_1(48296) <= 10049189;
srom_1(48297) <= 9482551;
srom_1(48298) <= 8910784;
srom_1(48299) <= 8336569;
srom_1(48300) <= 7762597;
srom_1(48301) <= 7191561;
srom_1(48302) <= 6626138;
srom_1(48303) <= 6068980;
srom_1(48304) <= 5522700;
srom_1(48305) <= 4989858;
srom_1(48306) <= 4472955;
srom_1(48307) <= 3974414;
srom_1(48308) <= 3496572;
srom_1(48309) <= 3041670;
srom_1(48310) <= 2611843;
srom_1(48311) <= 2209104;
srom_1(48312) <= 1835343;
srom_1(48313) <= 1492313;
srom_1(48314) <= 1181622;
srom_1(48315) <= 904727;
srom_1(48316) <= 662926;
srom_1(48317) <= 457354;
srom_1(48318) <= 288974;
srom_1(48319) <= 158576;
srom_1(48320) <= 66772;
srom_1(48321) <= 13991;
srom_1(48322) <= 482;
srom_1(48323) <= 26308;
srom_1(48324) <= 91347;
srom_1(48325) <= 195295;
srom_1(48326) <= 337665;
srom_1(48327) <= 517788;
srom_1(48328) <= 734820;
srom_1(48329) <= 987743;
srom_1(48330) <= 1275371;
srom_1(48331) <= 1596356;
srom_1(48332) <= 1949192;
srom_1(48333) <= 2332225;
srom_1(48334) <= 2743658;
srom_1(48335) <= 3181562;
srom_1(48336) <= 3643884;
srom_1(48337) <= 4128455;
srom_1(48338) <= 4633004;
srom_1(48339) <= 5155164;
srom_1(48340) <= 5692487;
srom_1(48341) <= 6242452;
srom_1(48342) <= 6802482;
srom_1(48343) <= 7369950;
srom_1(48344) <= 7942195;
srom_1(48345) <= 8516532;
srom_1(48346) <= 9090271;
srom_1(48347) <= 9660718;
srom_1(48348) <= 10225201;
srom_1(48349) <= 10781071;
srom_1(48350) <= 11325721;
srom_1(48351) <= 11856599;
srom_1(48352) <= 12371214;
srom_1(48353) <= 12867153;
srom_1(48354) <= 13342091;
srom_1(48355) <= 13793801;
srom_1(48356) <= 14220163;
srom_1(48357) <= 14619179;
srom_1(48358) <= 14988978;
srom_1(48359) <= 15327826;
srom_1(48360) <= 15634133;
srom_1(48361) <= 15906463;
srom_1(48362) <= 16143540;
srom_1(48363) <= 16344251;
srom_1(48364) <= 16507655;
srom_1(48365) <= 16632987;
srom_1(48366) <= 16719657;
srom_1(48367) <= 16767261;
srom_1(48368) <= 16775574;
srom_1(48369) <= 16744557;
srom_1(48370) <= 16674357;
srom_1(48371) <= 16565302;
srom_1(48372) <= 16417904;
srom_1(48373) <= 16232853;
srom_1(48374) <= 16011018;
srom_1(48375) <= 15753439;
srom_1(48376) <= 15461324;
srom_1(48377) <= 15136042;
srom_1(48378) <= 14779120;
srom_1(48379) <= 14392230;
srom_1(48380) <= 13977187;
srom_1(48381) <= 13535937;
srom_1(48382) <= 13070550;
srom_1(48383) <= 12583207;
srom_1(48384) <= 12076195;
srom_1(48385) <= 11551890;
srom_1(48386) <= 11012751;
srom_1(48387) <= 10461307;
srom_1(48388) <= 9900143;
srom_1(48389) <= 9331891;
srom_1(48390) <= 8759216;
srom_1(48391) <= 8184803;
srom_1(48392) <= 7611345;
srom_1(48393) <= 7041533;
srom_1(48394) <= 6478037;
srom_1(48395) <= 5923501;
srom_1(48396) <= 5380524;
srom_1(48397) <= 4851653;
srom_1(48398) <= 4339369;
srom_1(48399) <= 3846072;
srom_1(48400) <= 3374077;
srom_1(48401) <= 2925597;
srom_1(48402) <= 2502735;
srom_1(48403) <= 2107473;
srom_1(48404) <= 1741666;
srom_1(48405) <= 1407029;
srom_1(48406) <= 1105131;
srom_1(48407) <= 837388;
srom_1(48408) <= 605055;
srom_1(48409) <= 409221;
srom_1(48410) <= 250806;
srom_1(48411) <= 130551;
srom_1(48412) <= 49022;
srom_1(48413) <= 6600;
srom_1(48414) <= 3483;
srom_1(48415) <= 39688;
srom_1(48416) <= 115043;
srom_1(48417) <= 229196;
srom_1(48418) <= 381612;
srom_1(48419) <= 571574;
srom_1(48420) <= 798194;
srom_1(48421) <= 1060408;
srom_1(48422) <= 1356986;
srom_1(48423) <= 1686537;
srom_1(48424) <= 2047517;
srom_1(48425) <= 2438233;
srom_1(48426) <= 2856852;
srom_1(48427) <= 3301411;
srom_1(48428) <= 3769826;
srom_1(48429) <= 4259900;
srom_1(48430) <= 4769335;
srom_1(48431) <= 5295742;
srom_1(48432) <= 5836652;
srom_1(48433) <= 6389529;
srom_1(48434) <= 6951781;
srom_1(48435) <= 7520771;
srom_1(48436) <= 8093830;
srom_1(48437) <= 8668271;
srom_1(48438) <= 9241401;
srom_1(48439) <= 9810532;
srom_1(48440) <= 10372995;
srom_1(48441) <= 10926152;
srom_1(48442) <= 11467410;
srom_1(48443) <= 11994231;
srom_1(48444) <= 12504143;
srom_1(48445) <= 12994757;
srom_1(48446) <= 13463770;
srom_1(48447) <= 13908984;
srom_1(48448) <= 14328312;
srom_1(48449) <= 14719786;
srom_1(48450) <= 15081571;
srom_1(48451) <= 15411970;
srom_1(48452) <= 15709435;
srom_1(48453) <= 15972569;
srom_1(48454) <= 16200140;
srom_1(48455) <= 16391080;
srom_1(48456) <= 16544493;
srom_1(48457) <= 16659661;
srom_1(48458) <= 16736042;
srom_1(48459) <= 16773280;
srom_1(48460) <= 16771200;
srom_1(48461) <= 16729810;
srom_1(48462) <= 16649306;
srom_1(48463) <= 16530064;
srom_1(48464) <= 16372644;
srom_1(48465) <= 16177784;
srom_1(48466) <= 15946399;
srom_1(48467) <= 15679572;
srom_1(48468) <= 15378555;
srom_1(48469) <= 15044760;
srom_1(48470) <= 14679752;
srom_1(48471) <= 14285243;
srom_1(48472) <= 13863082;
srom_1(48473) <= 13415250;
srom_1(48474) <= 12943846;
srom_1(48475) <= 12451081;
srom_1(48476) <= 11939265;
srom_1(48477) <= 11410800;
srom_1(48478) <= 10868162;
srom_1(48479) <= 10313897;
srom_1(48480) <= 9750603;
srom_1(48481) <= 9180922;
srom_1(48482) <= 8607526;
srom_1(48483) <= 8033104;
srom_1(48484) <= 7460348;
srom_1(48485) <= 6891946;
srom_1(48486) <= 6330562;
srom_1(48487) <= 5778828;
srom_1(48488) <= 5239333;
srom_1(48489) <= 4714606;
srom_1(48490) <= 4207108;
srom_1(48491) <= 3719218;
srom_1(48492) <= 3253224;
srom_1(48493) <= 2811312;
srom_1(48494) <= 2395554;
srom_1(48495) <= 2007899;
srom_1(48496) <= 1650166;
srom_1(48497) <= 1324031;
srom_1(48498) <= 1031025;
srom_1(48499) <= 772521;
srom_1(48500) <= 549731;
srom_1(48501) <= 363701;
srom_1(48502) <= 215302;
srom_1(48503) <= 105230;
srom_1(48504) <= 34002;
srom_1(48505) <= 1952;
srom_1(48506) <= 9230;
srom_1(48507) <= 55801;
srom_1(48508) <= 141448;
srom_1(48509) <= 265768;
srom_1(48510) <= 428180;
srom_1(48511) <= 627920;
srom_1(48512) <= 864053;
srom_1(48513) <= 1135472;
srom_1(48514) <= 1440902;
srom_1(48515) <= 1778913;
srom_1(48516) <= 2147919;
srom_1(48517) <= 2546190;
srom_1(48518) <= 2971858;
srom_1(48519) <= 3422926;
srom_1(48520) <= 3897281;
srom_1(48521) <= 4392697;
srom_1(48522) <= 4906851;
srom_1(48523) <= 5437332;
srom_1(48524) <= 5981653;
srom_1(48525) <= 6537261;
srom_1(48526) <= 7101551;
srom_1(48527) <= 7671875;
srom_1(48528) <= 8245561;
srom_1(48529) <= 8819918;
srom_1(48530) <= 9392252;
srom_1(48531) <= 9959880;
srom_1(48532) <= 10520139;
srom_1(48533) <= 11070403;
srom_1(48534) <= 11608091;
srom_1(48535) <= 12130682;
srom_1(48536) <= 12635725;
srom_1(48537) <= 13120852;
srom_1(48538) <= 13583787;
srom_1(48539) <= 14022361;
srom_1(48540) <= 14434516;
srom_1(48541) <= 14818320;
srom_1(48542) <= 15171972;
srom_1(48543) <= 15493815;
srom_1(48544) <= 15782339;
srom_1(48545) <= 16036192;
srom_1(48546) <= 16254182;
srom_1(48547) <= 16435288;
srom_1(48548) <= 16578661;
srom_1(48549) <= 16683627;
srom_1(48550) <= 16749695;
srom_1(48551) <= 16776555;
srom_1(48552) <= 16764081;
srom_1(48553) <= 16712332;
srom_1(48554) <= 16621550;
srom_1(48555) <= 16492160;
srom_1(48556) <= 16324771;
srom_1(48557) <= 16120166;
srom_1(48558) <= 15879305;
srom_1(48559) <= 15603317;
srom_1(48560) <= 15293498;
srom_1(48561) <= 14951299;
srom_1(48562) <= 14578325;
srom_1(48563) <= 14176325;
srom_1(48564) <= 13747185;
srom_1(48565) <= 13292917;
srom_1(48566) <= 12815651;
srom_1(48567) <= 12317624;
srom_1(48568) <= 11801174;
srom_1(48569) <= 11268720;
srom_1(48570) <= 10722761;
srom_1(48571) <= 10165856;
srom_1(48572) <= 9600617;
srom_1(48573) <= 9029694;
srom_1(48574) <= 8455765;
srom_1(48575) <= 7881521;
srom_1(48576) <= 7309655;
srom_1(48577) <= 6742849;
srom_1(48578) <= 6183760;
srom_1(48579) <= 5635011;
srom_1(48580) <= 5099174;
srom_1(48581) <= 4578762;
srom_1(48582) <= 4076216;
srom_1(48583) <= 3593892;
srom_1(48584) <= 3134052;
srom_1(48585) <= 2698853;
srom_1(48586) <= 2290335;
srom_1(48587) <= 1910414;
srom_1(48588) <= 1560871;
srom_1(48589) <= 1243346;
srom_1(48590) <= 959327;
srom_1(48591) <= 710147;
srom_1(48592) <= 496974;
srom_1(48593) <= 320807;
srom_1(48594) <= 182474;
srom_1(48595) <= 82621;
srom_1(48596) <= 21718;
srom_1(48597) <= 50;
srom_1(48598) <= 17719;
srom_1(48599) <= 74643;
srom_1(48600) <= 170553;
srom_1(48601) <= 305000;
srom_1(48602) <= 477354;
srom_1(48603) <= 686807;
srom_1(48604) <= 932376;
srom_1(48605) <= 1212910;
srom_1(48606) <= 1527093;
srom_1(48607) <= 1873453;
srom_1(48608) <= 2250364;
srom_1(48609) <= 2656059;
srom_1(48610) <= 3088637;
srom_1(48611) <= 3546067;
srom_1(48612) <= 4026206;
srom_1(48613) <= 4526802;
srom_1(48614) <= 5045507;
srom_1(48615) <= 5579889;
srom_1(48616) <= 6127442;
srom_1(48617) <= 6685599;
srom_1(48618) <= 7251741;
srom_1(48619) <= 7823215;
srom_1(48620) <= 8397340;
srom_1(48621) <= 8971424;
srom_1(48622) <= 9542775;
srom_1(48623) <= 10108713;
srom_1(48624) <= 10666586;
srom_1(48625) <= 11213776;
srom_1(48626) <= 11747718;
srom_1(48627) <= 12265908;
srom_1(48628) <= 12765916;
srom_1(48629) <= 13245398;
srom_1(48630) <= 13702104;
srom_1(48631) <= 14133893;
srom_1(48632) <= 14538741;
srom_1(48633) <= 14914749;
srom_1(48634) <= 15260153;
srom_1(48635) <= 15573334;
srom_1(48636) <= 15852824;
srom_1(48637) <= 16097311;
srom_1(48638) <= 16305650;
srom_1(48639) <= 16476862;
srom_1(48640) <= 16610147;
srom_1(48641) <= 16704877;
srom_1(48642) <= 16760610;
srom_1(48643) <= 16777084;
srom_1(48644) <= 16754221;
srom_1(48645) <= 16692129;
srom_1(48646) <= 16591098;
srom_1(48647) <= 16451604;
srom_1(48648) <= 16274299;
srom_1(48649) <= 16060016;
srom_1(48650) <= 15809759;
srom_1(48651) <= 15524701;
srom_1(48652) <= 15206180;
srom_1(48653) <= 14855689;
srom_1(48654) <= 14474871;
srom_1(48655) <= 14065513;
srom_1(48656) <= 13629534;
srom_1(48657) <= 13168978;
srom_1(48658) <= 12686006;
srom_1(48659) <= 12182882;
srom_1(48660) <= 11661965;
srom_1(48661) <= 11125698;
srom_1(48662) <= 10576596;
srom_1(48663) <= 10017233;
srom_1(48664) <= 9450234;
srom_1(48665) <= 8878256;
srom_1(48666) <= 8303982;
srom_1(48667) <= 7730105;
srom_1(48668) <= 7159316;
srom_1(48669) <= 6594291;
srom_1(48670) <= 6037680;
srom_1(48671) <= 5492094;
srom_1(48672) <= 4960091;
srom_1(48673) <= 4444165;
srom_1(48674) <= 3946736;
srom_1(48675) <= 3470136;
srom_1(48676) <= 3016601;
srom_1(48677) <= 2588257;
srom_1(48678) <= 2187113;
srom_1(48679) <= 1815049;
srom_1(48680) <= 1473812;
srom_1(48681) <= 1165000;
srom_1(48682) <= 890062;
srom_1(48683) <= 650288;
srom_1(48684) <= 446801;
srom_1(48685) <= 280556;
srom_1(48686) <= 152332;
srom_1(48687) <= 62731;
srom_1(48688) <= 12173;
srom_1(48689) <= 895;
srom_1(48690) <= 28950;
srom_1(48691) <= 96206;
srom_1(48692) <= 202348;
srom_1(48693) <= 346878;
srom_1(48694) <= 529119;
srom_1(48695) <= 748215;
srom_1(48696) <= 1003140;
srom_1(48697) <= 1292698;
srom_1(48698) <= 1615531;
srom_1(48699) <= 1970125;
srom_1(48700) <= 2354818;
srom_1(48701) <= 2767806;
srom_1(48702) <= 3207151;
srom_1(48703) <= 3670793;
srom_1(48704) <= 4156560;
srom_1(48705) <= 4662171;
srom_1(48706) <= 5185258;
srom_1(48707) <= 5723366;
srom_1(48708) <= 6273972;
srom_1(48709) <= 6834494;
srom_1(48710) <= 7402304;
srom_1(48711) <= 7974739;
srom_1(48712) <= 8549115;
srom_1(48713) <= 9122739;
srom_1(48714) <= 9692920;
srom_1(48715) <= 10256984;
srom_1(48716) <= 10812287;
srom_1(48717) <= 11356224;
srom_1(48718) <= 11886245;
srom_1(48719) <= 12399865;
srom_1(48720) <= 12894674;
srom_1(48721) <= 13368353;
srom_1(48722) <= 13818681;
srom_1(48723) <= 14243544;
srom_1(48724) <= 14640952;
srom_1(48725) <= 15009041;
srom_1(48726) <= 15346084;
srom_1(48727) <= 15650501;
srom_1(48728) <= 15920864;
srom_1(48729) <= 16155906;
srom_1(48730) <= 16354525;
srom_1(48731) <= 16515789;
srom_1(48732) <= 16638941;
srom_1(48733) <= 16723405;
srom_1(48734) <= 16768784;
srom_1(48735) <= 16774866;
srom_1(48736) <= 16741621;
srom_1(48737) <= 16669207;
srom_1(48738) <= 16557962;
srom_1(48739) <= 16408408;
srom_1(48740) <= 16221246;
srom_1(48741) <= 15997354;
srom_1(48742) <= 15737783;
srom_1(48743) <= 15443748;
srom_1(48744) <= 15116630;
srom_1(48745) <= 14757961;
srom_1(48746) <= 14369425;
srom_1(48747) <= 13952842;
srom_1(48748) <= 13510167;
srom_1(48749) <= 13043475;
srom_1(48750) <= 12554954;
srom_1(48751) <= 12046897;
srom_1(48752) <= 11521684;
srom_1(48753) <= 10981779;
srom_1(48754) <= 10429714;
srom_1(48755) <= 9868077;
srom_1(48756) <= 9299503;
srom_1(48757) <= 8726657;
srom_1(48758) <= 8152226;
srom_1(48759) <= 7578904;
srom_1(48760) <= 7009378;
srom_1(48761) <= 6446320;
srom_1(48762) <= 5892370;
srom_1(48763) <= 5350126;
srom_1(48764) <= 4822131;
srom_1(48765) <= 4310859;
srom_1(48766) <= 3818710;
srom_1(48767) <= 3347991;
srom_1(48768) <= 2900908;
srom_1(48769) <= 2479560;
srom_1(48770) <= 2085921;
srom_1(48771) <= 1721837;
srom_1(48772) <= 1389016;
srom_1(48773) <= 1089019;
srom_1(48774) <= 823252;
srom_1(48775) <= 592961;
srom_1(48776) <= 399227;
srom_1(48777) <= 242958;
srom_1(48778) <= 124887;
srom_1(48779) <= 45567;
srom_1(48780) <= 5370;
srom_1(48781) <= 4486;
srom_1(48782) <= 42917;
srom_1(48783) <= 120484;
srom_1(48784) <= 236823;
srom_1(48785) <= 391389;
srom_1(48786) <= 583457;
srom_1(48787) <= 812125;
srom_1(48788) <= 1076322;
srom_1(48789) <= 1374809;
srom_1(48790) <= 1706186;
srom_1(48791) <= 2068899;
srom_1(48792) <= 2461248;
srom_1(48793) <= 2881392;
srom_1(48794) <= 3327361;
srom_1(48795) <= 3797064;
srom_1(48796) <= 4288299;
srom_1(48797) <= 4798761;
srom_1(48798) <= 5326057;
srom_1(48799) <= 5867715;
srom_1(48800) <= 6421193;
srom_1(48801) <= 6983898;
srom_1(48802) <= 7553190;
srom_1(48803) <= 8126400;
srom_1(48804) <= 8700839;
srom_1(48805) <= 9273813;
srom_1(48806) <= 9842637;
srom_1(48807) <= 10404643;
srom_1(48808) <= 10957194;
srom_1(48809) <= 11497701;
srom_1(48810) <= 12023628;
srom_1(48811) <= 12532509;
srom_1(48812) <= 13021957;
srom_1(48813) <= 13489679;
srom_1(48814) <= 13933480;
srom_1(48815) <= 14351279;
srom_1(48816) <= 14741117;
srom_1(48817) <= 15101165;
srom_1(48818) <= 15429737;
srom_1(48819) <= 15725290;
srom_1(48820) <= 15986439;
srom_1(48821) <= 16211959;
srom_1(48822) <= 16400792;
srom_1(48823) <= 16552054;
srom_1(48824) <= 16665035;
srom_1(48825) <= 16739204;
srom_1(48826) <= 16774215;
srom_1(48827) <= 16769903;
srom_1(48828) <= 16726287;
srom_1(48829) <= 16643574;
srom_1(48830) <= 16522150;
srom_1(48831) <= 16362586;
srom_1(48832) <= 16165628;
srom_1(48833) <= 15932202;
srom_1(48834) <= 15663401;
srom_1(48835) <= 15360486;
srom_1(48836) <= 15024877;
srom_1(48837) <= 14658149;
srom_1(48838) <= 14262020;
srom_1(48839) <= 13838349;
srom_1(48840) <= 13389123;
srom_1(48841) <= 12916447;
srom_1(48842) <= 12422539;
srom_1(48843) <= 11909714;
srom_1(48844) <= 11380377;
srom_1(48845) <= 10837012;
srom_1(48846) <= 10282164;
srom_1(48847) <= 9718437;
srom_1(48848) <= 9148474;
srom_1(48849) <= 8574948;
srom_1(48850) <= 8000548;
srom_1(48851) <= 7427968;
srom_1(48852) <= 6859892;
srom_1(48853) <= 6298986;
srom_1(48854) <= 5747878;
srom_1(48855) <= 5209153;
srom_1(48856) <= 4685338;
srom_1(48857) <= 4178889;
srom_1(48858) <= 3692180;
srom_1(48859) <= 3227495;
srom_1(48860) <= 2787012;
srom_1(48861) <= 2372797;
srom_1(48862) <= 1986792;
srom_1(48863) <= 1630807;
srom_1(48864) <= 1306512;
srom_1(48865) <= 1015428;
srom_1(48866) <= 758918;
srom_1(48867) <= 538187;
srom_1(48868) <= 354270;
srom_1(48869) <= 208028;
srom_1(48870) <= 100147;
srom_1(48871) <= 31134;
srom_1(48872) <= 1312;
srom_1(48873) <= 10821;
srom_1(48874) <= 59617;
srom_1(48875) <= 147469;
srom_1(48876) <= 273968;
srom_1(48877) <= 438518;
srom_1(48878) <= 640350;
srom_1(48879) <= 878515;
srom_1(48880) <= 1151898;
srom_1(48881) <= 1459216;
srom_1(48882) <= 1799029;
srom_1(48883) <= 2169743;
srom_1(48884) <= 2569618;
srom_1(48885) <= 2996781;
srom_1(48886) <= 3449229;
srom_1(48887) <= 3924838;
srom_1(48888) <= 4421380;
srom_1(48889) <= 4936526;
srom_1(48890) <= 5467859;
srom_1(48891) <= 6012889;
srom_1(48892) <= 6569059;
srom_1(48893) <= 7133762;
srom_1(48894) <= 7704349;
srom_1(48895) <= 8278145;
srom_1(48896) <= 8852459;
srom_1(48897) <= 9424598;
srom_1(48898) <= 9991879;
srom_1(48899) <= 10551641;
srom_1(48900) <= 11101261;
srom_1(48901) <= 11638159;
srom_1(48902) <= 12159820;
srom_1(48903) <= 12663795;
srom_1(48904) <= 13147723;
srom_1(48905) <= 13609334;
srom_1(48906) <= 14046463;
srom_1(48907) <= 14457061;
srom_1(48908) <= 14839201;
srom_1(48909) <= 15191093;
srom_1(48910) <= 15511085;
srom_1(48911) <= 15797677;
srom_1(48912) <= 16049526;
srom_1(48913) <= 16265450;
srom_1(48914) <= 16444437;
srom_1(48915) <= 16585647;
srom_1(48916) <= 16688418;
srom_1(48917) <= 16752269;
srom_1(48918) <= 16776900;
srom_1(48919) <= 16762195;
srom_1(48920) <= 16708224;
srom_1(48921) <= 16615239;
srom_1(48922) <= 16483676;
srom_1(48923) <= 16314153;
srom_1(48924) <= 16107464;
srom_1(48925) <= 15864579;
srom_1(48926) <= 15586637;
srom_1(48927) <= 15274940;
srom_1(48928) <= 14930952;
srom_1(48929) <= 14556283;
srom_1(48930) <= 14152693;
srom_1(48931) <= 13722072;
srom_1(48932) <= 13266442;
srom_1(48933) <= 12787937;
srom_1(48934) <= 12288802;
srom_1(48935) <= 11771378;
srom_1(48936) <= 11238092;
srom_1(48937) <= 10691442;
srom_1(48938) <= 10133994;
srom_1(48939) <= 9568362;
srom_1(48940) <= 8997197;
srom_1(48941) <= 8423178;
srom_1(48942) <= 7848997;
srom_1(48943) <= 7277346;
srom_1(48944) <= 6710907;
srom_1(48945) <= 6152335;
srom_1(48946) <= 5604249;
srom_1(48947) <= 5069221;
srom_1(48948) <= 4549758;
srom_1(48949) <= 4048296;
srom_1(48950) <= 3567188;
srom_1(48951) <= 3108690;
srom_1(48952) <= 2674950;
srom_1(48953) <= 2268004;
srom_1(48954) <= 1889759;
srom_1(48955) <= 1541990;
srom_1(48956) <= 1226327;
srom_1(48957) <= 944250;
srom_1(48958) <= 697083;
srom_1(48959) <= 485984;
srom_1(48960) <= 311942;
srom_1(48961) <= 175775;
srom_1(48962) <= 78121;
srom_1(48963) <= 19438;
srom_1(48964) <= 0;
srom_1(48965) <= 19900;
srom_1(48966) <= 79043;
srom_1(48967) <= 177153;
srom_1(48968) <= 313769;
srom_1(48969) <= 488250;
srom_1(48970) <= 699779;
srom_1(48971) <= 947364;
srom_1(48972) <= 1229843;
srom_1(48973) <= 1545892;
srom_1(48974) <= 1894029;
srom_1(48975) <= 2272622;
srom_1(48976) <= 2679894;
srom_1(48977) <= 3113936;
srom_1(48978) <= 3572713;
srom_1(48979) <= 4054074;
srom_1(48980) <= 4555760;
srom_1(48981) <= 5075420;
srom_1(48982) <= 5610617;
srom_1(48983) <= 6158841;
srom_1(48984) <= 6717521;
srom_1(48985) <= 7284037;
srom_1(48986) <= 7855733;
srom_1(48987) <= 8429927;
srom_1(48988) <= 9003928;
srom_1(48989) <= 9575044;
srom_1(48990) <= 10140596;
srom_1(48991) <= 10697932;
srom_1(48992) <= 11244439;
srom_1(48993) <= 11777554;
srom_1(48994) <= 12294777;
srom_1(48995) <= 12793683;
srom_1(48996) <= 13271931;
srom_1(48997) <= 13727280;
srom_1(48998) <= 14157595;
srom_1(48999) <= 14560856;
srom_1(49000) <= 14935174;
srom_1(49001) <= 15278793;
srom_1(49002) <= 15590101;
srom_1(49003) <= 15867639;
srom_1(49004) <= 16110105;
srom_1(49005) <= 16316362;
srom_1(49006) <= 16485444;
srom_1(49007) <= 16616556;
srom_1(49008) <= 16709085;
srom_1(49009) <= 16762596;
srom_1(49010) <= 16776839;
srom_1(49011) <= 16751746;
srom_1(49012) <= 16687436;
srom_1(49013) <= 16584210;
srom_1(49014) <= 16442552;
srom_1(49015) <= 16263126;
srom_1(49016) <= 16046774;
srom_1(49017) <= 15794510;
srom_1(49018) <= 15507517;
srom_1(49019) <= 15187141;
srom_1(49020) <= 14834884;
srom_1(49021) <= 14452399;
srom_1(49022) <= 14041478;
srom_1(49023) <= 13604049;
srom_1(49024) <= 13142164;
srom_1(49025) <= 12657987;
srom_1(49026) <= 12153789;
srom_1(49027) <= 11631936;
srom_1(49028) <= 11094873;
srom_1(49029) <= 10545119;
srom_1(49030) <= 9985253;
srom_1(49031) <= 9417900;
srom_1(49032) <= 8845720;
srom_1(49033) <= 8271396;
srom_1(49034) <= 7697623;
srom_1(49035) <= 7127089;
srom_1(49036) <= 6562471;
srom_1(49037) <= 6006416;
srom_1(49038) <= 5461533;
srom_1(49039) <= 4930375;
srom_1(49040) <= 4415434;
srom_1(49041) <= 3919125;
srom_1(49042) <= 3443775;
srom_1(49043) <= 2991613;
srom_1(49044) <= 2564759;
srom_1(49045) <= 2165215;
srom_1(49046) <= 1794854;
srom_1(49047) <= 1455415;
srom_1(49048) <= 1148487;
srom_1(49049) <= 875510;
srom_1(49050) <= 637766;
srom_1(49051) <= 436367;
srom_1(49052) <= 272259;
srom_1(49053) <= 146212;
srom_1(49054) <= 58816;
srom_1(49055) <= 10481;
srom_1(49056) <= 1434;
srom_1(49057) <= 31718;
srom_1(49058) <= 101190;
srom_1(49059) <= 209524;
srom_1(49060) <= 356213;
srom_1(49061) <= 540569;
srom_1(49062) <= 761726;
srom_1(49063) <= 1018649;
srom_1(49064) <= 1310132;
srom_1(49065) <= 1634809;
srom_1(49066) <= 1991156;
srom_1(49067) <= 2377503;
srom_1(49068) <= 2792038;
srom_1(49069) <= 3232818;
srom_1(49070) <= 3697775;
srom_1(49071) <= 4184728;
srom_1(49072) <= 4691395;
srom_1(49073) <= 5215400;
srom_1(49074) <= 5754285;
srom_1(49075) <= 6305523;
srom_1(49076) <= 6866529;
srom_1(49077) <= 7434673;
srom_1(49078) <= 8007291;
srom_1(49079) <= 8581696;
srom_1(49080) <= 9155196;
srom_1(49081) <= 9725101;
srom_1(49082) <= 10288739;
srom_1(49083) <= 10843466;
srom_1(49084) <= 11386682;
srom_1(49085) <= 11915839;
srom_1(49086) <= 12428455;
srom_1(49087) <= 12922127;
srom_1(49088) <= 13394540;
srom_1(49089) <= 13843479;
srom_1(49090) <= 14266837;
srom_1(49091) <= 14662631;
srom_1(49092) <= 15029003;
srom_1(49093) <= 15364237;
srom_1(49094) <= 15666759;
srom_1(49095) <= 15935152;
srom_1(49096) <= 16168156;
srom_1(49097) <= 16364679;
srom_1(49098) <= 16523799;
srom_1(49099) <= 16644771;
srom_1(49100) <= 16727027;
srom_1(49101) <= 16770182;
srom_1(49102) <= 16774032;
srom_1(49103) <= 16738560;
srom_1(49104) <= 16663932;
srom_1(49105) <= 16550498;
srom_1(49106) <= 16398791;
srom_1(49107) <= 16209521;
srom_1(49108) <= 15983576;
srom_1(49109) <= 15722015;
srom_1(49110) <= 15426066;
srom_1(49111) <= 15097115;
srom_1(49112) <= 14736706;
srom_1(49113) <= 14346529;
srom_1(49114) <= 13928413;
srom_1(49115) <= 13484319;
srom_1(49116) <= 13016329;
srom_1(49117) <= 12526639;
srom_1(49118) <= 12017543;
srom_1(49119) <= 11491431;
srom_1(49120) <= 10950768;
srom_1(49121) <= 10398090;
srom_1(49122) <= 9835989;
srom_1(49123) <= 9267101;
srom_1(49124) <= 8694094;
srom_1(49125) <= 8119653;
srom_1(49126) <= 7546474;
srom_1(49127) <= 6977244;
srom_1(49128) <= 6414633;
srom_1(49129) <= 5861278;
srom_1(49130) <= 5319774;
srom_1(49131) <= 4792662;
srom_1(49132) <= 4282412;
srom_1(49133) <= 3791417;
srom_1(49134) <= 3321980;
srom_1(49135) <= 2876302;
srom_1(49136) <= 2456474;
srom_1(49137) <= 2064463;
srom_1(49138) <= 1702108;
srom_1(49139) <= 1371109;
srom_1(49140) <= 1073017;
srom_1(49141) <= 809230;
srom_1(49142) <= 580986;
srom_1(49143) <= 389354;
srom_1(49144) <= 235234;
srom_1(49145) <= 119347;
srom_1(49146) <= 42238;
srom_1(49147) <= 4268;
srom_1(49148) <= 5615;
srom_1(49149) <= 46272;
srom_1(49150) <= 126050;
srom_1(49151) <= 244574;
srom_1(49152) <= 401287;
srom_1(49153) <= 595456;
srom_1(49154) <= 826170;
srom_1(49155) <= 1092347;
srom_1(49156) <= 1392738;
srom_1(49157) <= 1725936;
srom_1(49158) <= 2090377;
srom_1(49159) <= 2484352;
srom_1(49160) <= 2906015;
srom_1(49161) <= 3353387;
srom_1(49162) <= 3824372;
srom_1(49163) <= 4316759;
srom_1(49164) <= 4828241;
srom_1(49165) <= 5356418;
srom_1(49166) <= 5898815;
srom_1(49167) <= 6452887;
srom_1(49168) <= 7016036;
srom_1(49169) <= 7585622;
srom_1(49170) <= 8158973;
srom_1(49171) <= 8733401;
srom_1(49172) <= 9306213;
srom_1(49173) <= 9874721;
srom_1(49174) <= 10436260;
srom_1(49175) <= 10988197;
srom_1(49176) <= 11527944;
srom_1(49177) <= 12052969;
srom_1(49178) <= 12560811;
srom_1(49179) <= 13049088;
srom_1(49180) <= 13515511;
srom_1(49181) <= 13957891;
srom_1(49182) <= 14374155;
srom_1(49183) <= 14762351;
srom_1(49184) <= 15120659;
srom_1(49185) <= 15447397;
srom_1(49186) <= 15741035;
srom_1(49187) <= 16000194;
srom_1(49188) <= 16223660;
srom_1(49189) <= 16410384;
srom_1(49190) <= 16559492;
srom_1(49191) <= 16670284;
srom_1(49192) <= 16742240;
srom_1(49193) <= 16775023;
srom_1(49194) <= 16768479;
srom_1(49195) <= 16722639;
srom_1(49196) <= 16637718;
srom_1(49197) <= 16514114;
srom_1(49198) <= 16352407;
srom_1(49199) <= 16153355;
srom_1(49200) <= 15917891;
srom_1(49201) <= 15647120;
srom_1(49202) <= 15342311;
srom_1(49203) <= 15004894;
srom_1(49204) <= 14636450;
srom_1(49205) <= 14238709;
srom_1(49206) <= 13813534;
srom_1(49207) <= 13362920;
srom_1(49208) <= 12888980;
srom_1(49209) <= 12393936;
srom_1(49210) <= 11880109;
srom_1(49211) <= 11349910;
srom_1(49212) <= 10805824;
srom_1(49213) <= 10250403;
srom_1(49214) <= 9686252;
srom_1(49215) <= 9116015;
srom_1(49216) <= 8542367;
srom_1(49217) <= 7967998;
srom_1(49218) <= 7395602;
srom_1(49219) <= 6827862;
srom_1(49220) <= 6267441;
srom_1(49221) <= 5716967;
srom_1(49222) <= 5179021;
srom_1(49223) <= 4656126;
srom_1(49224) <= 4150733;
srom_1(49225) <= 3665214;
srom_1(49226) <= 3201844;
srom_1(49227) <= 2762797;
srom_1(49228) <= 2350131;
srom_1(49229) <= 1965782;
srom_1(49230) <= 1611551;
srom_1(49231) <= 1289101;
srom_1(49232) <= 999942;
srom_1(49233) <= 745431;
srom_1(49234) <= 526762;
srom_1(49235) <= 344960;
srom_1(49236) <= 200877;
srom_1(49237) <= 95189;
srom_1(49238) <= 28392;
srom_1(49239) <= 799;
srom_1(49240) <= 12539;
srom_1(49241) <= 63558;
srom_1(49242) <= 153615;
srom_1(49243) <= 282289;
srom_1(49244) <= 448977;
srom_1(49245) <= 652896;
srom_1(49246) <= 893090;
srom_1(49247) <= 1168434;
srom_1(49248) <= 1477635;
srom_1(49249) <= 1819245;
srom_1(49250) <= 2191660;
srom_1(49251) <= 2593135;
srom_1(49252) <= 3021787;
srom_1(49253) <= 3475605;
srom_1(49254) <= 3952463;
srom_1(49255) <= 4450123;
srom_1(49256) <= 4966252;
srom_1(49257) <= 5498430;
srom_1(49258) <= 6044160;
srom_1(49259) <= 6600885;
srom_1(49260) <= 7165993;
srom_1(49261) <= 7736834;
srom_1(49262) <= 8310731;
srom_1(49263) <= 8884994;
srom_1(49264) <= 9456929;
srom_1(49265) <= 10023854;
srom_1(49266) <= 10583111;
srom_1(49267) <= 11132077;
srom_1(49268) <= 11668178;
srom_1(49269) <= 12188900;
srom_1(49270) <= 12691801;
srom_1(49271) <= 13174523;
srom_1(49272) <= 13634802;
srom_1(49273) <= 14070480;
srom_1(49274) <= 14479514;
srom_1(49275) <= 14859985;
srom_1(49276) <= 15210110;
srom_1(49277) <= 15528247;
srom_1(49278) <= 15812903;
srom_1(49279) <= 16062744;
srom_1(49280) <= 16276599;
srom_1(49281) <= 16453464;
srom_1(49282) <= 16592510;
srom_1(49283) <= 16693085;
srom_1(49284) <= 16754717;
srom_1(49285) <= 16777118;
srom_1(49286) <= 16760183;
srom_1(49287) <= 16703990;
srom_1(49288) <= 16608804;
srom_1(49289) <= 16475070;
srom_1(49290) <= 16303416;
srom_1(49291) <= 16094647;
srom_1(49292) <= 15849741;
srom_1(49293) <= 15569848;
srom_1(49294) <= 15256279;
srom_1(49295) <= 14910506;
srom_1(49296) <= 14534149;
srom_1(49297) <= 14128973;
srom_1(49298) <= 13696879;
srom_1(49299) <= 13239893;
srom_1(49300) <= 12760157;
srom_1(49301) <= 12259922;
srom_1(49302) <= 11741532;
srom_1(49303) <= 11207420;
srom_1(49304) <= 10660089;
srom_1(49305) <= 10102107;
srom_1(49306) <= 9536089;
srom_1(49307) <= 8964690;
srom_1(49308) <= 8390590;
srom_1(49309) <= 7816481;
srom_1(49310) <= 7245054;
srom_1(49311) <= 6678990;
srom_1(49312) <= 6120943;
srom_1(49313) <= 5573530;
srom_1(49314) <= 5039318;
srom_1(49315) <= 4520811;
srom_1(49316) <= 4020443;
srom_1(49317) <= 3540557;
srom_1(49318) <= 3083406;
srom_1(49319) <= 2651133;
srom_1(49320) <= 2245765;
srom_1(49321) <= 1869203;
srom_1(49322) <= 1523213;
srom_1(49323) <= 1209417;
srom_1(49324) <= 929286;
srom_1(49325) <= 684135;
srom_1(49326) <= 475112;
srom_1(49327) <= 303199;
srom_1(49328) <= 169201;
srom_1(49329) <= 73747;
srom_1(49330) <= 17284;
srom_1(49331) <= 77;
srom_1(49332) <= 22206;
srom_1(49333) <= 83569;
srom_1(49334) <= 183876;
srom_1(49335) <= 322659;
srom_1(49336) <= 499265;
srom_1(49337) <= 712868;
srom_1(49338) <= 962464;
srom_1(49339) <= 1246884;
srom_1(49340) <= 1564794;
srom_1(49341) <= 1914704;
srom_1(49342) <= 2294972;
srom_1(49343) <= 2703815;
srom_1(49344) <= 3139315;
srom_1(49345) <= 3599432;
srom_1(49346) <= 4082007;
srom_1(49347) <= 4584776;
srom_1(49348) <= 5105384;
srom_1(49349) <= 5641387;
srom_1(49350) <= 6190273;
srom_1(49351) <= 6749468;
srom_1(49352) <= 7316349;
srom_1(49353) <= 7888259;
srom_1(49354) <= 8462515;
srom_1(49355) <= 9036424;
srom_1(49356) <= 9607295;
srom_1(49357) <= 10172452;
srom_1(49358) <= 10729243;
srom_1(49359) <= 11275058;
srom_1(49360) <= 11807338;
srom_1(49361) <= 12323586;
srom_1(49362) <= 12821382;
srom_1(49363) <= 13298391;
srom_1(49364) <= 13752376;
srom_1(49365) <= 14181209;
srom_1(49366) <= 14582878;
srom_1(49367) <= 14955501;
srom_1(49368) <= 15297328;
srom_1(49369) <= 15606759;
srom_1(49370) <= 15882341;
srom_1(49371) <= 16122782;
srom_1(49372) <= 16326955;
srom_1(49373) <= 16493902;
srom_1(49374) <= 16622841;
srom_1(49375) <= 16713167;
srom_1(49376) <= 16764456;
srom_1(49377) <= 16776468;
srom_1(49378) <= 16749146;
srom_1(49379) <= 16682619;
srom_1(49380) <= 16577198;
srom_1(49381) <= 16433378;
srom_1(49382) <= 16251834;
srom_1(49383) <= 16033416;
srom_1(49384) <= 15779149;
srom_1(49385) <= 15490225;
srom_1(49386) <= 15167999;
srom_1(49387) <= 14813983;
srom_1(49388) <= 14429835;
srom_1(49389) <= 14017358;
srom_1(49390) <= 13578486;
srom_1(49391) <= 13115277;
srom_1(49392) <= 12629903;
srom_1(49393) <= 12124640;
srom_1(49394) <= 11601858;
srom_1(49395) <= 11064007;
srom_1(49396) <= 10513611;
srom_1(49397) <= 9953249;
srom_1(49398) <= 9385551;
srom_1(49399) <= 8813177;
srom_1(49400) <= 8238813;
srom_1(49401) <= 7665151;
srom_1(49402) <= 7094881;
srom_1(49403) <= 6530679;
srom_1(49404) <= 5975188;
srom_1(49405) <= 5431015;
srom_1(49406) <= 4900711;
srom_1(49407) <= 4386764;
srom_1(49408) <= 3891582;
srom_1(49409) <= 3417488;
srom_1(49410) <= 2966706;
srom_1(49411) <= 2541348;
srom_1(49412) <= 2143411;
srom_1(49413) <= 1774759;
srom_1(49414) <= 1437122;
srom_1(49415) <= 1132083;
srom_1(49416) <= 861072;
srom_1(49417) <= 625361;
srom_1(49418) <= 426054;
srom_1(49419) <= 264086;
srom_1(49420) <= 140216;
srom_1(49421) <= 55027;
srom_1(49422) <= 8916;
srom_1(49423) <= 2100;
srom_1(49424) <= 34612;
srom_1(49425) <= 106299;
srom_1(49426) <= 216824;
srom_1(49427) <= 365669;
srom_1(49428) <= 552137;
srom_1(49429) <= 775352;
srom_1(49430) <= 1034269;
srom_1(49431) <= 1327673;
srom_1(49432) <= 1654188;
srom_1(49433) <= 2012283;
srom_1(49434) <= 2400278;
srom_1(49435) <= 2816356;
srom_1(49436) <= 3258563;
srom_1(49437) <= 3724826;
srom_1(49438) <= 4212960;
srom_1(49439) <= 4720675;
srom_1(49440) <= 5245590;
srom_1(49441) <= 5785244;
srom_1(49442) <= 6337106;
srom_1(49443) <= 6898588;
srom_1(49444) <= 7467057;
srom_1(49445) <= 8039848;
srom_1(49446) <= 8614274;
srom_1(49447) <= 9187642;
srom_1(49448) <= 9757262;
srom_1(49449) <= 10320465;
srom_1(49450) <= 10874609;
srom_1(49451) <= 11417095;
srom_1(49452) <= 11945379;
srom_1(49453) <= 12456985;
srom_1(49454) <= 12949512;
srom_1(49455) <= 13420652;
srom_1(49456) <= 13868195;
srom_1(49457) <= 14290042;
srom_1(49458) <= 14684215;
srom_1(49459) <= 15048866;
srom_1(49460) <= 15382284;
srom_1(49461) <= 15682907;
srom_1(49462) <= 15949325;
srom_1(49463) <= 16180288;
srom_1(49464) <= 16374712;
srom_1(49465) <= 16531688;
srom_1(49466) <= 16650477;
srom_1(49467) <= 16730524;
srom_1(49468) <= 16771452;
srom_1(49469) <= 16773071;
srom_1(49470) <= 16735372;
srom_1(49471) <= 16658532;
srom_1(49472) <= 16542912;
srom_1(49473) <= 16389053;
srom_1(49474) <= 16197677;
srom_1(49475) <= 15969682;
srom_1(49476) <= 15706137;
srom_1(49477) <= 15408277;
srom_1(49478) <= 15077500;
srom_1(49479) <= 14715356;
srom_1(49480) <= 14323544;
srom_1(49481) <= 13903901;
srom_1(49482) <= 13458394;
srom_1(49483) <= 12989114;
srom_1(49484) <= 12498261;
srom_1(49485) <= 11988135;
srom_1(49486) <= 11461131;
srom_1(49487) <= 10919718;
srom_1(49488) <= 10366436;
srom_1(49489) <= 9803879;
srom_1(49490) <= 9234686;
srom_1(49491) <= 8661525;
srom_1(49492) <= 8087084;
srom_1(49493) <= 7514058;
srom_1(49494) <= 6945132;
srom_1(49495) <= 6382975;
srom_1(49496) <= 5830223;
srom_1(49497) <= 5289469;
srom_1(49498) <= 4763247;
srom_1(49499) <= 4254026;
srom_1(49500) <= 3764193;
srom_1(49501) <= 3296046;
srom_1(49502) <= 2851780;
srom_1(49503) <= 2433477;
srom_1(49504) <= 2043101;
srom_1(49505) <= 1682480;
srom_1(49506) <= 1353307;
srom_1(49507) <= 1057125;
srom_1(49508) <= 795323;
srom_1(49509) <= 569128;
srom_1(49510) <= 379601;
srom_1(49511) <= 227632;
srom_1(49512) <= 113932;
srom_1(49513) <= 39035;
srom_1(49514) <= 3292;
srom_1(49515) <= 6870;
srom_1(49516) <= 49753;
srom_1(49517) <= 131740;
srom_1(49518) <= 252447;
srom_1(49519) <= 411306;
srom_1(49520) <= 607574;
srom_1(49521) <= 840330;
srom_1(49522) <= 1108482;
srom_1(49523) <= 1410773;
srom_1(49524) <= 1745786;
srom_1(49525) <= 2111949;
srom_1(49526) <= 2507546;
srom_1(49527) <= 2930721;
srom_1(49528) <= 3379490;
srom_1(49529) <= 3851748;
srom_1(49530) <= 4345281;
srom_1(49531) <= 4857775;
srom_1(49532) <= 5386826;
srom_1(49533) <= 5929953;
srom_1(49534) <= 6484610;
srom_1(49535) <= 7048195;
srom_1(49536) <= 7618066;
srom_1(49537) <= 8191551;
srom_1(49538) <= 8765959;
srom_1(49539) <= 9338598;
srom_1(49540) <= 9906782;
srom_1(49541) <= 10467847;
srom_1(49542) <= 11019161;
srom_1(49543) <= 11558140;
srom_1(49544) <= 12082256;
srom_1(49545) <= 12589051;
srom_1(49546) <= 13076149;
srom_1(49547) <= 13541265;
srom_1(49548) <= 13982219;
srom_1(49549) <= 14396942;
srom_1(49550) <= 14783490;
srom_1(49551) <= 15140051;
srom_1(49552) <= 15464951;
srom_1(49553) <= 15756668;
srom_1(49554) <= 16013834;
srom_1(49555) <= 16235242;
srom_1(49556) <= 16419855;
srom_1(49557) <= 16566807;
srom_1(49558) <= 16675408;
srom_1(49559) <= 16745149;
srom_1(49560) <= 16775704;
srom_1(49561) <= 16766929;
srom_1(49562) <= 16718865;
srom_1(49563) <= 16631738;
srom_1(49564) <= 16505955;
srom_1(49565) <= 16342108;
srom_1(49566) <= 16140964;
srom_1(49567) <= 15903466;
srom_1(49568) <= 15630729;
srom_1(49569) <= 15324031;
srom_1(49570) <= 14984810;
srom_1(49571) <= 14614658;
srom_1(49572) <= 14215309;
srom_1(49573) <= 13788637;
srom_1(49574) <= 13336643;
srom_1(49575) <= 12861445;
srom_1(49576) <= 12365272;
srom_1(49577) <= 11850452;
srom_1(49578) <= 11319398;
srom_1(49579) <= 10774601;
srom_1(49580) <= 10218614;
srom_1(49581) <= 9654046;
srom_1(49582) <= 9083544;
srom_1(49583) <= 8509784;
srom_1(49584) <= 7935455;
srom_1(49585) <= 7363251;
srom_1(49586) <= 6795855;
srom_1(49587) <= 6235928;
srom_1(49588) <= 5686096;
srom_1(49589) <= 5148937;
srom_1(49590) <= 4626970;
srom_1(49591) <= 4122642;
srom_1(49592) <= 3638319;
srom_1(49593) <= 3176272;
srom_1(49594) <= 2738667;
srom_1(49595) <= 2327556;
srom_1(49596) <= 1944868;
srom_1(49597) <= 1592397;
srom_1(49598) <= 1271796;
srom_1(49599) <= 984568;
srom_1(49600) <= 732059;
srom_1(49601) <= 515456;
srom_1(49602) <= 335772;
srom_1(49603) <= 193850;
srom_1(49604) <= 90357;
srom_1(49605) <= 25776;
srom_1(49606) <= 412;
srom_1(49607) <= 14384;
srom_1(49608) <= 67624;
srom_1(49609) <= 159885;
srom_1(49610) <= 290733;
srom_1(49611) <= 459555;
srom_1(49612) <= 665559;
srom_1(49613) <= 907778;
srom_1(49614) <= 1185078;
srom_1(49615) <= 1496158;
srom_1(49616) <= 1839559;
srom_1(49617) <= 2213671;
srom_1(49618) <= 2616739;
srom_1(49619) <= 3046873;
srom_1(49620) <= 3502056;
srom_1(49621) <= 3980155;
srom_1(49622) <= 4478925;
srom_1(49623) <= 4996030;
srom_1(49624) <= 5529044;
srom_1(49625) <= 6075467;
srom_1(49626) <= 6632737;
srom_1(49627) <= 7198242;
srom_1(49628) <= 7769328;
srom_1(49629) <= 8343318;
srom_1(49630) <= 8917521;
srom_1(49631) <= 9489243;
srom_1(49632) <= 10055804;
srom_1(49633) <= 10614547;
srom_1(49634) <= 11162852;
srom_1(49635) <= 11698147;
srom_1(49636) <= 12217923;
srom_1(49637) <= 12719742;
srom_1(49638) <= 13201251;
srom_1(49639) <= 13660191;
srom_1(49640) <= 14094411;
srom_1(49641) <= 14501875;
srom_1(49642) <= 14880672;
srom_1(49643) <= 15229025;
srom_1(49644) <= 15545301;
srom_1(49645) <= 15828017;
srom_1(49646) <= 16075846;
srom_1(49647) <= 16287628;
srom_1(49648) <= 16462369;
srom_1(49649) <= 16599248;
srom_1(49650) <= 16697626;
srom_1(49651) <= 16757039;
srom_1(49652) <= 16777210;
srom_1(49653) <= 16758044;
srom_1(49654) <= 16699631;
srom_1(49655) <= 16602245;
srom_1(49656) <= 16466342;
srom_1(49657) <= 16292559;
srom_1(49658) <= 16081713;
srom_1(49659) <= 15834790;
srom_1(49660) <= 15552950;
srom_1(49661) <= 15237514;
srom_1(49662) <= 14889961;
srom_1(49663) <= 14511921;
srom_1(49664) <= 14105167;
srom_1(49665) <= 13671606;
srom_1(49666) <= 13213271;
srom_1(49667) <= 12732311;
srom_1(49668) <= 12230983;
srom_1(49669) <= 11711636;
srom_1(49670) <= 11176706;
srom_1(49671) <= 10628702;
srom_1(49672) <= 10070193;
srom_1(49673) <= 9503799;
srom_1(49674) <= 8932175;
srom_1(49675) <= 8358002;
srom_1(49676) <= 7783973;
srom_1(49677) <= 7212779;
srom_1(49678) <= 6647099;
srom_1(49679) <= 6089586;
srom_1(49680) <= 5542853;
srom_1(49681) <= 5009465;
srom_1(49682) <= 4491924;
srom_1(49683) <= 3992655;
srom_1(49684) <= 3514000;
srom_1(49685) <= 3058203;
srom_1(49686) <= 2627403;
srom_1(49687) <= 2223620;
srom_1(49688) <= 1848745;
srom_1(49689) <= 1504539;
srom_1(49690) <= 1192614;
srom_1(49691) <= 914434;
srom_1(49692) <= 671303;
srom_1(49693) <= 464361;
srom_1(49694) <= 294578;
srom_1(49695) <= 162751;
srom_1(49696) <= 69498;
srom_1(49697) <= 15256;
srom_1(49698) <= 280;
srom_1(49699) <= 24639;
srom_1(49700) <= 88220;
srom_1(49701) <= 190724;
srom_1(49702) <= 331671;
srom_1(49703) <= 510399;
srom_1(49704) <= 726072;
srom_1(49705) <= 977676;
srom_1(49706) <= 1264033;
srom_1(49707) <= 1583800;
srom_1(49708) <= 1935476;
srom_1(49709) <= 2317414;
srom_1(49710) <= 2727821;
srom_1(49711) <= 3164774;
srom_1(49712) <= 3626223;
srom_1(49713) <= 4110005;
srom_1(49714) <= 4613850;
srom_1(49715) <= 5135397;
srom_1(49716) <= 5672198;
srom_1(49717) <= 6221739;
srom_1(49718) <= 6781440;
srom_1(49719) <= 7348678;
srom_1(49720) <= 7920792;
srom_1(49721) <= 8495100;
srom_1(49722) <= 9068909;
srom_1(49723) <= 9639528;
srom_1(49724) <= 10204281;
srom_1(49725) <= 10760519;
srom_1(49726) <= 11305634;
srom_1(49727) <= 11837071;
srom_1(49728) <= 12352337;
srom_1(49729) <= 12849015;
srom_1(49730) <= 13324777;
srom_1(49731) <= 13777392;
srom_1(49732) <= 14204736;
srom_1(49733) <= 14604807;
srom_1(49734) <= 14975728;
srom_1(49735) <= 15315760;
srom_1(49736) <= 15623308;
srom_1(49737) <= 15896929;
srom_1(49738) <= 16135342;
srom_1(49739) <= 16337428;
srom_1(49740) <= 16502239;
srom_1(49741) <= 16629002;
srom_1(49742) <= 16717123;
srom_1(49743) <= 16766189;
srom_1(49744) <= 16775970;
srom_1(49745) <= 16746419;
srom_1(49746) <= 16677676;
srom_1(49747) <= 16570062;
srom_1(49748) <= 16424083;
srom_1(49749) <= 16240423;
srom_1(49750) <= 16019943;
srom_1(49751) <= 15763677;
srom_1(49752) <= 15472826;
srom_1(49753) <= 15148755;
srom_1(49754) <= 14792984;
srom_1(49755) <= 14407180;
srom_1(49756) <= 13993153;
srom_1(49757) <= 13552845;
srom_1(49758) <= 13088319;
srom_1(49759) <= 12601755;
srom_1(49760) <= 12095435;
srom_1(49761) <= 11571731;
srom_1(49762) <= 11033101;
srom_1(49763) <= 10482070;
srom_1(49764) <= 9921222;
srom_1(49765) <= 9353186;
srom_1(49766) <= 8780628;
srom_1(49767) <= 8206231;
srom_1(49768) <= 7632690;
srom_1(49769) <= 7062693;
srom_1(49770) <= 6498914;
srom_1(49771) <= 5943996;
srom_1(49772) <= 5400542;
srom_1(49773) <= 4871101;
srom_1(49774) <= 4358153;
srom_1(49775) <= 3864106;
srom_1(49776) <= 3391276;
srom_1(49777) <= 2941880;
srom_1(49778) <= 2518026;
srom_1(49779) <= 2121701;
srom_1(49780) <= 1754764;
srom_1(49781) <= 1418935;
srom_1(49782) <= 1115789;
srom_1(49783) <= 846748;
srom_1(49784) <= 613073;
srom_1(49785) <= 415860;
srom_1(49786) <= 256034;
srom_1(49787) <= 134345;
srom_1(49788) <= 51363;
srom_1(49789) <= 7477;
srom_1(49790) <= 2893;
srom_1(49791) <= 37633;
srom_1(49792) <= 111533;
srom_1(49793) <= 224247;
srom_1(49794) <= 375246;
srom_1(49795) <= 563823;
srom_1(49796) <= 789093;
srom_1(49797) <= 1050000;
srom_1(49798) <= 1345320;
srom_1(49799) <= 1673669;
srom_1(49800) <= 2033506;
srom_1(49801) <= 2423144;
srom_1(49802) <= 2840757;
srom_1(49803) <= 3284385;
srom_1(49804) <= 3751949;
srom_1(49805) <= 4241255;
srom_1(49806) <= 4750010;
srom_1(49807) <= 5275828;
srom_1(49808) <= 5816242;
srom_1(49809) <= 6368719;
srom_1(49810) <= 6930669;
srom_1(49811) <= 7499454;
srom_1(49812) <= 8072410;
srom_1(49813) <= 8646848;
srom_1(49814) <= 9220075;
srom_1(49815) <= 9789403;
srom_1(49816) <= 10352163;
srom_1(49817) <= 10905714;
srom_1(49818) <= 11447462;
srom_1(49819) <= 11974866;
srom_1(49820) <= 12485453;
srom_1(49821) <= 12976828;
srom_1(49822) <= 13446687;
srom_1(49823) <= 13892828;
srom_1(49824) <= 14313157;
srom_1(49825) <= 14705704;
srom_1(49826) <= 15068628;
srom_1(49827) <= 15400227;
srom_1(49828) <= 15698946;
srom_1(49829) <= 15963384;
srom_1(49830) <= 16192302;
srom_1(49831) <= 16384625;
srom_1(49832) <= 16539453;
srom_1(49833) <= 16656058;
srom_1(49834) <= 16733894;
srom_1(49835) <= 16772597;
srom_1(49836) <= 16771984;
srom_1(49837) <= 16732058;
srom_1(49838) <= 16653007;
srom_1(49839) <= 16535202;
srom_1(49840) <= 16379194;
srom_1(49841) <= 16185716;
srom_1(49842) <= 15955674;
srom_1(49843) <= 15690148;
srom_1(49844) <= 15390383;
srom_1(49845) <= 15057783;
srom_1(49846) <= 14693910;
srom_1(49847) <= 14300469;
srom_1(49848) <= 13879305;
srom_1(49849) <= 13432393;
srom_1(49850) <= 12961830;
srom_1(49851) <= 12469820;
srom_1(49852) <= 11958673;
srom_1(49853) <= 11430784;
srom_1(49854) <= 10888630;
srom_1(49855) <= 10334752;
srom_1(49856) <= 9771748;
srom_1(49857) <= 9202258;
srom_1(49858) <= 8628953;
srom_1(49859) <= 8054520;
srom_1(49860) <= 7481654;
srom_1(49861) <= 6913041;
srom_1(49862) <= 6351347;
srom_1(49863) <= 5799207;
srom_1(49864) <= 5259210;
srom_1(49865) <= 4733887;
srom_1(49866) <= 4225703;
srom_1(49867) <= 3737039;
srom_1(49868) <= 3270189;
srom_1(49869) <= 2827341;
srom_1(49870) <= 2410571;
srom_1(49871) <= 2021834;
srom_1(49872) <= 1662954;
srom_1(49873) <= 1335612;
srom_1(49874) <= 1041344;
srom_1(49875) <= 781530;
srom_1(49876) <= 557388;
srom_1(49877) <= 369970;
srom_1(49878) <= 220153;
srom_1(49879) <= 108642;
srom_1(49880) <= 35958;
srom_1(49881) <= 2442;
srom_1(49882) <= 8252;
srom_1(49883) <= 53360;
srom_1(49884) <= 137555;
srom_1(49885) <= 260442;
srom_1(49886) <= 421445;
srom_1(49887) <= 619809;
srom_1(49888) <= 854603;
srom_1(49889) <= 1124727;
srom_1(49890) <= 1428914;
srom_1(49891) <= 1765737;
srom_1(49892) <= 2133616;
srom_1(49893) <= 2530828;
srom_1(49894) <= 2955509;
srom_1(49895) <= 3405667;
srom_1(49896) <= 3879193;
srom_1(49897) <= 4373864;
srom_1(49898) <= 4887362;
srom_1(49899) <= 5417278;
srom_1(49900) <= 5961128;
srom_1(49901) <= 6516362;
srom_1(49902) <= 7080374;
srom_1(49903) <= 7650522;
srom_1(49904) <= 8224131;
srom_1(49905) <= 8798511;
srom_1(49906) <= 9370969;
srom_1(49907) <= 9938820;
srom_1(49908) <= 10499402;
srom_1(49909) <= 11050085;
srom_1(49910) <= 11588288;
srom_1(49911) <= 12111487;
srom_1(49912) <= 12617227;
srom_1(49913) <= 13103138;
srom_1(49914) <= 13566942;
srom_1(49915) <= 14006462;
srom_1(49916) <= 14419638;
srom_1(49917) <= 14804532;
srom_1(49918) <= 15159340;
srom_1(49919) <= 15482398;
srom_1(49920) <= 15772191;
srom_1(49921) <= 16027359;
srom_1(49922) <= 16246707;
srom_1(49923) <= 16429205;
srom_1(49924) <= 16573998;
srom_1(49925) <= 16680407;
srom_1(49926) <= 16747933;
srom_1(49927) <= 16776259;
srom_1(49928) <= 16765253;
srom_1(49929) <= 16714965;
srom_1(49930) <= 16625633;
srom_1(49931) <= 16497674;
srom_1(49932) <= 16331689;
srom_1(49933) <= 16128456;
srom_1(49934) <= 15888929;
srom_1(49935) <= 15614229;
srom_1(49936) <= 15305647;
srom_1(49937) <= 14964628;
srom_1(49938) <= 14592771;
srom_1(49939) <= 14191822;
srom_1(49940) <= 13763659;
srom_1(49941) <= 13310290;
srom_1(49942) <= 12833842;
srom_1(49943) <= 12336549;
srom_1(49944) <= 11820743;
srom_1(49945) <= 11288842;
srom_1(49946) <= 10743341;
srom_1(49947) <= 10186798;
srom_1(49948) <= 9621822;
srom_1(49949) <= 9051063;
srom_1(49950) <= 8477198;
srom_1(49951) <= 7902918;
srom_1(49952) <= 7330915;
srom_1(49953) <= 6763872;
srom_1(49954) <= 6204448;
srom_1(49955) <= 5655266;
srom_1(49956) <= 5118902;
srom_1(49957) <= 4597870;
srom_1(49958) <= 4094615;
srom_1(49959) <= 3611495;
srom_1(49960) <= 3150778;
srom_1(49961) <= 2714622;
srom_1(49962) <= 2305073;
srom_1(49963) <= 1924052;
srom_1(49964) <= 1573346;
srom_1(49965) <= 1254598;
srom_1(49966) <= 969305;
srom_1(49967) <= 718803;
srom_1(49968) <= 504268;
srom_1(49969) <= 326705;
srom_1(49970) <= 186947;
srom_1(49971) <= 85649;
srom_1(49972) <= 23287;
srom_1(49973) <= 152;
srom_1(49974) <= 16354;
srom_1(49975) <= 71817;
srom_1(49976) <= 166279;
srom_1(49977) <= 299299;
srom_1(49978) <= 470253;
srom_1(49979) <= 678338;
srom_1(49980) <= 922580;
srom_1(49981) <= 1201832;
srom_1(49982) <= 1514785;
srom_1(49983) <= 1859972;
srom_1(49984) <= 2235775;
srom_1(49985) <= 2640430;
srom_1(49986) <= 3072040;
srom_1(49987) <= 3528581;
srom_1(49988) <= 4007913;
srom_1(49989) <= 4507787;
srom_1(49990) <= 5025860;
srom_1(49991) <= 5559701;
srom_1(49992) <= 6106809;
srom_1(49993) <= 6664617;
srom_1(49994) <= 7230509;
srom_1(49995) <= 7801831;
srom_1(49996) <= 8375906;
srom_1(49997) <= 8950040;
srom_1(49998) <= 9521541;
srom_1(49999) <= 10087729;
srom_1(50000) <= 10645950;
srom_1(50001) <= 11193585;
srom_1(50002) <= 11728067;
srom_1(50003) <= 12246889;
srom_1(50004) <= 12747618;
srom_1(50005) <= 13227906;
srom_1(50006) <= 13685501;
srom_1(50007) <= 14118257;
srom_1(50008) <= 14524144;
srom_1(50009) <= 14901260;
srom_1(50010) <= 15247836;
srom_1(50011) <= 15562247;
srom_1(50012) <= 15843018;
srom_1(50013) <= 16088833;
srom_1(50014) <= 16298539;
srom_1(50015) <= 16471152;
srom_1(50016) <= 16605863;
srom_1(50017) <= 16702041;
srom_1(50018) <= 16759235;
srom_1(50019) <= 16777176;
srom_1(50020) <= 16755779;
srom_1(50021) <= 16695147;
srom_1(50022) <= 16595562;
srom_1(50023) <= 16457491;
srom_1(50024) <= 16281583;
srom_1(50025) <= 16068663;
srom_1(50026) <= 15819727;
srom_1(50027) <= 15535945;
srom_1(50028) <= 15218646;
srom_1(50029) <= 14869319;
srom_1(50030) <= 14489602;
srom_1(50031) <= 14081275;
srom_1(50032) <= 13646253;
srom_1(50033) <= 13186576;
srom_1(50034) <= 12704400;
srom_1(50035) <= 12201985;
srom_1(50036) <= 11681689;
srom_1(50037) <= 11145950;
srom_1(50038) <= 10597281;
srom_1(50039) <= 10038254;
srom_1(50040) <= 9471492;
srom_1(50041) <= 8899652;
srom_1(50042) <= 8325415;
srom_1(50043) <= 7751475;
srom_1(50044) <= 7180522;
srom_1(50045) <= 6615235;
srom_1(50046) <= 6058263;
srom_1(50047) <= 5512220;
srom_1(50048) <= 4979664;
srom_1(50049) <= 4463095;
srom_1(50050) <= 3964933;
srom_1(50051) <= 3487515;
srom_1(50052) <= 3033081;
srom_1(50053) <= 2603760;
srom_1(50054) <= 2201567;
srom_1(50055) <= 1828386;
srom_1(50056) <= 1485969;
srom_1(50057) <= 1175921;
srom_1(50058) <= 899695;
srom_1(50059) <= 658587;
srom_1(50060) <= 453729;
srom_1(50061) <= 286079;
srom_1(50062) <= 156425;
srom_1(50063) <= 65375;
srom_1(50064) <= 13355;
srom_1(50065) <= 609;
srom_1(50066) <= 27198;
srom_1(50067) <= 92996;
srom_1(50068) <= 197695;
srom_1(50069) <= 340804;
srom_1(50070) <= 521653;
srom_1(50071) <= 739391;
srom_1(50072) <= 993000;
srom_1(50073) <= 1281289;
srom_1(50074) <= 1602907;
srom_1(50075) <= 1956346;
srom_1(50076) <= 2339947;
srom_1(50077) <= 2751913;
srom_1(50078) <= 3190311;
srom_1(50079) <= 3653086;
srom_1(50080) <= 4138067;
srom_1(50081) <= 4642980;
srom_1(50082) <= 5165458;
srom_1(50083) <= 5703051;
srom_1(50084) <= 6253237;
srom_1(50085) <= 6813436;
srom_1(50086) <= 7381022;
srom_1(50087) <= 7953333;
srom_1(50088) <= 8527685;
srom_1(50089) <= 9101385;
srom_1(50090) <= 9671742;
srom_1(50091) <= 10236082;
srom_1(50092) <= 10791759;
srom_1(50093) <= 11336166;
srom_1(50094) <= 11866752;
srom_1(50095) <= 12381027;
srom_1(50096) <= 12876581;
srom_1(50097) <= 13351088;
srom_1(50098) <= 13802325;
srom_1(50099) <= 14228176;
srom_1(50100) <= 14626642;
srom_1(50101) <= 14995856;
srom_1(50102) <= 15334087;
srom_1(50103) <= 15639747;
srom_1(50104) <= 15911405;
srom_1(50105) <= 16147786;
srom_1(50106) <= 16347781;
srom_1(50107) <= 16510453;
srom_1(50108) <= 16635039;
srom_1(50109) <= 16720954;
srom_1(50110) <= 16767796;
srom_1(50111) <= 16775346;
srom_1(50112) <= 16743567;
srom_1(50113) <= 16672608;
srom_1(50114) <= 16562803;
srom_1(50115) <= 16414667;
srom_1(50116) <= 16228894;
srom_1(50117) <= 16006354;
srom_1(50118) <= 15748093;
srom_1(50119) <= 15455320;
srom_1(50120) <= 15129410;
srom_1(50121) <= 14771889;
srom_1(50122) <= 14384435;
srom_1(50123) <= 13968864;
srom_1(50124) <= 13527126;
srom_1(50125) <= 13061291;
srom_1(50126) <= 12573544;
srom_1(50127) <= 12066173;
srom_1(50128) <= 11541557;
srom_1(50129) <= 11002155;
srom_1(50130) <= 10450497;
srom_1(50131) <= 9889171;
srom_1(50132) <= 9320808;
srom_1(50133) <= 8748073;
srom_1(50134) <= 8173653;
srom_1(50135) <= 7600240;
srom_1(50136) <= 7030525;
srom_1(50137) <= 6467178;
srom_1(50138) <= 5912842;
srom_1(50139) <= 5370115;
srom_1(50140) <= 4841543;
srom_1(50141) <= 4329604;
srom_1(50142) <= 3836699;
srom_1(50143) <= 3365140;
srom_1(50144) <= 2917138;
srom_1(50145) <= 2494793;
srom_1(50146) <= 2100086;
srom_1(50147) <= 1734868;
srom_1(50148) <= 1400852;
srom_1(50149) <= 1099604;
srom_1(50150) <= 832537;
srom_1(50151) <= 600902;
srom_1(50152) <= 405787;
srom_1(50153) <= 248106;
srom_1(50154) <= 128599;
srom_1(50155) <= 47825;
srom_1(50156) <= 6165;
srom_1(50157) <= 3812;
srom_1(50158) <= 40779;
srom_1(50159) <= 116891;
srom_1(50160) <= 231793;
srom_1(50161) <= 384944;
srom_1(50162) <= 575628;
srom_1(50163) <= 802949;
srom_1(50164) <= 1065842;
srom_1(50165) <= 1363074;
srom_1(50166) <= 1693251;
srom_1(50167) <= 2054825;
srom_1(50168) <= 2446100;
srom_1(50169) <= 2865242;
srom_1(50170) <= 3310284;
srom_1(50171) <= 3779141;
srom_1(50172) <= 4269613;
srom_1(50173) <= 4779400;
srom_1(50174) <= 5306112;
srom_1(50175) <= 5847279;
srom_1(50176) <= 6400364;
srom_1(50177) <= 6962771;
srom_1(50178) <= 7531865;
srom_1(50179) <= 8104977;
srom_1(50180) <= 8679418;
srom_1(50181) <= 9252496;
srom_1(50182) <= 9821523;
srom_1(50183) <= 10383830;
srom_1(50184) <= 10936781;
srom_1(50185) <= 11477783;
srom_1(50186) <= 12004298;
srom_1(50187) <= 12513859;
srom_1(50188) <= 13004074;
srom_1(50189) <= 13472646;
srom_1(50190) <= 13917378;
srom_1(50191) <= 14336183;
srom_1(50192) <= 14727097;
srom_1(50193) <= 15088289;
srom_1(50194) <= 15418063;
srom_1(50195) <= 15714874;
srom_1(50196) <= 15977329;
srom_1(50197) <= 16204198;
srom_1(50198) <= 16394418;
srom_1(50199) <= 16547095;
srom_1(50200) <= 16661514;
srom_1(50201) <= 16737139;
srom_1(50202) <= 16773614;
srom_1(50203) <= 16770770;
srom_1(50204) <= 16728618;
srom_1(50205) <= 16647358;
srom_1(50206) <= 16527369;
srom_1(50207) <= 16369215;
srom_1(50208) <= 16173637;
srom_1(50209) <= 15941552;
srom_1(50210) <= 15674049;
srom_1(50211) <= 15372382;
srom_1(50212) <= 15037966;
srom_1(50213) <= 14672369;
srom_1(50214) <= 14277305;
srom_1(50215) <= 13854626;
srom_1(50216) <= 13406316;
srom_1(50217) <= 12934476;
srom_1(50218) <= 12441319;
srom_1(50219) <= 11929157;
srom_1(50220) <= 11400392;
srom_1(50221) <= 10857504;
srom_1(50222) <= 10303039;
srom_1(50223) <= 9739596;
srom_1(50224) <= 9169818;
srom_1(50225) <= 8596376;
srom_1(50226) <= 8021961;
srom_1(50227) <= 7449264;
srom_1(50228) <= 6880973;
srom_1(50229) <= 6319751;
srom_1(50230) <= 5768231;
srom_1(50231) <= 5228998;
srom_1(50232) <= 4704582;
srom_1(50233) <= 4197442;
srom_1(50234) <= 3709956;
srom_1(50235) <= 3244409;
srom_1(50236) <= 2802986;
srom_1(50237) <= 2387755;
srom_1(50238) <= 2000664;
srom_1(50239) <= 1643529;
srom_1(50240) <= 1318023;
srom_1(50241) <= 1025674;
srom_1(50242) <= 767852;
srom_1(50243) <= 545767;
srom_1(50244) <= 360459;
srom_1(50245) <= 212798;
srom_1(50246) <= 103476;
srom_1(50247) <= 33007;
srom_1(50248) <= 1719;
srom_1(50249) <= 9760;
srom_1(50250) <= 57093;
srom_1(50251) <= 143495;
srom_1(50252) <= 268561;
srom_1(50253) <= 431705;
srom_1(50254) <= 632161;
srom_1(50255) <= 868990;
srom_1(50256) <= 1141081;
srom_1(50257) <= 1447159;
srom_1(50258) <= 1785787;
srom_1(50259) <= 2155378;
srom_1(50260) <= 2554199;
srom_1(50261) <= 2980379;
srom_1(50262) <= 3431920;
srom_1(50263) <= 3906705;
srom_1(50264) <= 4402507;
srom_1(50265) <= 4917002;
srom_1(50266) <= 5447776;
srom_1(50267) <= 5992340;
srom_1(50268) <= 6548141;
srom_1(50269) <= 7112573;
srom_1(50270) <= 7682989;
srom_1(50271) <= 8256714;
srom_1(50272) <= 8831057;
srom_1(50273) <= 9403325;
srom_1(50274) <= 9970835;
srom_1(50275) <= 10530925;
srom_1(50276) <= 11080969;
srom_1(50277) <= 11618388;
srom_1(50278) <= 12140661;
srom_1(50279) <= 12645340;
srom_1(50280) <= 13130057;
srom_1(50281) <= 13592540;
srom_1(50282) <= 14030620;
srom_1(50283) <= 14442243;
srom_1(50284) <= 14825478;
srom_1(50285) <= 15178528;
srom_1(50286) <= 15499738;
srom_1(50287) <= 15787602;
srom_1(50288) <= 16040769;
srom_1(50289) <= 16258052;
srom_1(50290) <= 16438433;
srom_1(50291) <= 16581066;
srom_1(50292) <= 16685281;
srom_1(50293) <= 16750590;
srom_1(50294) <= 16776687;
srom_1(50295) <= 16763450;
srom_1(50296) <= 16710940;
srom_1(50297) <= 16619404;
srom_1(50298) <= 16489270;
srom_1(50299) <= 16321150;
srom_1(50300) <= 16115832;
srom_1(50301) <= 15874278;
srom_1(50302) <= 15597620;
srom_1(50303) <= 15287158;
srom_1(50304) <= 14944346;
srom_1(50305) <= 14570791;
srom_1(50306) <= 14168247;
srom_1(50307) <= 13738599;
srom_1(50308) <= 13283864;
srom_1(50309) <= 12806173;
srom_1(50310) <= 12307766;
srom_1(50311) <= 11790981;
srom_1(50312) <= 11258242;
srom_1(50313) <= 10712045;
srom_1(50314) <= 10154954;
srom_1(50315) <= 9589579;
srom_1(50316) <= 9018572;
srom_1(50317) <= 8444612;
srom_1(50318) <= 7870388;
srom_1(50319) <= 7298595;
srom_1(50320) <= 6731914;
srom_1(50321) <= 6173001;
srom_1(50322) <= 5624477;
srom_1(50323) <= 5088916;
srom_1(50324) <= 4568828;
srom_1(50325) <= 4066653;
srom_1(50326) <= 3584744;
srom_1(50327) <= 3125363;
srom_1(50328) <= 2690662;
srom_1(50329) <= 2282681;
srom_1(50330) <= 1903333;
srom_1(50331) <= 1554397;
srom_1(50332) <= 1237509;
srom_1(50333) <= 954154;
srom_1(50334) <= 705663;
srom_1(50335) <= 493199;
srom_1(50336) <= 317760;
srom_1(50337) <= 180167;
srom_1(50338) <= 81067;
srom_1(50339) <= 20923;
srom_1(50340) <= 19;
srom_1(50341) <= 18451;
srom_1(50342) <= 76135;
srom_1(50343) <= 172798;
srom_1(50344) <= 307987;
srom_1(50345) <= 481070;
srom_1(50346) <= 691234;
srom_1(50347) <= 937493;
srom_1(50348) <= 1218694;
srom_1(50349) <= 1533516;
srom_1(50350) <= 1880484;
srom_1(50351) <= 2257972;
srom_1(50352) <= 2664207;
srom_1(50353) <= 3097287;
srom_1(50354) <= 3555179;
srom_1(50355) <= 4035737;
srom_1(50356) <= 4536707;
srom_1(50357) <= 5055740;
srom_1(50358) <= 5590402;
srom_1(50359) <= 6138185;
srom_1(50360) <= 6696522;
srom_1(50361) <= 7262793;
srom_1(50362) <= 7834344;
srom_1(50363) <= 8408494;
srom_1(50364) <= 8982550;
srom_1(50365) <= 9553821;
srom_1(50366) <= 10119629;
srom_1(50367) <= 10677318;
srom_1(50368) <= 11224276;
srom_1(50369) <= 11757936;
srom_1(50370) <= 12275796;
srom_1(50371) <= 12775427;
srom_1(50372) <= 13254487;
srom_1(50373) <= 13710730;
srom_1(50374) <= 14142015;
srom_1(50375) <= 14546321;
srom_1(50376) <= 14921751;
srom_1(50377) <= 15266544;
srom_1(50378) <= 15579085;
srom_1(50379) <= 15857907;
srom_1(50380) <= 16101703;
srom_1(50381) <= 16309330;
srom_1(50382) <= 16479813;
srom_1(50383) <= 16612354;
srom_1(50384) <= 16706332;
srom_1(50385) <= 16761304;
srom_1(50386) <= 16777014;
srom_1(50387) <= 16753388;
srom_1(50388) <= 16690537;
srom_1(50389) <= 16588755;
srom_1(50390) <= 16448519;
srom_1(50391) <= 16270488;
srom_1(50392) <= 16055496;
srom_1(50393) <= 15804552;
srom_1(50394) <= 15518831;
srom_1(50395) <= 15199675;
srom_1(50396) <= 14848579;
srom_1(50397) <= 14467190;
srom_1(50398) <= 14057296;
srom_1(50399) <= 13620820;
srom_1(50400) <= 13159809;
srom_1(50401) <= 12676423;
srom_1(50402) <= 12172931;
srom_1(50403) <= 11651692;
srom_1(50404) <= 11115152;
srom_1(50405) <= 10565826;
srom_1(50406) <= 10006290;
srom_1(50407) <= 9439169;
srom_1(50408) <= 8867121;
srom_1(50409) <= 8292829;
srom_1(50410) <= 7718986;
srom_1(50411) <= 7148283;
srom_1(50412) <= 6583397;
srom_1(50413) <= 6026976;
srom_1(50414) <= 5481629;
srom_1(50415) <= 4949914;
srom_1(50416) <= 4434325;
srom_1(50417) <= 3937278;
srom_1(50418) <= 3461105;
srom_1(50419) <= 3008039;
srom_1(50420) <= 2580204;
srom_1(50421) <= 2179607;
srom_1(50422) <= 1808126;
srom_1(50423) <= 1467503;
srom_1(50424) <= 1159336;
srom_1(50425) <= 885069;
srom_1(50426) <= 645989;
srom_1(50427) <= 443216;
srom_1(50428) <= 277702;
srom_1(50429) <= 150223;
srom_1(50430) <= 61377;
srom_1(50431) <= 11580;
srom_1(50432) <= 1065;
srom_1(50433) <= 29883;
srom_1(50434) <= 97898;
srom_1(50435) <= 204790;
srom_1(50436) <= 350060;
srom_1(50437) <= 533024;
srom_1(50438) <= 752827;
srom_1(50439) <= 1008436;
srom_1(50440) <= 1298653;
srom_1(50441) <= 1622118;
srom_1(50442) <= 1977313;
srom_1(50443) <= 2362572;
srom_1(50444) <= 2776090;
srom_1(50445) <= 3215927;
srom_1(50446) <= 3680020;
srom_1(50447) <= 4166194;
srom_1(50448) <= 4672167;
srom_1(50449) <= 5195569;
srom_1(50450) <= 5733944;
srom_1(50451) <= 6284767;
srom_1(50452) <= 6845456;
srom_1(50453) <= 7413381;
srom_1(50454) <= 7985880;
srom_1(50455) <= 8560267;
srom_1(50456) <= 9133849;
srom_1(50457) <= 9703936;
srom_1(50458) <= 10267856;
srom_1(50459) <= 10822963;
srom_1(50460) <= 11366654;
srom_1(50461) <= 11896380;
srom_1(50462) <= 12409657;
srom_1(50463) <= 12904078;
srom_1(50464) <= 13377325;
srom_1(50465) <= 13827177;
srom_1(50466) <= 14251527;
srom_1(50467) <= 14648383;
srom_1(50468) <= 15015885;
srom_1(50469) <= 15352309;
srom_1(50470) <= 15656078;
srom_1(50471) <= 15925767;
srom_1(50472) <= 16160112;
srom_1(50473) <= 16358014;
srom_1(50474) <= 16518544;
srom_1(50475) <= 16640951;
srom_1(50476) <= 16724659;
srom_1(50477) <= 16769277;
srom_1(50478) <= 16774595;
srom_1(50479) <= 16740588;
srom_1(50480) <= 16667415;
srom_1(50481) <= 16555421;
srom_1(50482) <= 16405130;
srom_1(50483) <= 16217246;
srom_1(50484) <= 15992651;
srom_1(50485) <= 15732398;
srom_1(50486) <= 15437708;
srom_1(50487) <= 15109962;
srom_1(50488) <= 14750697;
srom_1(50489) <= 14361598;
srom_1(50490) <= 13944490;
srom_1(50491) <= 13501329;
srom_1(50492) <= 13034192;
srom_1(50493) <= 12545270;
srom_1(50494) <= 12036856;
srom_1(50495) <= 11511335;
srom_1(50496) <= 10971169;
srom_1(50497) <= 10418894;
srom_1(50498) <= 9857097;
srom_1(50499) <= 9288415;
srom_1(50500) <= 8715512;
srom_1(50501) <= 8141077;
srom_1(50502) <= 7567803;
srom_1(50503) <= 6998377;
srom_1(50504) <= 6435471;
srom_1(50505) <= 5881724;
srom_1(50506) <= 5339733;
srom_1(50507) <= 4812038;
srom_1(50508) <= 4301116;
srom_1(50509) <= 3809361;
srom_1(50510) <= 3339079;
srom_1(50511) <= 2892477;
srom_1(50512) <= 2471648;
srom_1(50513) <= 2078566;
srom_1(50514) <= 1715073;
srom_1(50515) <= 1382875;
srom_1(50516) <= 1083530;
srom_1(50517) <= 818440;
srom_1(50518) <= 588849;
srom_1(50519) <= 395834;
srom_1(50520) <= 240300;
srom_1(50521) <= 122977;
srom_1(50522) <= 44413;
srom_1(50523) <= 4979;
srom_1(50524) <= 4858;
srom_1(50525) <= 44051;
srom_1(50526) <= 122375;
srom_1(50527) <= 239462;
srom_1(50528) <= 394763;
srom_1(50529) <= 587550;
srom_1(50530) <= 816919;
srom_1(50531) <= 1081795;
srom_1(50532) <= 1380934;
srom_1(50533) <= 1712935;
srom_1(50534) <= 2076240;
srom_1(50535) <= 2469146;
srom_1(50536) <= 2889810;
srom_1(50537) <= 3336260;
srom_1(50538) <= 3806403;
srom_1(50539) <= 4298033;
srom_1(50540) <= 4808845;
srom_1(50541) <= 5336444;
srom_1(50542) <= 5878355;
srom_1(50543) <= 6432038;
srom_1(50544) <= 6994896;
srom_1(50545) <= 7564289;
srom_1(50546) <= 8137548;
srom_1(50547) <= 8711984;
srom_1(50548) <= 9284904;
srom_1(50549) <= 9853621;
srom_1(50550) <= 10415468;
srom_1(50551) <= 10967810;
srom_1(50552) <= 11508057;
srom_1(50553) <= 12033676;
srom_1(50554) <= 12542203;
srom_1(50555) <= 13031251;
srom_1(50556) <= 13498529;
srom_1(50557) <= 13941844;
srom_1(50558) <= 14359119;
srom_1(50559) <= 14748395;
srom_1(50560) <= 15107849;
srom_1(50561) <= 15435793;
srom_1(50562) <= 15730691;
srom_1(50563) <= 15991160;
srom_1(50564) <= 16215977;
srom_1(50565) <= 16404089;
srom_1(50566) <= 16554614;
srom_1(50567) <= 16666845;
srom_1(50568) <= 16740257;
srom_1(50569) <= 16774506;
srom_1(50570) <= 16769430;
srom_1(50571) <= 16725053;
srom_1(50572) <= 16641584;
srom_1(50573) <= 16519414;
srom_1(50574) <= 16359115;
srom_1(50575) <= 16161441;
srom_1(50576) <= 15927316;
srom_1(50577) <= 15657841;
srom_1(50578) <= 15354277;
srom_1(50579) <= 15018049;
srom_1(50580) <= 14650733;
srom_1(50581) <= 14254051;
srom_1(50582) <= 13829865;
srom_1(50583) <= 13380163;
srom_1(50584) <= 12907054;
srom_1(50585) <= 12412756;
srom_1(50586) <= 11899587;
srom_1(50587) <= 11369955;
srom_1(50588) <= 10826341;
srom_1(50589) <= 10271297;
srom_1(50590) <= 9707423;
srom_1(50591) <= 9137366;
srom_1(50592) <= 8563797;
srom_1(50593) <= 7989407;
srom_1(50594) <= 7416888;
srom_1(50595) <= 6848927;
srom_1(50596) <= 6288185;
srom_1(50597) <= 5737293;
srom_1(50598) <= 5198834;
srom_1(50599) <= 4675333;
srom_1(50600) <= 4169245;
srom_1(50601) <= 3682943;
srom_1(50602) <= 3218707;
srom_1(50603) <= 2778715;
srom_1(50604) <= 2365029;
srom_1(50605) <= 1979590;
srom_1(50606) <= 1624205;
srom_1(50607) <= 1300541;
srom_1(50608) <= 1010115;
srom_1(50609) <= 754289;
srom_1(50610) <= 534264;
srom_1(50611) <= 351070;
srom_1(50612) <= 205566;
srom_1(50613) <= 98436;
srom_1(50614) <= 30182;
srom_1(50615) <= 1122;
srom_1(50616) <= 11395;
srom_1(50617) <= 60951;
srom_1(50618) <= 149559;
srom_1(50619) <= 276802;
srom_1(50620) <= 442084;
srom_1(50621) <= 644631;
srom_1(50622) <= 883491;
srom_1(50623) <= 1157545;
srom_1(50624) <= 1465509;
srom_1(50625) <= 1805937;
srom_1(50626) <= 2177234;
srom_1(50627) <= 2577657;
srom_1(50628) <= 3005331;
srom_1(50629) <= 3458248;
srom_1(50630) <= 3934286;
srom_1(50631) <= 4431211;
srom_1(50632) <= 4946694;
srom_1(50633) <= 5478317;
srom_1(50634) <= 6023588;
srom_1(50635) <= 6579949;
srom_1(50636) <= 7144791;
srom_1(50637) <= 7715467;
srom_1(50638) <= 8289298;
srom_1(50639) <= 8863596;
srom_1(50640) <= 9435666;
srom_1(50641) <= 10002826;
srom_1(50642) <= 10562416;
srom_1(50643) <= 11111813;
srom_1(50644) <= 11648439;
srom_1(50645) <= 12169779;
srom_1(50646) <= 12673388;
srom_1(50647) <= 13156904;
srom_1(50648) <= 13618060;
srom_1(50649) <= 14054693;
srom_1(50650) <= 14464756;
srom_1(50651) <= 14846326;
srom_1(50652) <= 15197613;
srom_1(50653) <= 15516971;
srom_1(50654) <= 15802901;
srom_1(50655) <= 16054063;
srom_1(50656) <= 16269279;
srom_1(50657) <= 16447540;
srom_1(50658) <= 16588010;
srom_1(50659) <= 16690030;
srom_1(50660) <= 16753121;
srom_1(50661) <= 16776989;
srom_1(50662) <= 16761521;
srom_1(50663) <= 16706789;
srom_1(50664) <= 16613050;
srom_1(50665) <= 16480744;
srom_1(50666) <= 16310492;
srom_1(50667) <= 16103090;
srom_1(50668) <= 15859513;
srom_1(50669) <= 15580903;
srom_1(50670) <= 15268565;
srom_1(50671) <= 14923965;
srom_1(50672) <= 14548718;
srom_1(50673) <= 14144584;
srom_1(50674) <= 13713459;
srom_1(50675) <= 13257363;
srom_1(50676) <= 12778436;
srom_1(50677) <= 12278924;
srom_1(50678) <= 11761169;
srom_1(50679) <= 11227599;
srom_1(50680) <= 10680715;
srom_1(50681) <= 10123083;
srom_1(50682) <= 9557318;
srom_1(50683) <= 8986072;
srom_1(50684) <= 8412024;
srom_1(50685) <= 7837867;
srom_1(50686) <= 7266292;
srom_1(50687) <= 6699980;
srom_1(50688) <= 6141587;
srom_1(50689) <= 5593730;
srom_1(50690) <= 5058980;
srom_1(50691) <= 4539844;
srom_1(50692) <= 4038756;
srom_1(50693) <= 3558065;
srom_1(50694) <= 3100027;
srom_1(50695) <= 2666789;
srom_1(50696) <= 2260382;
srom_1(50697) <= 1882713;
srom_1(50698) <= 1535552;
srom_1(50699) <= 1220527;
srom_1(50700) <= 939116;
srom_1(50701) <= 692638;
srom_1(50702) <= 482249;
srom_1(50703) <= 308936;
srom_1(50704) <= 173511;
srom_1(50705) <= 76610;
srom_1(50706) <= 18686;
srom_1(50707) <= 12;
srom_1(50708) <= 20675;
srom_1(50709) <= 80578;
srom_1(50710) <= 179440;
srom_1(50711) <= 316798;
srom_1(50712) <= 492007;
srom_1(50713) <= 704246;
srom_1(50714) <= 952520;
srom_1(50715) <= 1235664;
srom_1(50716) <= 1552350;
srom_1(50717) <= 1901095;
srom_1(50718) <= 2280261;
srom_1(50719) <= 2688071;
srom_1(50720) <= 3122614;
srom_1(50721) <= 3581850;
srom_1(50722) <= 4063627;
srom_1(50723) <= 4565685;
srom_1(50724) <= 5085670;
srom_1(50725) <= 5621144;
srom_1(50726) <= 6169595;
srom_1(50727) <= 6728452;
srom_1(50728) <= 7295095;
srom_1(50729) <= 7866864;
srom_1(50730) <= 8441081;
srom_1(50731) <= 9015052;
srom_1(50732) <= 9586084;
srom_1(50733) <= 10151502;
srom_1(50734) <= 10708653;
srom_1(50735) <= 11254924;
srom_1(50736) <= 11787754;
srom_1(50737) <= 12304644;
srom_1(50738) <= 12803171;
srom_1(50739) <= 13280996;
srom_1(50740) <= 13735879;
srom_1(50741) <= 14165687;
srom_1(50742) <= 14568404;
srom_1(50743) <= 14942142;
srom_1(50744) <= 15285148;
srom_1(50745) <= 15595814;
srom_1(50746) <= 15872683;
srom_1(50747) <= 16114457;
srom_1(50748) <= 16320001;
srom_1(50749) <= 16488352;
srom_1(50750) <= 16618721;
srom_1(50751) <= 16710496;
srom_1(50752) <= 16763247;
srom_1(50753) <= 16776726;
srom_1(50754) <= 16750871;
srom_1(50755) <= 16685802;
srom_1(50756) <= 16581824;
srom_1(50757) <= 16439426;
srom_1(50758) <= 16259274;
srom_1(50759) <= 16042215;
srom_1(50760) <= 15789265;
srom_1(50761) <= 15501610;
srom_1(50762) <= 15180601;
srom_1(50763) <= 14827741;
srom_1(50764) <= 14444686;
srom_1(50765) <= 14033232;
srom_1(50766) <= 13595309;
srom_1(50767) <= 13132969;
srom_1(50768) <= 12648382;
srom_1(50769) <= 12143819;
srom_1(50770) <= 11621646;
srom_1(50771) <= 11084313;
srom_1(50772) <= 10534339;
srom_1(50773) <= 9974302;
srom_1(50774) <= 9406830;
srom_1(50775) <= 8834582;
srom_1(50776) <= 8260244;
srom_1(50777) <= 7686507;
srom_1(50778) <= 7116063;
srom_1(50779) <= 6551586;
srom_1(50780) <= 5995724;
srom_1(50781) <= 5451083;
srom_1(50782) <= 4920216;
srom_1(50783) <= 4405615;
srom_1(50784) <= 3909690;
srom_1(50785) <= 3434769;
srom_1(50786) <= 2983079;
srom_1(50787) <= 2556736;
srom_1(50788) <= 2157741;
srom_1(50789) <= 1787965;
srom_1(50790) <= 1449142;
srom_1(50791) <= 1142860;
srom_1(50792) <= 870556;
srom_1(50793) <= 633507;
srom_1(50794) <= 432824;
srom_1(50795) <= 269448;
srom_1(50796) <= 144146;
srom_1(50797) <= 57505;
srom_1(50798) <= 9931;
srom_1(50799) <= 1648;
srom_1(50800) <= 32694;
srom_1(50801) <= 102924;
srom_1(50802) <= 212009;
srom_1(50803) <= 359436;
srom_1(50804) <= 544515;
srom_1(50805) <= 766377;
srom_1(50806) <= 1023983;
srom_1(50807) <= 1316124;
srom_1(50808) <= 1641430;
srom_1(50809) <= 1998376;
srom_1(50810) <= 2385288;
srom_1(50811) <= 2800352;
srom_1(50812) <= 3241621;
srom_1(50813) <= 3707026;
srom_1(50814) <= 4194384;
srom_1(50815) <= 4701411;
srom_1(50816) <= 5225728;
srom_1(50817) <= 5764877;
srom_1(50818) <= 6316329;
srom_1(50819) <= 6877499;
srom_1(50820) <= 7445756;
srom_1(50821) <= 8018433;
srom_1(50822) <= 8592847;
srom_1(50823) <= 9166302;
srom_1(50824) <= 9736111;
srom_1(50825) <= 10299601;
srom_1(50826) <= 10854130;
srom_1(50827) <= 11397097;
srom_1(50828) <= 11925956;
srom_1(50829) <= 12438227;
srom_1(50830) <= 12931508;
srom_1(50831) <= 13403486;
srom_1(50832) <= 13851947;
srom_1(50833) <= 14274789;
srom_1(50834) <= 14670029;
srom_1(50835) <= 15035813;
srom_1(50836) <= 15370426;
srom_1(50837) <= 15672298;
srom_1(50838) <= 15940015;
srom_1(50839) <= 16172321;
srom_1(50840) <= 16368127;
srom_1(50841) <= 16526513;
srom_1(50842) <= 16646738;
srom_1(50843) <= 16728238;
srom_1(50844) <= 16770631;
srom_1(50845) <= 16773717;
srom_1(50846) <= 16737483;
srom_1(50847) <= 16662098;
srom_1(50848) <= 16547915;
srom_1(50849) <= 16395471;
srom_1(50850) <= 16205480;
srom_1(50851) <= 15978833;
srom_1(50852) <= 15716593;
srom_1(50853) <= 15419989;
srom_1(50854) <= 15090413;
srom_1(50855) <= 14729410;
srom_1(50856) <= 14338672;
srom_1(50857) <= 13920033;
srom_1(50858) <= 13475454;
srom_1(50859) <= 13007022;
srom_1(50860) <= 12516933;
srom_1(50861) <= 12007484;
srom_1(50862) <= 11481065;
srom_1(50863) <= 10940145;
srom_1(50864) <= 10387259;
srom_1(50865) <= 9825002;
srom_1(50866) <= 9256008;
srom_1(50867) <= 8682947;
srom_1(50868) <= 8108506;
srom_1(50869) <= 7535378;
srom_1(50870) <= 6966251;
srom_1(50871) <= 6403794;
srom_1(50872) <= 5850645;
srom_1(50873) <= 5309396;
srom_1(50874) <= 4782588;
srom_1(50875) <= 4272689;
srom_1(50876) <= 3782091;
srom_1(50877) <= 3313095;
srom_1(50878) <= 2867900;
srom_1(50879) <= 2448593;
srom_1(50880) <= 2057141;
srom_1(50881) <= 1695379;
srom_1(50882) <= 1365004;
srom_1(50883) <= 1067565;
srom_1(50884) <= 804457;
srom_1(50885) <= 576914;
srom_1(50886) <= 386002;
srom_1(50887) <= 232618;
srom_1(50888) <= 117480;
srom_1(50889) <= 41127;
srom_1(50890) <= 3919;
srom_1(50891) <= 6030;
srom_1(50892) <= 47449;
srom_1(50893) <= 127983;
srom_1(50894) <= 247254;
srom_1(50895) <= 404703;
srom_1(50896) <= 599591;
srom_1(50897) <= 831004;
srom_1(50898) <= 1097857;
srom_1(50899) <= 1398899;
srom_1(50900) <= 1732719;
srom_1(50901) <= 2097750;
srom_1(50902) <= 2492281;
srom_1(50903) <= 2914462;
srom_1(50904) <= 3362313;
srom_1(50905) <= 3833734;
srom_1(50906) <= 4326514;
srom_1(50907) <= 4838343;
srom_1(50908) <= 5366821;
srom_1(50909) <= 5909468;
srom_1(50910) <= 6463741;
srom_1(50911) <= 7027041;
srom_1(50912) <= 7596725;
srom_1(50913) <= 8170123;
srom_1(50914) <= 8744545;
srom_1(50915) <= 9317298;
srom_1(50916) <= 9885697;
srom_1(50917) <= 10447075;
srom_1(50918) <= 10998800;
srom_1(50919) <= 11538284;
srom_1(50920) <= 12062999;
srom_1(50921) <= 12570484;
srom_1(50922) <= 13058358;
srom_1(50923) <= 13524334;
srom_1(50924) <= 13966227;
srom_1(50925) <= 14381965;
srom_1(50926) <= 14769597;
srom_1(50927) <= 15127307;
srom_1(50928) <= 15453417;
srom_1(50929) <= 15746398;
srom_1(50930) <= 16004875;
srom_1(50931) <= 16227637;
srom_1(50932) <= 16413640;
srom_1(50933) <= 16562010;
srom_1(50934) <= 16672052;
srom_1(50935) <= 16743250;
srom_1(50936) <= 16775270;
srom_1(50937) <= 16767963;
srom_1(50938) <= 16721362;
srom_1(50939) <= 16635685;
srom_1(50940) <= 16511335;
srom_1(50941) <= 16348895;
srom_1(50942) <= 16149127;
srom_1(50943) <= 15912967;
srom_1(50944) <= 15641522;
srom_1(50945) <= 15336066;
srom_1(50946) <= 14998031;
srom_1(50947) <= 14629002;
srom_1(50948) <= 14230710;
srom_1(50949) <= 13805022;
srom_1(50950) <= 13353935;
srom_1(50951) <= 12879563;
srom_1(50952) <= 12384132;
srom_1(50953) <= 11869965;
srom_1(50954) <= 11339472;
srom_1(50955) <= 10795141;
srom_1(50956) <= 10239526;
srom_1(50957) <= 9675231;
srom_1(50958) <= 9104903;
srom_1(50959) <= 8531215;
srom_1(50960) <= 7956859;
srom_1(50961) <= 7384527;
srom_1(50962) <= 6816904;
srom_1(50963) <= 6256651;
srom_1(50964) <= 5706396;
srom_1(50965) <= 5168718;
srom_1(50966) <= 4646140;
srom_1(50967) <= 4141111;
srom_1(50968) <= 3656001;
srom_1(50969) <= 3193083;
srom_1(50970) <= 2754528;
srom_1(50971) <= 2342394;
srom_1(50972) <= 1958613;
srom_1(50973) <= 1604984;
srom_1(50974) <= 1283166;
srom_1(50975) <= 994667;
srom_1(50976) <= 740842;
srom_1(50977) <= 522879;
srom_1(50978) <= 341801;
srom_1(50979) <= 198458;
srom_1(50980) <= 93521;
srom_1(50981) <= 27483;
srom_1(50982) <= 652;
srom_1(50983) <= 13156;
srom_1(50984) <= 64935;
srom_1(50985) <= 155747;
srom_1(50986) <= 285166;
srom_1(50987) <= 452584;
srom_1(50988) <= 657217;
srom_1(50989) <= 898105;
srom_1(50990) <= 1174118;
srom_1(50991) <= 1483963;
srom_1(50992) <= 1826186;
srom_1(50993) <= 2199183;
srom_1(50994) <= 2601204;
srom_1(50995) <= 3030364;
srom_1(50996) <= 3484650;
srom_1(50997) <= 3961933;
srom_1(50998) <= 4459974;
srom_1(50999) <= 4976438;
srom_1(51000) <= 5508903;
srom_1(51001) <= 6054872;
srom_1(51002) <= 6611784;
srom_1(51003) <= 7177028;
srom_1(51004) <= 7747954;
srom_1(51005) <= 8321884;
srom_1(51006) <= 8896128;
srom_1(51007) <= 9467991;
srom_1(51008) <= 10034792;
srom_1(51009) <= 10593874;
srom_1(51010) <= 11142615;
srom_1(51011) <= 11678441;
srom_1(51012) <= 12198840;
srom_1(51013) <= 12701372;
srom_1(51014) <= 13183679;
srom_1(51015) <= 13643501;
srom_1(51016) <= 14078681;
srom_1(51017) <= 14487178;
srom_1(51018) <= 14867077;
srom_1(51019) <= 15216596;
srom_1(51020) <= 15534096;
srom_1(51021) <= 15818088;
srom_1(51022) <= 16067242;
srom_1(51023) <= 16280387;
srom_1(51024) <= 16456525;
srom_1(51025) <= 16594830;
srom_1(51026) <= 16694653;
srom_1(51027) <= 16755526;
srom_1(51028) <= 16777164;
srom_1(51029) <= 16759465;
srom_1(51030) <= 16702512;
srom_1(51031) <= 16606573;
srom_1(51032) <= 16472096;
srom_1(51033) <= 16299714;
srom_1(51034) <= 16090233;
srom_1(51035) <= 15844637;
srom_1(51036) <= 15564077;
srom_1(51037) <= 15249868;
srom_1(51038) <= 14903485;
srom_1(51039) <= 14526552;
srom_1(51040) <= 14120835;
srom_1(51041) <= 13688238;
srom_1(51042) <= 13230789;
srom_1(51043) <= 12750634;
srom_1(51044) <= 12250023;
srom_1(51045) <= 11731305;
srom_1(51046) <= 11196912;
srom_1(51047) <= 10649350;
srom_1(51048) <= 10091187;
srom_1(51049) <= 9525039;
srom_1(51050) <= 8953562;
srom_1(51051) <= 8379437;
srom_1(51052) <= 7805354;
srom_1(51053) <= 7234006;
srom_1(51054) <= 6668072;
srom_1(51055) <= 6110207;
srom_1(51056) <= 5563026;
srom_1(51057) <= 5029095;
srom_1(51058) <= 4510918;
srom_1(51059) <= 4010924;
srom_1(51060) <= 3531459;
srom_1(51061) <= 3074771;
srom_1(51062) <= 2643002;
srom_1(51063) <= 2238175;
srom_1(51064) <= 1862190;
srom_1(51065) <= 1516810;
srom_1(51066) <= 1203653;
srom_1(51067) <= 924190;
srom_1(51068) <= 679730;
srom_1(51069) <= 471419;
srom_1(51070) <= 300235;
srom_1(51071) <= 166980;
srom_1(51072) <= 72278;
srom_1(51073) <= 16575;
srom_1(51074) <= 132;
srom_1(51075) <= 23025;
srom_1(51076) <= 85146;
srom_1(51077) <= 186206;
srom_1(51078) <= 325730;
srom_1(51079) <= 503063;
srom_1(51080) <= 717374;
srom_1(51081) <= 967658;
srom_1(51082) <= 1252742;
srom_1(51083) <= 1571288;
srom_1(51084) <= 1921803;
srom_1(51085) <= 2302642;
srom_1(51086) <= 2712022;
srom_1(51087) <= 3148020;
srom_1(51088) <= 3608594;
srom_1(51089) <= 4091582;
srom_1(51090) <= 4594721;
srom_1(51091) <= 5115651;
srom_1(51092) <= 5651928;
srom_1(51093) <= 6201039;
srom_1(51094) <= 6760408;
srom_1(51095) <= 7327412;
srom_1(51096) <= 7899393;
srom_1(51097) <= 8473668;
srom_1(51098) <= 9047544;
srom_1(51099) <= 9618329;
srom_1(51100) <= 10183349;
srom_1(51101) <= 10739952;
srom_1(51102) <= 11285529;
srom_1(51103) <= 11817521;
srom_1(51104) <= 12333433;
srom_1(51105) <= 12830848;
srom_1(51106) <= 13307431;
srom_1(51107) <= 13760947;
srom_1(51108) <= 14189272;
srom_1(51109) <= 14590394;
srom_1(51110) <= 14962435;
srom_1(51111) <= 15303648;
srom_1(51112) <= 15612435;
srom_1(51113) <= 15887347;
srom_1(51114) <= 16127094;
srom_1(51115) <= 16330553;
srom_1(51116) <= 16496769;
srom_1(51117) <= 16624964;
srom_1(51118) <= 16714535;
srom_1(51119) <= 16765063;
srom_1(51120) <= 16776312;
srom_1(51121) <= 16748227;
srom_1(51122) <= 16680941;
srom_1(51123) <= 16574770;
srom_1(51124) <= 16430211;
srom_1(51125) <= 16247942;
srom_1(51126) <= 16028817;
srom_1(51127) <= 15773866;
srom_1(51128) <= 15484282;
srom_1(51129) <= 15161424;
srom_1(51130) <= 14806806;
srom_1(51131) <= 14422091;
srom_1(51132) <= 14009083;
srom_1(51133) <= 13569719;
srom_1(51134) <= 13106058;
srom_1(51135) <= 12620276;
srom_1(51136) <= 12114650;
srom_1(51137) <= 11591552;
srom_1(51138) <= 11053433;
srom_1(51139) <= 10502819;
srom_1(51140) <= 9942290;
srom_1(51141) <= 9374475;
srom_1(51142) <= 8802037;
srom_1(51143) <= 8227661;
srom_1(51144) <= 7654039;
srom_1(51145) <= 7083862;
srom_1(51146) <= 6519803;
srom_1(51147) <= 5964508;
srom_1(51148) <= 5420580;
srom_1(51149) <= 4890571;
srom_1(51150) <= 4376964;
srom_1(51151) <= 3882170;
srom_1(51152) <= 3408508;
srom_1(51153) <= 2958200;
srom_1(51154) <= 2533356;
srom_1(51155) <= 2135970;
srom_1(51156) <= 1767904;
srom_1(51157) <= 1430885;
srom_1(51158) <= 1126494;
srom_1(51159) <= 856157;
srom_1(51160) <= 621142;
srom_1(51161) <= 422551;
srom_1(51162) <= 261316;
srom_1(51163) <= 138193;
srom_1(51164) <= 53759;
srom_1(51165) <= 8409;
srom_1(51166) <= 2357;
srom_1(51167) <= 35632;
srom_1(51168) <= 108076;
srom_1(51169) <= 219351;
srom_1(51170) <= 368933;
srom_1(51171) <= 556123;
srom_1(51172) <= 780043;
srom_1(51173) <= 1039641;
srom_1(51174) <= 1333701;
srom_1(51175) <= 1660844;
srom_1(51176) <= 2019536;
srom_1(51177) <= 2408095;
srom_1(51178) <= 2824698;
srom_1(51179) <= 3267392;
srom_1(51180) <= 3734102;
srom_1(51181) <= 4222638;
srom_1(51182) <= 4730709;
srom_1(51183) <= 5255934;
srom_1(51184) <= 5795849;
srom_1(51185) <= 6347923;
srom_1(51186) <= 6909565;
srom_1(51187) <= 7478144;
srom_1(51188) <= 8050992;
srom_1(51189) <= 8625423;
srom_1(51190) <= 9198744;
srom_1(51191) <= 9768266;
srom_1(51192) <= 10331318;
srom_1(51193) <= 10885259;
srom_1(51194) <= 11427494;
srom_1(51195) <= 11955478;
srom_1(51196) <= 12466735;
srom_1(51197) <= 12958869;
srom_1(51198) <= 13429571;
srom_1(51199) <= 13876635;
srom_1(51200) <= 14297963;
srom_1(51201) <= 14691581;
srom_1(51202) <= 15055641;
srom_1(51203) <= 15388437;
srom_1(51204) <= 15688409;
srom_1(51205) <= 15954150;
srom_1(51206) <= 16184413;
srom_1(51207) <= 16378119;
srom_1(51208) <= 16534359;
srom_1(51209) <= 16652401;
srom_1(51210) <= 16731692;
srom_1(51211) <= 16771858;
srom_1(51212) <= 16772713;
srom_1(51213) <= 16734252;
srom_1(51214) <= 16656655;
srom_1(51215) <= 16540287;
srom_1(51216) <= 16385692;
srom_1(51217) <= 16193596;
srom_1(51218) <= 15964901;
srom_1(51219) <= 15700677;
srom_1(51220) <= 15402164;
srom_1(51221) <= 15070763;
srom_1(51222) <= 14708026;
srom_1(51223) <= 14315656;
srom_1(51224) <= 13895492;
srom_1(51225) <= 13449504;
srom_1(51226) <= 12979783;
srom_1(51227) <= 12488533;
srom_1(51228) <= 11978058;
srom_1(51229) <= 11450749;
srom_1(51230) <= 10909082;
srom_1(51231) <= 10355595;
srom_1(51232) <= 9792884;
srom_1(51233) <= 9223588;
srom_1(51234) <= 8650377;
srom_1(51235) <= 8075938;
srom_1(51236) <= 7502965;
srom_1(51237) <= 6934146;
srom_1(51238) <= 6372147;
srom_1(51239) <= 5819603;
srom_1(51240) <= 5279107;
srom_1(51241) <= 4753192;
srom_1(51242) <= 4244325;
srom_1(51243) <= 3754892;
srom_1(51244) <= 3287187;
srom_1(51245) <= 2843406;
srom_1(51246) <= 2425627;
srom_1(51247) <= 2035811;
srom_1(51248) <= 1675786;
srom_1(51249) <= 1347239;
srom_1(51250) <= 1051711;
srom_1(51251) <= 790589;
srom_1(51252) <= 565097;
srom_1(51253) <= 376291;
srom_1(51254) <= 225058;
srom_1(51255) <= 112107;
srom_1(51256) <= 37967;
srom_1(51257) <= 2986;
srom_1(51258) <= 7329;
srom_1(51259) <= 50974;
srom_1(51260) <= 133717;
srom_1(51261) <= 255169;
srom_1(51262) <= 414763;
srom_1(51263) <= 611748;
srom_1(51264) <= 845202;
srom_1(51265) <= 1114030;
srom_1(51266) <= 1416970;
srom_1(51267) <= 1752603;
srom_1(51268) <= 2119355;
srom_1(51269) <= 2515505;
srom_1(51270) <= 2939196;
srom_1(51271) <= 3388441;
srom_1(51272) <= 3861134;
srom_1(51273) <= 4355057;
srom_1(51274) <= 4867895;
srom_1(51275) <= 5397244;
srom_1(51276) <= 5940619;
srom_1(51277) <= 6495474;
srom_1(51278) <= 7059207;
srom_1(51279) <= 7629174;
srom_1(51280) <= 8202701;
srom_1(51281) <= 8777101;
srom_1(51282) <= 9349679;
srom_1(51283) <= 9917750;
srom_1(51284) <= 10478650;
srom_1(51285) <= 11029750;
srom_1(51286) <= 11568464;
srom_1(51287) <= 12092267;
srom_1(51288) <= 12598702;
srom_1(51289) <= 13085394;
srom_1(51290) <= 13550062;
srom_1(51291) <= 13990526;
srom_1(51292) <= 14404720;
srom_1(51293) <= 14790703;
srom_1(51294) <= 15146664;
srom_1(51295) <= 15470935;
srom_1(51296) <= 15761993;
srom_1(51297) <= 16018476;
srom_1(51298) <= 16239179;
srom_1(51299) <= 16423069;
srom_1(51300) <= 16569282;
srom_1(51301) <= 16677133;
srom_1(51302) <= 16746116;
srom_1(51303) <= 16775908;
srom_1(51304) <= 16766370;
srom_1(51305) <= 16717544;
srom_1(51306) <= 16629662;
srom_1(51307) <= 16503135;
srom_1(51308) <= 16338555;
srom_1(51309) <= 16136696;
srom_1(51310) <= 15898503;
srom_1(51311) <= 15625094;
srom_1(51312) <= 15317750;
srom_1(51313) <= 14977914;
srom_1(51314) <= 14607177;
srom_1(51315) <= 14207280;
srom_1(51316) <= 13780097;
srom_1(51317) <= 13327631;
srom_1(51318) <= 12852005;
srom_1(51319) <= 12355448;
srom_1(51320) <= 11840289;
srom_1(51321) <= 11308945;
srom_1(51322) <= 10763905;
srom_1(51323) <= 10207727;
srom_1(51324) <= 9643019;
srom_1(51325) <= 9072428;
srom_1(51326) <= 8498631;
srom_1(51327) <= 7924318;
srom_1(51328) <= 7352181;
srom_1(51329) <= 6784905;
srom_1(51330) <= 6225150;
srom_1(51331) <= 5675539;
srom_1(51332) <= 5138651;
srom_1(51333) <= 4617003;
srom_1(51334) <= 4113042;
srom_1(51335) <= 3629130;
srom_1(51336) <= 3167537;
srom_1(51337) <= 2730427;
srom_1(51338) <= 2319851;
srom_1(51339) <= 1937733;
srom_1(51340) <= 1585865;
srom_1(51341) <= 1265898;
srom_1(51342) <= 979331;
srom_1(51343) <= 727509;
srom_1(51344) <= 511613;
srom_1(51345) <= 332655;
srom_1(51346) <= 191473;
srom_1(51347) <= 88731;
srom_1(51348) <= 24910;
srom_1(51349) <= 309;
srom_1(51350) <= 15044;
srom_1(51351) <= 69045;
srom_1(51352) <= 162060;
srom_1(51353) <= 293651;
srom_1(51354) <= 463203;
srom_1(51355) <= 669920;
srom_1(51356) <= 912832;
srom_1(51357) <= 1190800;
srom_1(51358) <= 1502522;
srom_1(51359) <= 1846535;
srom_1(51360) <= 2221226;
srom_1(51361) <= 2624837;
srom_1(51362) <= 3055478;
srom_1(51363) <= 3511127;
srom_1(51364) <= 3989648;
srom_1(51365) <= 4488797;
srom_1(51366) <= 5006234;
srom_1(51367) <= 5539532;
srom_1(51368) <= 6086191;
srom_1(51369) <= 6643646;
srom_1(51370) <= 7209284;
srom_1(51371) <= 7780452;
srom_1(51372) <= 8354472;
srom_1(51373) <= 8928652;
srom_1(51374) <= 9500299;
srom_1(51375) <= 10066734;
srom_1(51376) <= 10625299;
srom_1(51377) <= 11173376;
srom_1(51378) <= 11708393;
srom_1(51379) <= 12227844;
srom_1(51380) <= 12729290;
srom_1(51381) <= 13210382;
srom_1(51382) <= 13668863;
srom_1(51383) <= 14102583;
srom_1(51384) <= 14509508;
srom_1(51385) <= 14887730;
srom_1(51386) <= 15235475;
srom_1(51387) <= 15551113;
srom_1(51388) <= 15833164;
srom_1(51389) <= 16080304;
srom_1(51390) <= 16291376;
srom_1(51391) <= 16465389;
srom_1(51392) <= 16601527;
srom_1(51393) <= 16699151;
srom_1(51394) <= 16757805;
srom_1(51395) <= 16777213;
srom_1(51396) <= 16757283;
srom_1(51397) <= 16698110;
srom_1(51398) <= 16599971;
srom_1(51399) <= 16463326;
srom_1(51400) <= 16288816;
srom_1(51401) <= 16077259;
srom_1(51402) <= 15829647;
srom_1(51403) <= 15547142;
srom_1(51404) <= 15231068;
srom_1(51405) <= 14882907;
srom_1(51406) <= 14504293;
srom_1(51407) <= 14096999;
srom_1(51408) <= 13662937;
srom_1(51409) <= 13204142;
srom_1(51410) <= 12722765;
srom_1(51411) <= 12221064;
srom_1(51412) <= 11701391;
srom_1(51413) <= 11166184;
srom_1(51414) <= 10617951;
srom_1(51415) <= 10059264;
srom_1(51416) <= 9492743;
srom_1(51417) <= 8921044;
srom_1(51418) <= 8346849;
srom_1(51419) <= 7772849;
srom_1(51420) <= 7201737;
srom_1(51421) <= 6636190;
srom_1(51422) <= 6078861;
srom_1(51423) <= 5532364;
srom_1(51424) <= 4999260;
srom_1(51425) <= 4482050;
srom_1(51426) <= 3983159;
srom_1(51427) <= 3504927;
srom_1(51428) <= 3049596;
srom_1(51429) <= 2619301;
srom_1(51430) <= 2216061;
srom_1(51431) <= 1841766;
srom_1(51432) <= 1498171;
srom_1(51433) <= 1186888;
srom_1(51434) <= 909377;
srom_1(51435) <= 666938;
srom_1(51436) <= 460708;
srom_1(51437) <= 291655;
srom_1(51438) <= 160572;
srom_1(51439) <= 68073;
srom_1(51440) <= 14591;
srom_1(51441) <= 378;
srom_1(51442) <= 25501;
srom_1(51443) <= 89840;
srom_1(51444) <= 193096;
srom_1(51445) <= 334783;
srom_1(51446) <= 514238;
srom_1(51447) <= 730618;
srom_1(51448) <= 982909;
srom_1(51449) <= 1269927;
srom_1(51450) <= 1590328;
srom_1(51451) <= 1942608;
srom_1(51452) <= 2325116;
srom_1(51453) <= 2736057;
srom_1(51454) <= 3173506;
srom_1(51455) <= 3635409;
srom_1(51456) <= 4119602;
srom_1(51457) <= 4623814;
srom_1(51458) <= 5145680;
srom_1(51459) <= 5682754;
srom_1(51460) <= 6232516;
srom_1(51461) <= 6792388;
srom_1(51462) <= 7359746;
srom_1(51463) <= 7931929;
srom_1(51464) <= 8506253;
srom_1(51465) <= 9080026;
srom_1(51466) <= 9650556;
srom_1(51467) <= 10215168;
srom_1(51468) <= 10771215;
srom_1(51469) <= 11316090;
srom_1(51470) <= 11847236;
srom_1(51471) <= 12362163;
srom_1(51472) <= 12858457;
srom_1(51473) <= 13333791;
srom_1(51474) <= 13785935;
srom_1(51475) <= 14212769;
srom_1(51476) <= 14612291;
srom_1(51477) <= 14982628;
srom_1(51478) <= 15322044;
srom_1(51479) <= 15628947;
srom_1(51480) <= 15901897;
srom_1(51481) <= 16139614;
srom_1(51482) <= 16340985;
srom_1(51483) <= 16505064;
srom_1(51484) <= 16631082;
srom_1(51485) <= 16718449;
srom_1(51486) <= 16766754;
srom_1(51487) <= 16775770;
srom_1(51488) <= 16745457;
srom_1(51489) <= 16675956;
srom_1(51490) <= 16567592;
srom_1(51491) <= 16420874;
srom_1(51492) <= 16236490;
srom_1(51493) <= 16015305;
srom_1(51494) <= 15758355;
srom_1(51495) <= 15466847;
srom_1(51496) <= 15142145;
srom_1(51497) <= 14785775;
srom_1(51498) <= 14399405;
srom_1(51499) <= 13984849;
srom_1(51500) <= 13544051;
srom_1(51501) <= 13079076;
srom_1(51502) <= 12592107;
srom_1(51503) <= 12085426;
srom_1(51504) <= 11561409;
srom_1(51505) <= 11022514;
srom_1(51506) <= 10471267;
srom_1(51507) <= 9910254;
srom_1(51508) <= 9342106;
srom_1(51509) <= 8769486;
srom_1(51510) <= 8195080;
srom_1(51511) <= 7621582;
srom_1(51512) <= 7051681;
srom_1(51513) <= 6488049;
srom_1(51514) <= 5933329;
srom_1(51515) <= 5390123;
srom_1(51516) <= 4860978;
srom_1(51517) <= 4348375;
srom_1(51518) <= 3854718;
srom_1(51519) <= 3382322;
srom_1(51520) <= 2933403;
srom_1(51521) <= 2510064;
srom_1(51522) <= 2114292;
srom_1(51523) <= 1747943;
srom_1(51524) <= 1412734;
srom_1(51525) <= 1110237;
srom_1(51526) <= 841871;
srom_1(51527) <= 608894;
srom_1(51528) <= 412399;
srom_1(51529) <= 253307;
srom_1(51530) <= 132364;
srom_1(51531) <= 50138;
srom_1(51532) <= 7014;
srom_1(51533) <= 3193;
srom_1(51534) <= 38695;
srom_1(51535) <= 113353;
srom_1(51536) <= 226816;
srom_1(51537) <= 378552;
srom_1(51538) <= 567850;
srom_1(51539) <= 793823;
srom_1(51540) <= 1055410;
srom_1(51541) <= 1351385;
srom_1(51542) <= 1680360;
srom_1(51543) <= 2040792;
srom_1(51544) <= 2430991;
srom_1(51545) <= 2849128;
srom_1(51546) <= 3293241;
srom_1(51547) <= 3761248;
srom_1(51548) <= 4250954;
srom_1(51549) <= 4760063;
srom_1(51550) <= 5286188;
srom_1(51551) <= 5826861;
srom_1(51552) <= 6379547;
srom_1(51553) <= 6941654;
srom_1(51554) <= 7510546;
srom_1(51555) <= 8083556;
srom_1(51556) <= 8657996;
srom_1(51557) <= 9231173;
srom_1(51558) <= 9800399;
srom_1(51559) <= 10363005;
srom_1(51560) <= 10916352;
srom_1(51561) <= 11457845;
srom_1(51562) <= 11984946;
srom_1(51563) <= 12495182;
srom_1(51564) <= 12986161;
srom_1(51565) <= 13455581;
srom_1(51566) <= 13901240;
srom_1(51567) <= 14321048;
srom_1(51568) <= 14713037;
srom_1(51569) <= 15075368;
srom_1(51570) <= 15406343;
srom_1(51571) <= 15704410;
srom_1(51572) <= 15968170;
srom_1(51573) <= 16196387;
srom_1(51574) <= 16387990;
srom_1(51575) <= 16542082;
srom_1(51576) <= 16657939;
srom_1(51577) <= 16735019;
srom_1(51578) <= 16772959;
srom_1(51579) <= 16771582;
srom_1(51580) <= 16730895;
srom_1(51581) <= 16651088;
srom_1(51582) <= 16532535;
srom_1(51583) <= 16375792;
srom_1(51584) <= 16181595;
srom_1(51585) <= 15950854;
srom_1(51586) <= 15684650;
srom_1(51587) <= 15384234;
srom_1(51588) <= 15051012;
srom_1(51589) <= 14686548;
srom_1(51590) <= 14292550;
srom_1(51591) <= 13870868;
srom_1(51592) <= 13423476;
srom_1(51593) <= 12952475;
srom_1(51594) <= 12460072;
srom_1(51595) <= 11948577;
srom_1(51596) <= 11420387;
srom_1(51597) <= 10877981;
srom_1(51598) <= 10323901;
srom_1(51599) <= 9760746;
srom_1(51600) <= 9191156;
srom_1(51601) <= 8617803;
srom_1(51602) <= 8043375;
srom_1(51603) <= 7470566;
srom_1(51604) <= 6902063;
srom_1(51605) <= 6340530;
srom_1(51606) <= 5788601;
srom_1(51607) <= 5248864;
srom_1(51608) <= 4723851;
srom_1(51609) <= 4216023;
srom_1(51610) <= 3727762;
srom_1(51611) <= 3261357;
srom_1(51612) <= 2818995;
srom_1(51613) <= 2402752;
srom_1(51614) <= 2014578;
srom_1(51615) <= 1656294;
srom_1(51616) <= 1329580;
srom_1(51617) <= 1035968;
srom_1(51618) <= 776836;
srom_1(51619) <= 553397;
srom_1(51620) <= 366701;
srom_1(51621) <= 217622;
srom_1(51622) <= 106860;
srom_1(51623) <= 34933;
srom_1(51624) <= 2180;
srom_1(51625) <= 8754;
srom_1(51626) <= 54624;
srom_1(51627) <= 139574;
srom_1(51628) <= 263207;
srom_1(51629) <= 424943;
srom_1(51630) <= 624024;
srom_1(51631) <= 859515;
srom_1(51632) <= 1130312;
srom_1(51633) <= 1435146;
srom_1(51634) <= 1772588;
srom_1(51635) <= 2141054;
srom_1(51636) <= 2538817;
srom_1(51637) <= 2964012;
srom_1(51638) <= 3414644;
srom_1(51639) <= 3888602;
srom_1(51640) <= 4383661;
srom_1(51641) <= 4897501;
srom_1(51642) <= 5427711;
srom_1(51643) <= 5971807;
srom_1(51644) <= 6527236;
srom_1(51645) <= 7091393;
srom_1(51646) <= 7661633;
srom_1(51647) <= 8235283;
srom_1(51648) <= 8809651;
srom_1(51649) <= 9382045;
srom_1(51650) <= 9949780;
srom_1(51651) <= 10510195;
srom_1(51652) <= 11060660;
srom_1(51653) <= 11598596;
srom_1(51654) <= 12121478;
srom_1(51655) <= 12626856;
srom_1(51656) <= 13112360;
srom_1(51657) <= 13575712;
srom_1(51658) <= 14014740;
srom_1(51659) <= 14427385;
srom_1(51660) <= 14811712;
srom_1(51661) <= 15165919;
srom_1(51662) <= 15488345;
srom_1(51663) <= 15777478;
srom_1(51664) <= 16031962;
srom_1(51665) <= 16250603;
srom_1(51666) <= 16432377;
srom_1(51667) <= 16576431;
srom_1(51668) <= 16682089;
srom_1(51669) <= 16748857;
srom_1(51670) <= 16776420;
srom_1(51671) <= 16764650;
srom_1(51672) <= 16713602;
srom_1(51673) <= 16623515;
srom_1(51674) <= 16494811;
srom_1(51675) <= 16328095;
srom_1(51676) <= 16124148;
srom_1(51677) <= 15883927;
srom_1(51678) <= 15608557;
srom_1(51679) <= 15299330;
srom_1(51680) <= 14957697;
srom_1(51681) <= 14585259;
srom_1(51682) <= 14183763;
srom_1(51683) <= 13755091;
srom_1(51684) <= 13301254;
srom_1(51685) <= 12824379;
srom_1(51686) <= 12326704;
srom_1(51687) <= 11810562;
srom_1(51688) <= 11278373;
srom_1(51689) <= 10732633;
srom_1(51690) <= 10175901;
srom_1(51691) <= 9610788;
srom_1(51692) <= 9039944;
srom_1(51693) <= 8466045;
srom_1(51694) <= 7891783;
srom_1(51695) <= 7319851;
srom_1(51696) <= 6752931;
srom_1(51697) <= 6193681;
srom_1(51698) <= 5644723;
srom_1(51699) <= 5108633;
srom_1(51700) <= 4587924;
srom_1(51701) <= 4085037;
srom_1(51702) <= 3602331;
srom_1(51703) <= 3142070;
srom_1(51704) <= 2706411;
srom_1(51705) <= 2297399;
srom_1(51706) <= 1916950;
srom_1(51707) <= 1566849;
srom_1(51708) <= 1248737;
srom_1(51709) <= 964107;
srom_1(51710) <= 714293;
srom_1(51711) <= 500466;
srom_1(51712) <= 323629;
srom_1(51713) <= 184612;
srom_1(51714) <= 84067;
srom_1(51715) <= 22464;
srom_1(51716) <= 92;
srom_1(51717) <= 17058;
srom_1(51718) <= 73280;
srom_1(51719) <= 168496;
srom_1(51720) <= 302259;
srom_1(51721) <= 473942;
srom_1(51722) <= 682739;
srom_1(51723) <= 927671;
srom_1(51724) <= 1207591;
srom_1(51725) <= 1521185;
srom_1(51726) <= 1866982;
srom_1(51727) <= 2243361;
srom_1(51728) <= 2648558;
srom_1(51729) <= 3080672;
srom_1(51730) <= 3537676;
srom_1(51731) <= 4017429;
srom_1(51732) <= 4517679;
srom_1(51733) <= 5036081;
srom_1(51734) <= 5570204;
srom_1(51735) <= 6117544;
srom_1(51736) <= 6675534;
srom_1(51737) <= 7241557;
srom_1(51738) <= 7812958;
srom_1(51739) <= 8387059;
srom_1(51740) <= 8961168;
srom_1(51741) <= 9532591;
srom_1(51742) <= 10098650;
srom_1(51743) <= 10656690;
srom_1(51744) <= 11204094;
srom_1(51745) <= 11738296;
srom_1(51746) <= 12256789;
srom_1(51747) <= 12757143;
srom_1(51748) <= 13237012;
srom_1(51749) <= 13694145;
srom_1(51750) <= 14126398;
srom_1(51751) <= 14531745;
srom_1(51752) <= 14908285;
srom_1(51753) <= 15254251;
srom_1(51754) <= 15568022;
srom_1(51755) <= 15848127;
srom_1(51756) <= 16093251;
srom_1(51757) <= 16302245;
srom_1(51758) <= 16474130;
srom_1(51759) <= 16608099;
srom_1(51760) <= 16703524;
srom_1(51761) <= 16759957;
srom_1(51762) <= 16777135;
srom_1(51763) <= 16754975;
srom_1(51764) <= 16693583;
srom_1(51765) <= 16593246;
srom_1(51766) <= 16454434;
srom_1(51767) <= 16277799;
srom_1(51768) <= 16064169;
srom_1(51769) <= 15814546;
srom_1(51770) <= 15530100;
srom_1(51771) <= 15212165;
srom_1(51772) <= 14862231;
srom_1(51773) <= 14481941;
srom_1(51774) <= 14073077;
srom_1(51775) <= 13637557;
srom_1(51776) <= 13177423;
srom_1(51777) <= 12694832;
srom_1(51778) <= 12192047;
srom_1(51779) <= 11671427;
srom_1(51780) <= 11135413;
srom_1(51781) <= 10586518;
srom_1(51782) <= 10027317;
srom_1(51783) <= 9460431;
srom_1(51784) <= 8888518;
srom_1(51785) <= 8314262;
srom_1(51786) <= 7740354;
srom_1(51787) <= 7169486;
srom_1(51788) <= 6604335;
srom_1(51789) <= 6047551;
srom_1(51790) <= 5501745;
srom_1(51791) <= 4969476;
srom_1(51792) <= 4453241;
srom_1(51793) <= 3955460;
srom_1(51794) <= 3478468;
srom_1(51795) <= 3024501;
srom_1(51796) <= 2595688;
srom_1(51797) <= 2194040;
srom_1(51798) <= 1821441;
srom_1(51799) <= 1479637;
srom_1(51800) <= 1170232;
srom_1(51801) <= 894676;
srom_1(51802) <= 654262;
srom_1(51803) <= 450117;
srom_1(51804) <= 283198;
srom_1(51805) <= 154288;
srom_1(51806) <= 63992;
srom_1(51807) <= 12733;
srom_1(51808) <= 751;
srom_1(51809) <= 28103;
srom_1(51810) <= 94660;
srom_1(51811) <= 200110;
srom_1(51812) <= 343958;
srom_1(51813) <= 525531;
srom_1(51814) <= 743977;
srom_1(51815) <= 998271;
srom_1(51816) <= 1287220;
srom_1(51817) <= 1609471;
srom_1(51818) <= 1963511;
srom_1(51819) <= 2347681;
srom_1(51820) <= 2760178;
srom_1(51821) <= 3199070;
srom_1(51822) <= 3662297;
srom_1(51823) <= 4147687;
srom_1(51824) <= 4652964;
srom_1(51825) <= 5175759;
srom_1(51826) <= 5713620;
srom_1(51827) <= 6264025;
srom_1(51828) <= 6824393;
srom_1(51829) <= 7392096;
srom_1(51830) <= 7964472;
srom_1(51831) <= 8538837;
srom_1(51832) <= 9112497;
srom_1(51833) <= 9682763;
srom_1(51834) <= 10246960;
srom_1(51835) <= 10802443;
srom_1(51836) <= 11346606;
srom_1(51837) <= 11876899;
srom_1(51838) <= 12390833;
srom_1(51839) <= 12886000;
srom_1(51840) <= 13360077;
srom_1(51841) <= 13810841;
srom_1(51842) <= 14236178;
srom_1(51843) <= 14634094;
srom_1(51844) <= 15002722;
srom_1(51845) <= 15340335;
srom_1(51846) <= 15645349;
srom_1(51847) <= 15916333;
srom_1(51848) <= 16152018;
srom_1(51849) <= 16351297;
srom_1(51850) <= 16513236;
srom_1(51851) <= 16637076;
srom_1(51852) <= 16722236;
srom_1(51853) <= 16768317;
srom_1(51854) <= 16775103;
srom_1(51855) <= 16742561;
srom_1(51856) <= 16670845;
srom_1(51857) <= 16560291;
srom_1(51858) <= 16411416;
srom_1(51859) <= 16224920;
srom_1(51860) <= 16001677;
srom_1(51861) <= 15742734;
srom_1(51862) <= 15449304;
srom_1(51863) <= 15122765;
srom_1(51864) <= 14764646;
srom_1(51865) <= 14376629;
srom_1(51866) <= 13960531;
srom_1(51867) <= 13518305;
srom_1(51868) <= 13052024;
srom_1(51869) <= 12563874;
srom_1(51870) <= 12056145;
srom_1(51871) <= 11531218;
srom_1(51872) <= 10991554;
srom_1(51873) <= 10439684;
srom_1(51874) <= 9878196;
srom_1(51875) <= 9309722;
srom_1(51876) <= 8736929;
srom_1(51877) <= 8162503;
srom_1(51878) <= 7589137;
srom_1(51879) <= 7019520;
srom_1(51880) <= 6456323;
srom_1(51881) <= 5902187;
srom_1(51882) <= 5359711;
srom_1(51883) <= 4831438;
srom_1(51884) <= 4319846;
srom_1(51885) <= 3827334;
srom_1(51886) <= 3356212;
srom_1(51887) <= 2908688;
srom_1(51888) <= 2486861;
srom_1(51889) <= 2092710;
srom_1(51890) <= 1728082;
srom_1(51891) <= 1394687;
srom_1(51892) <= 1094090;
srom_1(51893) <= 827699;
srom_1(51894) <= 596764;
srom_1(51895) <= 402367;
srom_1(51896) <= 245421;
srom_1(51897) <= 126660;
srom_1(51898) <= 46643;
srom_1(51899) <= 5744;
srom_1(51900) <= 4156;
srom_1(51901) <= 41885;
srom_1(51902) <= 118754;
srom_1(51903) <= 234404;
srom_1(51904) <= 388292;
srom_1(51905) <= 579695;
srom_1(51906) <= 807718;
srom_1(51907) <= 1071290;
srom_1(51908) <= 1369175;
srom_1(51909) <= 1699977;
srom_1(51910) <= 2062144;
srom_1(51911) <= 2453978;
srom_1(51912) <= 2873641;
srom_1(51913) <= 3319167;
srom_1(51914) <= 3788464;
srom_1(51915) <= 4279333;
srom_1(51916) <= 4789472;
srom_1(51917) <= 5316489;
srom_1(51918) <= 5857911;
srom_1(51919) <= 6411201;
srom_1(51920) <= 6973764;
srom_1(51921) <= 7542961;
srom_1(51922) <= 8116124;
srom_1(51923) <= 8690565;
srom_1(51924) <= 9263590;
srom_1(51925) <= 9832511;
srom_1(51926) <= 10394662;
srom_1(51927) <= 10947406;
srom_1(51928) <= 11488150;
srom_1(51929) <= 12014360;
srom_1(51930) <= 12523567;
srom_1(51931) <= 13013384;
srom_1(51932) <= 13481514;
srom_1(51933) <= 13925761;
srom_1(51934) <= 14344043;
srom_1(51935) <= 14734398;
srom_1(51936) <= 15094995;
srom_1(51937) <= 15424144;
srom_1(51938) <= 15720300;
srom_1(51939) <= 15982076;
srom_1(51940) <= 16208243;
srom_1(51941) <= 16397741;
srom_1(51942) <= 16549682;
srom_1(51943) <= 16663353;
srom_1(51944) <= 16738220;
srom_1(51945) <= 16773934;
srom_1(51946) <= 16770325;
srom_1(51947) <= 16727412;
srom_1(51948) <= 16645396;
srom_1(51949) <= 16524660;
srom_1(51950) <= 16365772;
srom_1(51951) <= 16169476;
srom_1(51952) <= 15936693;
srom_1(51953) <= 15668514;
srom_1(51954) <= 15366197;
srom_1(51955) <= 15031160;
srom_1(51956) <= 14664974;
srom_1(51957) <= 14269356;
srom_1(51958) <= 13846161;
srom_1(51959) <= 13397373;
srom_1(51960) <= 12925098;
srom_1(51961) <= 12431549;
srom_1(51962) <= 11919042;
srom_1(51963) <= 11389980;
srom_1(51964) <= 10846842;
srom_1(51965) <= 10292178;
srom_1(51966) <= 9728587;
srom_1(51967) <= 9158712;
srom_1(51968) <= 8585226;
srom_1(51969) <= 8010818;
srom_1(51970) <= 7438181;
srom_1(51971) <= 6870002;
srom_1(51972) <= 6308943;
srom_1(51973) <= 5757637;
srom_1(51974) <= 5218669;
srom_1(51975) <= 4694565;
srom_1(51976) <= 4187784;
srom_1(51977) <= 3700702;
srom_1(51978) <= 3235603;
srom_1(51979) <= 2794669;
srom_1(51980) <= 2379966;
srom_1(51981) <= 1993440;
srom_1(51982) <= 1636903;
srom_1(51983) <= 1312027;
srom_1(51984) <= 1020336;
srom_1(51985) <= 763197;
srom_1(51986) <= 541816;
srom_1(51987) <= 357232;
srom_1(51988) <= 210309;
srom_1(51989) <= 101737;
srom_1(51990) <= 32025;
srom_1(51991) <= 1500;
srom_1(51992) <= 10306;
srom_1(51993) <= 58399;
srom_1(51994) <= 145556;
srom_1(51995) <= 271368;
srom_1(51996) <= 435244;
srom_1(51997) <= 636416;
srom_1(51998) <= 873941;
srom_1(51999) <= 1146704;
srom_1(52000) <= 1453428;
srom_1(52001) <= 1792672;
srom_1(52002) <= 2162848;
srom_1(52003) <= 2562218;
srom_1(52004) <= 2988910;
srom_1(52005) <= 3440923;
srom_1(52006) <= 3916138;
srom_1(52007) <= 4412325;
srom_1(52008) <= 4927159;
srom_1(52009) <= 5458224;
srom_1(52010) <= 6003031;
srom_1(52011) <= 6559025;
srom_1(52012) <= 7123598;
srom_1(52013) <= 7694104;
srom_1(52014) <= 8267866;
srom_1(52015) <= 8842194;
srom_1(52016) <= 9414396;
srom_1(52017) <= 9981787;
srom_1(52018) <= 10541707;
srom_1(52019) <= 11091530;
srom_1(52020) <= 11628679;
srom_1(52021) <= 12150634;
srom_1(52022) <= 12654947;
srom_1(52023) <= 13139254;
srom_1(52024) <= 13601284;
srom_1(52025) <= 14038869;
srom_1(52026) <= 14449959;
srom_1(52027) <= 14832624;
srom_1(52028) <= 15185072;
srom_1(52029) <= 15505648;
srom_1(52030) <= 15792851;
srom_1(52031) <= 16045332;
srom_1(52032) <= 16261908;
srom_1(52033) <= 16441564;
srom_1(52034) <= 16583456;
srom_1(52035) <= 16686920;
srom_1(52036) <= 16751471;
srom_1(52037) <= 16776805;
srom_1(52038) <= 16762804;
srom_1(52039) <= 16709533;
srom_1(52040) <= 16617243;
srom_1(52041) <= 16486366;
srom_1(52042) <= 16317516;
srom_1(52043) <= 16111484;
srom_1(52044) <= 15869237;
srom_1(52045) <= 15591911;
srom_1(52046) <= 15280806;
srom_1(52047) <= 14937381;
srom_1(52048) <= 14563247;
srom_1(52049) <= 14160157;
srom_1(52050) <= 13730003;
srom_1(52051) <= 13274802;
srom_1(52052) <= 12796687;
srom_1(52053) <= 12297901;
srom_1(52054) <= 11780783;
srom_1(52055) <= 11247758;
srom_1(52056) <= 10701326;
srom_1(52057) <= 10144049;
srom_1(52058) <= 9578539;
srom_1(52059) <= 9007450;
srom_1(52060) <= 8433458;
srom_1(52061) <= 7859257;
srom_1(52062) <= 7287537;
srom_1(52063) <= 6720981;
srom_1(52064) <= 6162245;
srom_1(52065) <= 5613949;
srom_1(52066) <= 5078664;
srom_1(52067) <= 4558901;
srom_1(52068) <= 4057097;
srom_1(52069) <= 3575605;
srom_1(52070) <= 3116682;
srom_1(52071) <= 2682481;
srom_1(52072) <= 2275039;
srom_1(52073) <= 1896265;
srom_1(52074) <= 1547935;
srom_1(52075) <= 1231684;
srom_1(52076) <= 948995;
srom_1(52077) <= 701192;
srom_1(52078) <= 489438;
srom_1(52079) <= 314726;
srom_1(52080) <= 177875;
srom_1(52081) <= 79527;
srom_1(52082) <= 20143;
srom_1(52083) <= 2;
srom_1(52084) <= 19198;
srom_1(52085) <= 77641;
srom_1(52086) <= 175057;
srom_1(52087) <= 310989;
srom_1(52088) <= 484800;
srom_1(52089) <= 695674;
srom_1(52090) <= 942624;
srom_1(52091) <= 1224490;
srom_1(52092) <= 1539951;
srom_1(52093) <= 1887527;
srom_1(52094) <= 2265590;
srom_1(52095) <= 2672365;
srom_1(52096) <= 3105946;
srom_1(52097) <= 3564299;
srom_1(52098) <= 4045275;
srom_1(52099) <= 4546619;
srom_1(52100) <= 5065978;
srom_1(52101) <= 5600919;
srom_1(52102) <= 6148932;
srom_1(52103) <= 6707448;
srom_1(52104) <= 7273847;
srom_1(52105) <= 7845474;
srom_1(52106) <= 8419647;
srom_1(52107) <= 8993675;
srom_1(52108) <= 9564866;
srom_1(52109) <= 10130541;
srom_1(52110) <= 10688047;
srom_1(52111) <= 11234770;
srom_1(52112) <= 11768147;
srom_1(52113) <= 12285676;
srom_1(52114) <= 12784930;
srom_1(52115) <= 13263569;
srom_1(52116) <= 13719347;
srom_1(52117) <= 14150127;
srom_1(52118) <= 14553890;
srom_1(52119) <= 14928741;
srom_1(52120) <= 15272924;
srom_1(52121) <= 15584823;
srom_1(52122) <= 15862977;
srom_1(52123) <= 16106081;
srom_1(52124) <= 16312996;
srom_1(52125) <= 16482750;
srom_1(52126) <= 16614548;
srom_1(52127) <= 16707771;
srom_1(52128) <= 16761983;
srom_1(52129) <= 16776930;
srom_1(52130) <= 16752541;
srom_1(52131) <= 16688930;
srom_1(52132) <= 16586396;
srom_1(52133) <= 16445421;
srom_1(52134) <= 16266664;
srom_1(52135) <= 16050964;
srom_1(52136) <= 15799332;
srom_1(52137) <= 15512949;
srom_1(52138) <= 15193158;
srom_1(52139) <= 14841458;
srom_1(52140) <= 14459498;
srom_1(52141) <= 14049070;
srom_1(52142) <= 13612097;
srom_1(52143) <= 13150631;
srom_1(52144) <= 12666833;
srom_1(52145) <= 12162973;
srom_1(52146) <= 11641414;
srom_1(52147) <= 11104601;
srom_1(52148) <= 10555053;
srom_1(52149) <= 9995345;
srom_1(52150) <= 9428102;
srom_1(52151) <= 8855985;
srom_1(52152) <= 8281676;
srom_1(52153) <= 7707869;
srom_1(52154) <= 7137253;
srom_1(52155) <= 6572506;
srom_1(52156) <= 6016275;
srom_1(52157) <= 5471169;
srom_1(52158) <= 4939744;
srom_1(52159) <= 4424491;
srom_1(52160) <= 3927828;
srom_1(52161) <= 3452083;
srom_1(52162) <= 2999487;
srom_1(52163) <= 2572162;
srom_1(52164) <= 2172113;
srom_1(52165) <= 1801215;
srom_1(52166) <= 1461207;
srom_1(52167) <= 1153684;
srom_1(52168) <= 880089;
srom_1(52169) <= 641703;
srom_1(52170) <= 439646;
srom_1(52171) <= 274863;
srom_1(52172) <= 148129;
srom_1(52173) <= 60037;
srom_1(52174) <= 11001;
srom_1(52175) <= 1251;
srom_1(52176) <= 30831;
srom_1(52177) <= 99604;
srom_1(52178) <= 207247;
srom_1(52179) <= 353255;
srom_1(52180) <= 536944;
srom_1(52181) <= 757452;
srom_1(52182) <= 1013745;
srom_1(52183) <= 1304621;
srom_1(52184) <= 1628716;
srom_1(52185) <= 1984511;
srom_1(52186) <= 2370337;
srom_1(52187) <= 2784384;
srom_1(52188) <= 3224712;
srom_1(52189) <= 3689255;
srom_1(52190) <= 4175835;
srom_1(52191) <= 4682170;
srom_1(52192) <= 5205886;
srom_1(52193) <= 5744527;
srom_1(52194) <= 6295566;
srom_1(52195) <= 6856421;
srom_1(52196) <= 7424460;
srom_1(52197) <= 7997021;
srom_1(52198) <= 8571418;
srom_1(52199) <= 9144958;
srom_1(52200) <= 9714951;
srom_1(52201) <= 10278724;
srom_1(52202) <= 10833634;
srom_1(52203) <= 11377079;
srom_1(52204) <= 11906509;
srom_1(52205) <= 12419443;
srom_1(52206) <= 12913474;
srom_1(52207) <= 13386287;
srom_1(52208) <= 13835665;
srom_1(52209) <= 14259499;
srom_1(52210) <= 14655802;
srom_1(52211) <= 15022717;
srom_1(52212) <= 15358521;
srom_1(52213) <= 15661642;
srom_1(52214) <= 15930657;
srom_1(52215) <= 16164304;
srom_1(52216) <= 16361489;
srom_1(52217) <= 16521286;
srom_1(52218) <= 16642946;
srom_1(52219) <= 16725898;
srom_1(52220) <= 16769754;
srom_1(52221) <= 16774309;
srom_1(52222) <= 16739539;
srom_1(52223) <= 16665609;
srom_1(52224) <= 16552866;
srom_1(52225) <= 16401838;
srom_1(52226) <= 16213232;
srom_1(52227) <= 15987935;
srom_1(52228) <= 15727001;
srom_1(52229) <= 15431655;
srom_1(52230) <= 15103282;
srom_1(52231) <= 14743422;
srom_1(52232) <= 14353762;
srom_1(52233) <= 13936129;
srom_1(52234) <= 13492481;
srom_1(52235) <= 13024900;
srom_1(52236) <= 12535578;
srom_1(52237) <= 12026809;
srom_1(52238) <= 11500980;
srom_1(52239) <= 10960555;
srom_1(52240) <= 10408070;
srom_1(52241) <= 9846114;
srom_1(52242) <= 9277324;
srom_1(52243) <= 8704367;
srom_1(52244) <= 8129929;
srom_1(52245) <= 7556703;
srom_1(52246) <= 6987379;
srom_1(52247) <= 6424626;
srom_1(52248) <= 5871082;
srom_1(52249) <= 5329344;
srom_1(52250) <= 4801952;
srom_1(52251) <= 4291379;
srom_1(52252) <= 3800020;
srom_1(52253) <= 3330177;
srom_1(52254) <= 2884056;
srom_1(52255) <= 2463747;
srom_1(52256) <= 2071222;
srom_1(52257) <= 1708321;
srom_1(52258) <= 1376747;
srom_1(52259) <= 1078053;
srom_1(52260) <= 813641;
srom_1(52261) <= 584751;
srom_1(52262) <= 392456;
srom_1(52263) <= 237657;
srom_1(52264) <= 121081;
srom_1(52265) <= 43274;
srom_1(52266) <= 4602;
srom_1(52267) <= 5245;
srom_1(52268) <= 45200;
srom_1(52269) <= 124281;
srom_1(52270) <= 242115;
srom_1(52271) <= 398152;
srom_1(52272) <= 591658;
srom_1(52273) <= 821727;
srom_1(52274) <= 1087280;
srom_1(52275) <= 1387071;
srom_1(52276) <= 1719695;
srom_1(52277) <= 2083591;
srom_1(52278) <= 2477054;
srom_1(52279) <= 2898238;
srom_1(52280) <= 3345169;
srom_1(52281) <= 3815750;
srom_1(52282) <= 4307774;
srom_1(52283) <= 4818935;
srom_1(52284) <= 5346835;
srom_1(52285) <= 5889000;
srom_1(52286) <= 6442886;
srom_1(52287) <= 7005896;
srom_1(52288) <= 7575390;
srom_1(52289) <= 8148697;
srom_1(52290) <= 8723129;
srom_1(52291) <= 9295993;
srom_1(52292) <= 9864602;
srom_1(52293) <= 10426289;
srom_1(52294) <= 10978421;
srom_1(52295) <= 11518408;
srom_1(52296) <= 12043719;
srom_1(52297) <= 12551889;
srom_1(52298) <= 13040537;
srom_1(52299) <= 13507370;
srom_1(52300) <= 13950199;
srom_1(52301) <= 14366948;
srom_1(52302) <= 14755663;
srom_1(52303) <= 15114520;
srom_1(52304) <= 15441837;
srom_1(52305) <= 15736080;
srom_1(52306) <= 15995867;
srom_1(52307) <= 16219981;
srom_1(52308) <= 16407371;
srom_1(52309) <= 16557159;
srom_1(52310) <= 16668641;
srom_1(52311) <= 16741296;
srom_1(52312) <= 16774782;
srom_1(52313) <= 16768942;
srom_1(52314) <= 16723804;
srom_1(52315) <= 16639579;
srom_1(52316) <= 16516663;
srom_1(52317) <= 16355631;
srom_1(52318) <= 16157239;
srom_1(52319) <= 15922418;
srom_1(52320) <= 15652268;
srom_1(52321) <= 15348056;
srom_1(52322) <= 15011208;
srom_1(52323) <= 14643306;
srom_1(52324) <= 14246072;
srom_1(52325) <= 13821371;
srom_1(52326) <= 13371194;
srom_1(52327) <= 12897652;
srom_1(52328) <= 12402966;
srom_1(52329) <= 11889454;
srom_1(52330) <= 11359526;
srom_1(52331) <= 10815667;
srom_1(52332) <= 10260426;
srom_1(52333) <= 9696407;
srom_1(52334) <= 9126256;
srom_1(52335) <= 8552646;
srom_1(52336) <= 7978266;
srom_1(52337) <= 7405811;
srom_1(52338) <= 6837964;
srom_1(52339) <= 6277389;
srom_1(52340) <= 5726714;
srom_1(52341) <= 5188521;
srom_1(52342) <= 4665335;
srom_1(52343) <= 4159609;
srom_1(52344) <= 3673713;
srom_1(52345) <= 3209928;
srom_1(52346) <= 2770427;
srom_1(52347) <= 2357272;
srom_1(52348) <= 1972399;
srom_1(52349) <= 1617615;
srom_1(52350) <= 1294582;
srom_1(52351) <= 1004815;
srom_1(52352) <= 749674;
srom_1(52353) <= 530354;
srom_1(52354) <= 347884;
srom_1(52355) <= 203120;
srom_1(52356) <= 96740;
srom_1(52357) <= 29244;
srom_1(52358) <= 947;
srom_1(52359) <= 11984;
srom_1(52360) <= 62301;
srom_1(52361) <= 151663;
srom_1(52362) <= 279651;
srom_1(52363) <= 445664;
srom_1(52364) <= 648925;
srom_1(52365) <= 888480;
srom_1(52366) <= 1163206;
srom_1(52367) <= 1471813;
srom_1(52368) <= 1812856;
srom_1(52369) <= 2184736;
srom_1(52370) <= 2585707;
srom_1(52371) <= 3013890;
srom_1(52372) <= 3467276;
srom_1(52373) <= 3943741;
srom_1(52374) <= 4441049;
srom_1(52375) <= 4956869;
srom_1(52376) <= 5488781;
srom_1(52377) <= 6034291;
srom_1(52378) <= 6590842;
srom_1(52379) <= 7155823;
srom_1(52380) <= 7726585;
srom_1(52381) <= 8300451;
srom_1(52382) <= 8874731;
srom_1(52383) <= 9446731;
srom_1(52384) <= 10013769;
srom_1(52385) <= 10573187;
srom_1(52386) <= 11122360;
srom_1(52387) <= 11658713;
srom_1(52388) <= 12179732;
srom_1(52389) <= 12682973;
srom_1(52390) <= 13166076;
srom_1(52391) <= 13626777;
srom_1(52392) <= 14062913;
srom_1(52393) <= 14472441;
srom_1(52394) <= 14853439;
srom_1(52395) <= 15204122;
srom_1(52396) <= 15522844;
srom_1(52397) <= 15808112;
srom_1(52398) <= 16058587;
srom_1(52399) <= 16273094;
srom_1(52400) <= 16450629;
srom_1(52401) <= 16590358;
srom_1(52402) <= 16691626;
srom_1(52403) <= 16753959;
srom_1(52404) <= 16777063;
srom_1(52405) <= 16760831;
srom_1(52406) <= 16705339;
srom_1(52407) <= 16610847;
srom_1(52408) <= 16477798;
srom_1(52409) <= 16306816;
srom_1(52410) <= 16098703;
srom_1(52411) <= 15854434;
srom_1(52412) <= 15575156;
srom_1(52413) <= 15262177;
srom_1(52414) <= 14916966;
srom_1(52415) <= 14541142;
srom_1(52416) <= 14136465;
srom_1(52417) <= 13704836;
srom_1(52418) <= 13248276;
srom_1(52419) <= 12768928;
srom_1(52420) <= 12269039;
srom_1(52421) <= 11750953;
srom_1(52422) <= 11217100;
srom_1(52423) <= 10669984;
srom_1(52424) <= 10112169;
srom_1(52425) <= 9546272;
srom_1(52426) <= 8974946;
srom_1(52427) <= 8400871;
srom_1(52428) <= 7826738;
srom_1(52429) <= 7255240;
srom_1(52430) <= 6689056;
srom_1(52431) <= 6130843;
srom_1(52432) <= 5583216;
srom_1(52433) <= 5048746;
srom_1(52434) <= 4529937;
srom_1(52435) <= 4029222;
srom_1(52436) <= 3548951;
srom_1(52437) <= 3091374;
srom_1(52438) <= 2658638;
srom_1(52439) <= 2252771;
srom_1(52440) <= 1875677;
srom_1(52441) <= 1529125;
srom_1(52442) <= 1214740;
srom_1(52443) <= 933995;
srom_1(52444) <= 688207;
srom_1(52445) <= 478529;
srom_1(52446) <= 305944;
srom_1(52447) <= 171262;
srom_1(52448) <= 75113;
srom_1(52449) <= 17950;
srom_1(52450) <= 39;
srom_1(52451) <= 21465;
srom_1(52452) <= 82127;
srom_1(52453) <= 181742;
srom_1(52454) <= 319841;
srom_1(52455) <= 495778;
srom_1(52456) <= 708726;
srom_1(52457) <= 957688;
srom_1(52458) <= 1241497;
srom_1(52459) <= 1558820;
srom_1(52460) <= 1908171;
srom_1(52461) <= 2287911;
srom_1(52462) <= 2696259;
srom_1(52463) <= 3131301;
srom_1(52464) <= 3590995;
srom_1(52465) <= 4073188;
srom_1(52466) <= 4575617;
srom_1(52467) <= 5095926;
srom_1(52468) <= 5631676;
srom_1(52469) <= 6180354;
srom_1(52470) <= 6739387;
srom_1(52471) <= 7306154;
srom_1(52472) <= 7877997;
srom_1(52473) <= 8452234;
srom_1(52474) <= 9026174;
srom_1(52475) <= 9597123;
srom_1(52476) <= 10162405;
srom_1(52477) <= 10719369;
srom_1(52478) <= 11265404;
srom_1(52479) <= 11797948;
srom_1(52480) <= 12314504;
srom_1(52481) <= 12812651;
srom_1(52482) <= 13290052;
srom_1(52483) <= 13744468;
srom_1(52484) <= 14173769;
srom_1(52485) <= 14575941;
srom_1(52486) <= 14949099;
srom_1(52487) <= 15291492;
srom_1(52488) <= 15601515;
srom_1(52489) <= 15877715;
srom_1(52490) <= 16118795;
srom_1(52491) <= 16323626;
srom_1(52492) <= 16491247;
srom_1(52493) <= 16620872;
srom_1(52494) <= 16711893;
srom_1(52495) <= 16763883;
srom_1(52496) <= 16776599;
srom_1(52497) <= 16749980;
srom_1(52498) <= 16684152;
srom_1(52499) <= 16579423;
srom_1(52500) <= 16436285;
srom_1(52501) <= 16255409;
srom_1(52502) <= 16037642;
srom_1(52503) <= 15784007;
srom_1(52504) <= 15495692;
srom_1(52505) <= 15174049;
srom_1(52506) <= 14820587;
srom_1(52507) <= 14436963;
srom_1(52508) <= 14024977;
srom_1(52509) <= 13586559;
srom_1(52510) <= 13123767;
srom_1(52511) <= 12638770;
srom_1(52512) <= 12133842;
srom_1(52513) <= 11611351;
srom_1(52514) <= 11073748;
srom_1(52515) <= 10523554;
srom_1(52516) <= 9963348;
srom_1(52517) <= 9395757;
srom_1(52518) <= 8823444;
srom_1(52519) <= 8249092;
srom_1(52520) <= 7675393;
srom_1(52521) <= 7105040;
srom_1(52522) <= 6540705;
srom_1(52523) <= 5985036;
srom_1(52524) <= 5440638;
srom_1(52525) <= 4910064;
srom_1(52526) <= 4395802;
srom_1(52527) <= 3900263;
srom_1(52528) <= 3425773;
srom_1(52529) <= 2974554;
srom_1(52530) <= 2548724;
srom_1(52531) <= 2150279;
srom_1(52532) <= 1781088;
srom_1(52533) <= 1442881;
srom_1(52534) <= 1137246;
srom_1(52535) <= 865615;
srom_1(52536) <= 629261;
srom_1(52537) <= 429294;
srom_1(52538) <= 266651;
srom_1(52539) <= 142094;
srom_1(52540) <= 56208;
srom_1(52541) <= 9396;
srom_1(52542) <= 1877;
srom_1(52543) <= 33686;
srom_1(52544) <= 104673;
srom_1(52545) <= 214508;
srom_1(52546) <= 362673;
srom_1(52547) <= 548475;
srom_1(52548) <= 771041;
srom_1(52549) <= 1029330;
srom_1(52550) <= 1322128;
srom_1(52551) <= 1648063;
srom_1(52552) <= 2005608;
srom_1(52553) <= 2393084;
srom_1(52554) <= 2808675;
srom_1(52555) <= 3250433;
srom_1(52556) <= 3716285;
srom_1(52557) <= 4204047;
srom_1(52558) <= 4711432;
srom_1(52559) <= 5236061;
srom_1(52560) <= 5775473;
srom_1(52561) <= 6327139;
srom_1(52562) <= 6888472;
srom_1(52563) <= 7456839;
srom_1(52564) <= 8029576;
srom_1(52565) <= 8603997;
srom_1(52566) <= 9177407;
srom_1(52567) <= 9747119;
srom_1(52568) <= 10310460;
srom_1(52569) <= 10864789;
srom_1(52570) <= 11407506;
srom_1(52571) <= 11936066;
srom_1(52572) <= 12447991;
srom_1(52573) <= 12940881;
srom_1(52574) <= 13412423;
srom_1(52575) <= 13860406;
srom_1(52576) <= 14282731;
srom_1(52577) <= 14677416;
srom_1(52578) <= 15042611;
srom_1(52579) <= 15376602;
srom_1(52580) <= 15677825;
srom_1(52581) <= 15944866;
srom_1(52582) <= 16176473;
srom_1(52583) <= 16371560;
srom_1(52584) <= 16529212;
srom_1(52585) <= 16648691;
srom_1(52586) <= 16729434;
srom_1(52587) <= 16771065;
srom_1(52588) <= 16773388;
srom_1(52589) <= 16736391;
srom_1(52590) <= 16660249;
srom_1(52591) <= 16545318;
srom_1(52592) <= 16392138;
srom_1(52593) <= 16201426;
srom_1(52594) <= 15974077;
srom_1(52595) <= 15711158;
srom_1(52596) <= 15413900;
srom_1(52597) <= 15083699;
srom_1(52598) <= 14722102;
srom_1(52599) <= 14330805;
srom_1(52600) <= 13911642;
srom_1(52601) <= 13466581;
srom_1(52602) <= 12997707;
srom_1(52603) <= 12507220;
srom_1(52604) <= 11997419;
srom_1(52605) <= 11470694;
srom_1(52606) <= 10929517;
srom_1(52607) <= 10376425;
srom_1(52608) <= 9814011;
srom_1(52609) <= 9244913;
srom_1(52610) <= 8671800;
srom_1(52611) <= 8097358;
srom_1(52612) <= 7524283;
srom_1(52613) <= 6955260;
srom_1(52614) <= 6392959;
srom_1(52615) <= 5840016;
srom_1(52616) <= 5299024;
srom_1(52617) <= 4772521;
srom_1(52618) <= 4262974;
srom_1(52619) <= 3772774;
srom_1(52620) <= 3304219;
srom_1(52621) <= 2859507;
srom_1(52622) <= 2440722;
srom_1(52623) <= 2049830;
srom_1(52624) <= 1688661;
srom_1(52625) <= 1358912;
srom_1(52626) <= 1062127;
srom_1(52627) <= 799698;
srom_1(52628) <= 572856;
srom_1(52629) <= 382665;
srom_1(52630) <= 230017;
srom_1(52631) <= 115627;
srom_1(52632) <= 40032;
srom_1(52633) <= 3586;
srom_1(52634) <= 6460;
srom_1(52635) <= 48641;
srom_1(52636) <= 129932;
srom_1(52637) <= 249950;
srom_1(52638) <= 408133;
srom_1(52639) <= 603739;
srom_1(52640) <= 835851;
srom_1(52641) <= 1103380;
srom_1(52642) <= 1405073;
srom_1(52643) <= 1739513;
srom_1(52644) <= 2105134;
srom_1(52645) <= 2500219;
srom_1(52646) <= 2922918;
srom_1(52647) <= 3371247;
srom_1(52648) <= 3843104;
srom_1(52649) <= 4336277;
srom_1(52650) <= 4848452;
srom_1(52651) <= 5377228;
srom_1(52652) <= 5920126;
srom_1(52653) <= 6474599;
srom_1(52654) <= 7038048;
srom_1(52655) <= 7607830;
srom_1(52656) <= 8181273;
srom_1(52657) <= 8755689;
srom_1(52658) <= 9328383;
srom_1(52659) <= 9896670;
srom_1(52660) <= 10457885;
srom_1(52661) <= 11009397;
srom_1(52662) <= 11548619;
srom_1(52663) <= 12073023;
srom_1(52664) <= 12580149;
srom_1(52665) <= 13067620;
srom_1(52666) <= 13533149;
srom_1(52667) <= 13974553;
srom_1(52668) <= 14389763;
srom_1(52669) <= 14776832;
srom_1(52670) <= 15133944;
srom_1(52671) <= 15459425;
srom_1(52672) <= 15751748;
srom_1(52673) <= 16009543;
srom_1(52674) <= 16231601;
srom_1(52675) <= 16416881;
srom_1(52676) <= 16564513;
srom_1(52677) <= 16673805;
srom_1(52678) <= 16744245;
srom_1(52679) <= 16775503;
srom_1(52680) <= 16767432;
srom_1(52681) <= 16720069;
srom_1(52682) <= 16633638;
srom_1(52683) <= 16508542;
srom_1(52684) <= 16345370;
srom_1(52685) <= 16144885;
srom_1(52686) <= 15908029;
srom_1(52687) <= 15635912;
srom_1(52688) <= 15329809;
srom_1(52689) <= 14991157;
srom_1(52690) <= 14621543;
srom_1(52691) <= 14222701;
srom_1(52692) <= 13796500;
srom_1(52693) <= 13344940;
srom_1(52694) <= 12870139;
srom_1(52695) <= 12374321;
srom_1(52696) <= 11859814;
srom_1(52697) <= 11329028;
srom_1(52698) <= 10784454;
srom_1(52699) <= 10228646;
srom_1(52700) <= 9664208;
srom_1(52701) <= 9093789;
srom_1(52702) <= 8520063;
srom_1(52703) <= 7945720;
srom_1(52704) <= 7373455;
srom_1(52705) <= 6805949;
srom_1(52706) <= 6245866;
srom_1(52707) <= 5695830;
srom_1(52708) <= 5158422;
srom_1(52709) <= 4636161;
srom_1(52710) <= 4131497;
srom_1(52711) <= 3646796;
srom_1(52712) <= 3184330;
srom_1(52713) <= 2746270;
srom_1(52714) <= 2334668;
srom_1(52715) <= 1951455;
srom_1(52716) <= 1598429;
srom_1(52717) <= 1277243;
srom_1(52718) <= 989406;
srom_1(52719) <= 736265;
srom_1(52720) <= 519010;
srom_1(52721) <= 338657;
srom_1(52722) <= 196053;
srom_1(52723) <= 91868;
srom_1(52724) <= 26588;
srom_1(52725) <= 521;
srom_1(52726) <= 13788;
srom_1(52727) <= 66328;
srom_1(52728) <= 157894;
srom_1(52729) <= 288056;
srom_1(52730) <= 456205;
srom_1(52731) <= 661551;
srom_1(52732) <= 903133;
srom_1(52733) <= 1179816;
srom_1(52734) <= 1490304;
srom_1(52735) <= 1833140;
srom_1(52736) <= 2206717;
srom_1(52737) <= 2609283;
srom_1(52738) <= 3038950;
srom_1(52739) <= 3493704;
srom_1(52740) <= 3971412;
srom_1(52741) <= 4469833;
srom_1(52742) <= 4986631;
srom_1(52743) <= 5519381;
srom_1(52744) <= 6065587;
srom_1(52745) <= 6622686;
srom_1(52746) <= 7188066;
srom_1(52747) <= 7759076;
srom_1(52748) <= 8333038;
srom_1(52749) <= 8907260;
srom_1(52750) <= 9479051;
srom_1(52751) <= 10045728;
srom_1(52752) <= 10604634;
srom_1(52753) <= 11153148;
srom_1(52754) <= 11688698;
srom_1(52755) <= 12208774;
srom_1(52756) <= 12710935;
srom_1(52757) <= 13192827;
srom_1(52758) <= 13652190;
srom_1(52759) <= 14086871;
srom_1(52760) <= 14494831;
srom_1(52761) <= 14874156;
srom_1(52762) <= 15223069;
srom_1(52763) <= 15539932;
srom_1(52764) <= 15823261;
srom_1(52765) <= 16071726;
srom_1(52766) <= 16284162;
srom_1(52767) <= 16459573;
srom_1(52768) <= 16597136;
srom_1(52769) <= 16696207;
srom_1(52770) <= 16756320;
srom_1(52771) <= 16777195;
srom_1(52772) <= 16758733;
srom_1(52773) <= 16701020;
srom_1(52774) <= 16604327;
srom_1(52775) <= 16469108;
srom_1(52776) <= 16295997;
srom_1(52777) <= 16085805;
srom_1(52778) <= 15839519;
srom_1(52779) <= 15558293;
srom_1(52780) <= 15243445;
srom_1(52781) <= 14896453;
srom_1(52782) <= 14518943;
srom_1(52783) <= 14112686;
srom_1(52784) <= 13679587;
srom_1(52785) <= 13221677;
srom_1(52786) <= 12741103;
srom_1(52787) <= 12240118;
srom_1(52788) <= 11721072;
srom_1(52789) <= 11186400;
srom_1(52790) <= 10638607;
srom_1(52791) <= 10080264;
srom_1(52792) <= 9513987;
srom_1(52793) <= 8942434;
srom_1(52794) <= 8368283;
srom_1(52795) <= 7794227;
srom_1(52796) <= 7222959;
srom_1(52797) <= 6657157;
srom_1(52798) <= 6099474;
srom_1(52799) <= 5552526;
srom_1(52800) <= 5018877;
srom_1(52801) <= 4501030;
srom_1(52802) <= 4001414;
srom_1(52803) <= 3522370;
srom_1(52804) <= 3066146;
srom_1(52805) <= 2634880;
srom_1(52806) <= 2230596;
srom_1(52807) <= 1855189;
srom_1(52808) <= 1510419;
srom_1(52809) <= 1197903;
srom_1(52810) <= 919107;
srom_1(52811) <= 675338;
srom_1(52812) <= 467740;
srom_1(52813) <= 297285;
srom_1(52814) <= 164772;
srom_1(52815) <= 70825;
srom_1(52816) <= 15882;
srom_1(52817) <= 202;
srom_1(52818) <= 23858;
srom_1(52819) <= 86739;
srom_1(52820) <= 188550;
srom_1(52821) <= 328815;
srom_1(52822) <= 506874;
srom_1(52823) <= 721894;
srom_1(52824) <= 972865;
srom_1(52825) <= 1258612;
srom_1(52826) <= 1577793;
srom_1(52827) <= 1928913;
srom_1(52828) <= 2310324;
srom_1(52829) <= 2720239;
srom_1(52830) <= 3156734;
srom_1(52831) <= 3617764;
srom_1(52832) <= 4101165;
srom_1(52833) <= 4604672;
srom_1(52834) <= 5125923;
srom_1(52835) <= 5662474;
srom_1(52836) <= 6211809;
srom_1(52837) <= 6771351;
srom_1(52838) <= 7338477;
srom_1(52839) <= 7910528;
srom_1(52840) <= 8484821;
srom_1(52841) <= 9058662;
srom_1(52842) <= 9629362;
srom_1(52843) <= 10194242;
srom_1(52844) <= 10750656;
srom_1(52845) <= 11295993;
srom_1(52846) <= 11827697;
srom_1(52847) <= 12343273;
srom_1(52848) <= 12840305;
srom_1(52849) <= 13316461;
srom_1(52850) <= 13769509;
srom_1(52851) <= 14197324;
srom_1(52852) <= 14597899;
srom_1(52853) <= 14969358;
srom_1(52854) <= 15309956;
srom_1(52855) <= 15618099;
srom_1(52856) <= 15892339;
srom_1(52857) <= 16131392;
srom_1(52858) <= 16334137;
srom_1(52859) <= 16499622;
srom_1(52860) <= 16627072;
srom_1(52861) <= 16715889;
srom_1(52862) <= 16765656;
srom_1(52863) <= 16776141;
srom_1(52864) <= 16747293;
srom_1(52865) <= 16679249;
srom_1(52866) <= 16572327;
srom_1(52867) <= 16427029;
srom_1(52868) <= 16244035;
srom_1(52869) <= 16024205;
srom_1(52870) <= 15768570;
srom_1(52871) <= 15478326;
srom_1(52872) <= 15154837;
srom_1(52873) <= 14799619;
srom_1(52874) <= 14414337;
srom_1(52875) <= 14000798;
srom_1(52876) <= 13560942;
srom_1(52877) <= 13096831;
srom_1(52878) <= 12610642;
srom_1(52879) <= 12104654;
srom_1(52880) <= 11581240;
srom_1(52881) <= 11042855;
srom_1(52882) <= 10492023;
srom_1(52883) <= 9931328;
srom_1(52884) <= 9363398;
srom_1(52885) <= 8790897;
srom_1(52886) <= 8216509;
srom_1(52887) <= 7642929;
srom_1(52888) <= 7072845;
srom_1(52889) <= 6508932;
srom_1(52890) <= 5953832;
srom_1(52891) <= 5410151;
srom_1(52892) <= 4880436;
srom_1(52893) <= 4367172;
srom_1(52894) <= 3872767;
srom_1(52895) <= 3399537;
srom_1(52896) <= 2949703;
srom_1(52897) <= 2525374;
srom_1(52898) <= 2128540;
srom_1(52899) <= 1761061;
srom_1(52900) <= 1424661;
srom_1(52901) <= 1120917;
srom_1(52902) <= 851254;
srom_1(52903) <= 616936;
srom_1(52904) <= 419063;
srom_1(52905) <= 258561;
srom_1(52906) <= 136184;
srom_1(52907) <= 52505;
srom_1(52908) <= 7917;
srom_1(52909) <= 2629;
srom_1(52910) <= 36666;
srom_1(52911) <= 109868;
srom_1(52912) <= 221892;
srom_1(52913) <= 372212;
srom_1(52914) <= 560124;
srom_1(52915) <= 784746;
srom_1(52916) <= 1045026;
srom_1(52917) <= 1339742;
srom_1(52918) <= 1667512;
srom_1(52919) <= 2026800;
srom_1(52920) <= 2415921;
srom_1(52921) <= 2833050;
srom_1(52922) <= 3276231;
srom_1(52923) <= 3743385;
srom_1(52924) <= 4232322;
srom_1(52925) <= 4740750;
srom_1(52926) <= 5266284;
srom_1(52927) <= 5806459;
srom_1(52928) <= 6358743;
srom_1(52929) <= 6920546;
srom_1(52930) <= 7489233;
srom_1(52931) <= 8062137;
srom_1(52932) <= 8636572;
srom_1(52933) <= 9209845;
srom_1(52934) <= 9779266;
srom_1(52935) <= 10342166;
srom_1(52936) <= 10895906;
srom_1(52937) <= 11437887;
srom_1(52938) <= 11965570;
srom_1(52939) <= 12476479;
srom_1(52940) <= 12968218;
srom_1(52941) <= 13438482;
srom_1(52942) <= 13885066;
srom_1(52943) <= 14305874;
srom_1(52944) <= 14698935;
srom_1(52945) <= 15062404;
srom_1(52946) <= 15394578;
srom_1(52947) <= 15693898;
srom_1(52948) <= 15958961;
srom_1(52949) <= 16188524;
srom_1(52950) <= 16381511;
srom_1(52951) <= 16537016;
srom_1(52952) <= 16654311;
srom_1(52953) <= 16732845;
srom_1(52954) <= 16772249;
srom_1(52955) <= 16772340;
srom_1(52956) <= 16733117;
srom_1(52957) <= 16654764;
srom_1(52958) <= 16537647;
srom_1(52959) <= 16382317;
srom_1(52960) <= 16189502;
srom_1(52961) <= 15960106;
srom_1(52962) <= 15695204;
srom_1(52963) <= 15396039;
srom_1(52964) <= 15064014;
srom_1(52965) <= 14700686;
srom_1(52966) <= 14307758;
srom_1(52967) <= 13887073;
srom_1(52968) <= 13440604;
srom_1(52969) <= 12970444;
srom_1(52970) <= 12478799;
srom_1(52971) <= 11967973;
srom_1(52972) <= 11440363;
srom_1(52973) <= 10898441;
srom_1(52974) <= 10344751;
srom_1(52975) <= 9781887;
srom_1(52976) <= 9212489;
srom_1(52977) <= 8639229;
srom_1(52978) <= 8064792;
srom_1(52979) <= 7491875;
srom_1(52980) <= 6923162;
srom_1(52981) <= 6361322;
srom_1(52982) <= 5808988;
srom_1(52983) <= 5268750;
srom_1(52984) <= 4743143;
srom_1(52985) <= 4234631;
srom_1(52986) <= 3745598;
srom_1(52987) <= 3278338;
srom_1(52988) <= 2835041;
srom_1(52989) <= 2417788;
srom_1(52990) <= 2028533;
srom_1(52991) <= 1669103;
srom_1(52992) <= 1341183;
srom_1(52993) <= 1046311;
srom_1(52994) <= 785869;
srom_1(52995) <= 561079;
srom_1(52996) <= 372995;
srom_1(52997) <= 222499;
srom_1(52998) <= 110297;
srom_1(52999) <= 36915;
srom_1(53000) <= 2696;
srom_1(53001) <= 7802;
srom_1(53002) <= 52209;
srom_1(53003) <= 135707;
srom_1(53004) <= 257907;
srom_1(53005) <= 418234;
srom_1(53006) <= 615937;
srom_1(53007) <= 850088;
srom_1(53008) <= 1119590;
srom_1(53009) <= 1423180;
srom_1(53010) <= 1759432;
srom_1(53011) <= 2126771;
srom_1(53012) <= 2523474;
srom_1(53013) <= 2947680;
srom_1(53014) <= 3397401;
srom_1(53015) <= 3870527;
srom_1(53016) <= 4364840;
srom_1(53017) <= 4878022;
srom_1(53018) <= 5407667;
srom_1(53019) <= 5951290;
srom_1(53020) <= 6506342;
srom_1(53021) <= 7070221;
srom_1(53022) <= 7640282;
srom_1(53023) <= 8213853;
srom_1(53024) <= 8788242;
srom_1(53025) <= 9360758;
srom_1(53026) <= 9928715;
srom_1(53027) <= 10489451;
srom_1(53028) <= 11040334;
srom_1(53029) <= 11578783;
srom_1(53030) <= 12102271;
srom_1(53031) <= 12608345;
srom_1(53032) <= 13094632;
srom_1(53033) <= 13558850;
srom_1(53034) <= 13998823;
srom_1(53035) <= 14412488;
srom_1(53036) <= 14797905;
srom_1(53037) <= 15153266;
srom_1(53038) <= 15476906;
srom_1(53039) <= 15767306;
srom_1(53040) <= 16023105;
srom_1(53041) <= 16243103;
srom_1(53042) <= 16426268;
srom_1(53043) <= 16571743;
srom_1(53044) <= 16678843;
srom_1(53045) <= 16747068;
srom_1(53046) <= 16776098;
srom_1(53047) <= 16765795;
srom_1(53048) <= 16716209;
srom_1(53049) <= 16627572;
srom_1(53050) <= 16500300;
srom_1(53051) <= 16334989;
srom_1(53052) <= 16132415;
srom_1(53053) <= 15893527;
srom_1(53054) <= 15619446;
srom_1(53055) <= 15311458;
srom_1(53056) <= 14971005;
srom_1(53057) <= 14599686;
srom_1(53058) <= 14199241;
srom_1(53059) <= 13771547;
srom_1(53060) <= 13318612;
srom_1(53061) <= 12842557;
srom_1(53062) <= 12345617;
srom_1(53063) <= 11830121;
srom_1(53064) <= 11298486;
srom_1(53065) <= 10753206;
srom_1(53066) <= 10196838;
srom_1(53067) <= 9631990;
srom_1(53068) <= 9061311;
srom_1(53069) <= 8487478;
srom_1(53070) <= 7913181;
srom_1(53071) <= 7341114;
srom_1(53072) <= 6773959;
srom_1(53073) <= 6214375;
srom_1(53074) <= 5664987;
srom_1(53075) <= 5128372;
srom_1(53076) <= 4607044;
srom_1(53077) <= 4103450;
srom_1(53078) <= 3619950;
srom_1(53079) <= 3158812;
srom_1(53080) <= 2722198;
srom_1(53081) <= 2312156;
srom_1(53082) <= 1930608;
srom_1(53083) <= 1579345;
srom_1(53084) <= 1260012;
srom_1(53085) <= 974108;
srom_1(53086) <= 722973;
srom_1(53087) <= 507784;
srom_1(53088) <= 329552;
srom_1(53089) <= 189111;
srom_1(53090) <= 87121;
srom_1(53091) <= 24059;
srom_1(53092) <= 221;
srom_1(53093) <= 15719;
srom_1(53094) <= 70481;
srom_1(53095) <= 164249;
srom_1(53096) <= 296584;
srom_1(53097) <= 466865;
srom_1(53098) <= 674294;
srom_1(53099) <= 917898;
srom_1(53100) <= 1196535;
srom_1(53101) <= 1508898;
srom_1(53102) <= 1853522;
srom_1(53103) <= 2228792;
srom_1(53104) <= 2632946;
srom_1(53105) <= 3064092;
srom_1(53106) <= 3520205;
srom_1(53107) <= 3999149;
srom_1(53108) <= 4498676;
srom_1(53109) <= 5016444;
srom_1(53110) <= 5550025;
srom_1(53111) <= 6096918;
srom_1(53112) <= 6654557;
srom_1(53113) <= 7220328;
srom_1(53114) <= 7791577;
srom_1(53115) <= 8365625;
srom_1(53116) <= 8939782;
srom_1(53117) <= 9511354;
srom_1(53118) <= 10077661;
srom_1(53119) <= 10636047;
srom_1(53120) <= 11183894;
srom_1(53121) <= 11718634;
srom_1(53122) <= 12237757;
srom_1(53123) <= 12738831;
srom_1(53124) <= 13219505;
srom_1(53125) <= 13677525;
srom_1(53126) <= 14110744;
srom_1(53127) <= 14517129;
srom_1(53128) <= 14894776;
srom_1(53129) <= 15241913;
srom_1(53130) <= 15556913;
srom_1(53131) <= 15838298;
srom_1(53132) <= 16084749;
srom_1(53133) <= 16295110;
srom_1(53134) <= 16468394;
srom_1(53135) <= 16603790;
srom_1(53136) <= 16700662;
srom_1(53137) <= 16758556;
srom_1(53138) <= 16777200;
srom_1(53139) <= 16756507;
srom_1(53140) <= 16696575;
srom_1(53141) <= 16597683;
srom_1(53142) <= 16460296;
srom_1(53143) <= 16285059;
srom_1(53144) <= 16072792;
srom_1(53145) <= 15824491;
srom_1(53146) <= 15541321;
srom_1(53147) <= 15224610;
srom_1(53148) <= 14875842;
srom_1(53149) <= 14496653;
srom_1(53150) <= 14088821;
srom_1(53151) <= 13654259;
srom_1(53152) <= 13195005;
srom_1(53153) <= 12713212;
srom_1(53154) <= 12211139;
srom_1(53155) <= 11691141;
srom_1(53156) <= 11155657;
srom_1(53157) <= 10607197;
srom_1(53158) <= 10048333;
srom_1(53159) <= 9481686;
srom_1(53160) <= 8909913;
srom_1(53161) <= 8335695;
srom_1(53162) <= 7761726;
srom_1(53163) <= 7190696;
srom_1(53164) <= 6625284;
srom_1(53165) <= 6068141;
srom_1(53166) <= 5521879;
srom_1(53167) <= 4989060;
srom_1(53168) <= 4472183;
srom_1(53169) <= 3973671;
srom_1(53170) <= 3495862;
srom_1(53171) <= 3040998;
srom_1(53172) <= 2611209;
srom_1(53173) <= 2208514;
srom_1(53174) <= 1834798;
srom_1(53175) <= 1491816;
srom_1(53176) <= 1181175;
srom_1(53177) <= 904332;
srom_1(53178) <= 662586;
srom_1(53179) <= 457070;
srom_1(53180) <= 288747;
srom_1(53181) <= 158407;
srom_1(53182) <= 66662;
srom_1(53183) <= 13941;
srom_1(53184) <= 492;
srom_1(53185) <= 26377;
srom_1(53186) <= 91476;
srom_1(53187) <= 195483;
srom_1(53188) <= 337910;
srom_1(53189) <= 518090;
srom_1(53190) <= 735177;
srom_1(53191) <= 988154;
srom_1(53192) <= 1275834;
srom_1(53193) <= 1596868;
srom_1(53194) <= 1949752;
srom_1(53195) <= 2332829;
srom_1(53196) <= 2744304;
srom_1(53197) <= 3182246;
srom_1(53198) <= 3644604;
srom_1(53199) <= 4129207;
srom_1(53200) <= 4633785;
srom_1(53201) <= 5155970;
srom_1(53202) <= 5693314;
srom_1(53203) <= 6243297;
srom_1(53204) <= 6803340;
srom_1(53205) <= 7370817;
srom_1(53206) <= 7943067;
srom_1(53207) <= 8517406;
srom_1(53208) <= 9091141;
srom_1(53209) <= 9661581;
srom_1(53210) <= 10226053;
srom_1(53211) <= 10781908;
srom_1(53212) <= 11326539;
srom_1(53213) <= 11857394;
srom_1(53214) <= 12371983;
srom_1(53215) <= 12867892;
srom_1(53216) <= 13342796;
srom_1(53217) <= 13794468;
srom_1(53218) <= 14220791;
srom_1(53219) <= 14619764;
srom_1(53220) <= 14989517;
srom_1(53221) <= 15328316;
srom_1(53222) <= 15634573;
srom_1(53223) <= 15906851;
srom_1(53224) <= 16143873;
srom_1(53225) <= 16344528;
srom_1(53226) <= 16507875;
srom_1(53227) <= 16633148;
srom_1(53228) <= 16719759;
srom_1(53229) <= 16767303;
srom_1(53230) <= 16775556;
srom_1(53231) <= 16744480;
srom_1(53232) <= 16674220;
srom_1(53233) <= 16565107;
srom_1(53234) <= 16417651;
srom_1(53235) <= 16232544;
srom_1(53236) <= 16010654;
srom_1(53237) <= 15753021;
srom_1(53238) <= 15460854;
srom_1(53239) <= 15135524;
srom_1(53240) <= 14778554;
srom_1(53241) <= 14391620;
srom_1(53242) <= 13976536;
srom_1(53243) <= 13535248;
srom_1(53244) <= 13069825;
srom_1(53245) <= 12582451;
srom_1(53246) <= 12075410;
srom_1(53247) <= 11551081;
srom_1(53248) <= 11011922;
srom_1(53249) <= 10460461;
srom_1(53250) <= 9899284;
srom_1(53251) <= 9331024;
srom_1(53252) <= 8758344;
srom_1(53253) <= 8183930;
srom_1(53254) <= 7610476;
srom_1(53255) <= 7040671;
srom_1(53256) <= 6477187;
srom_1(53257) <= 5922666;
srom_1(53258) <= 5379709;
srom_1(53259) <= 4850861;
srom_1(53260) <= 4338604;
srom_1(53261) <= 3845338;
srom_1(53262) <= 3373377;
srom_1(53263) <= 2924934;
srom_1(53264) <= 2502112;
srom_1(53265) <= 2106895;
srom_1(53266) <= 1741134;
srom_1(53267) <= 1406545;
srom_1(53268) <= 1104698;
srom_1(53269) <= 837007;
srom_1(53270) <= 604729;
srom_1(53271) <= 408952;
srom_1(53272) <= 250594;
srom_1(53273) <= 130398;
srom_1(53274) <= 48928;
srom_1(53275) <= 6565;
srom_1(53276) <= 3509;
srom_1(53277) <= 39773;
srom_1(53278) <= 115187;
srom_1(53279) <= 229399;
srom_1(53280) <= 381872;
srom_1(53281) <= 571891;
srom_1(53282) <= 798566;
srom_1(53283) <= 1060833;
srom_1(53284) <= 1357462;
srom_1(53285) <= 1687063;
srom_1(53286) <= 2048089;
srom_1(53287) <= 2438849;
srom_1(53288) <= 2857509;
srom_1(53289) <= 3302106;
srom_1(53290) <= 3770555;
srom_1(53291) <= 4260660;
srom_1(53292) <= 4770123;
srom_1(53293) <= 5296554;
srom_1(53294) <= 5837484;
srom_1(53295) <= 6390378;
srom_1(53296) <= 6952642;
srom_1(53297) <= 7521639;
srom_1(53298) <= 8094702;
srom_1(53299) <= 8669144;
srom_1(53300) <= 9242270;
srom_1(53301) <= 9811392;
srom_1(53302) <= 10373843;
srom_1(53303) <= 10926985;
srom_1(53304) <= 11468223;
srom_1(53305) <= 11995019;
srom_1(53306) <= 12504904;
srom_1(53307) <= 12995487;
srom_1(53308) <= 13464465;
srom_1(53309) <= 13909642;
srom_1(53310) <= 14328928;
srom_1(53311) <= 14720359;
srom_1(53312) <= 15082097;
srom_1(53313) <= 15412448;
srom_1(53314) <= 15709861;
srom_1(53315) <= 15972942;
srom_1(53316) <= 16200458;
srom_1(53317) <= 16391341;
srom_1(53318) <= 16544697;
srom_1(53319) <= 16659806;
srom_1(53320) <= 16736129;
srom_1(53321) <= 16773307;
srom_1(53322) <= 16771166;
srom_1(53323) <= 16729717;
srom_1(53324) <= 16649154;
srom_1(53325) <= 16529853;
srom_1(53326) <= 16372376;
srom_1(53327) <= 16177460;
srom_1(53328) <= 15946020;
srom_1(53329) <= 15679140;
srom_1(53330) <= 15378072;
srom_1(53331) <= 15044229;
srom_1(53332) <= 14679174;
srom_1(53333) <= 14284622;
srom_1(53334) <= 13862420;
srom_1(53335) <= 13414551;
srom_1(53336) <= 12943112;
srom_1(53337) <= 12450317;
srom_1(53338) <= 11938474;
srom_1(53339) <= 11409985;
srom_1(53340) <= 10867327;
srom_1(53341) <= 10313047;
srom_1(53342) <= 9749741;
srom_1(53343) <= 9180053;
srom_1(53344) <= 8606653;
srom_1(53345) <= 8032231;
srom_1(53346) <= 7459481;
srom_1(53347) <= 6891087;
srom_1(53348) <= 6329715;
srom_1(53349) <= 5777998;
srom_1(53350) <= 5238524;
srom_1(53351) <= 4713821;
srom_1(53352) <= 4206351;
srom_1(53353) <= 3718492;
srom_1(53354) <= 3252534;
srom_1(53355) <= 2810660;
srom_1(53356) <= 2394943;
srom_1(53357) <= 2007332;
srom_1(53358) <= 1649646;
srom_1(53359) <= 1323560;
srom_1(53360) <= 1030605;
srom_1(53361) <= 772155;
srom_1(53362) <= 549420;
srom_1(53363) <= 363446;
srom_1(53364) <= 215105;
srom_1(53365) <= 105092;
srom_1(53366) <= 33924;
srom_1(53367) <= 1933;
srom_1(53368) <= 9271;
srom_1(53369) <= 55902;
srom_1(53370) <= 141608;
srom_1(53371) <= 265987;
srom_1(53372) <= 428455;
srom_1(53373) <= 628252;
srom_1(53374) <= 864439;
srom_1(53375) <= 1135910;
srom_1(53376) <= 1441392;
srom_1(53377) <= 1779451;
srom_1(53378) <= 2148503;
srom_1(53379) <= 2546817;
srom_1(53380) <= 2972524;
srom_1(53381) <= 3423630;
srom_1(53382) <= 3898019;
srom_1(53383) <= 4393465;
srom_1(53384) <= 4907646;
srom_1(53385) <= 5438150;
srom_1(53386) <= 5982490;
srom_1(53387) <= 6538113;
srom_1(53388) <= 7102414;
srom_1(53389) <= 7672746;
srom_1(53390) <= 8246435;
srom_1(53391) <= 8820790;
srom_1(53392) <= 9393119;
srom_1(53393) <= 9960738;
srom_1(53394) <= 10520984;
srom_1(53395) <= 11071231;
srom_1(53396) <= 11608898;
srom_1(53397) <= 12131464;
srom_1(53398) <= 12636478;
srom_1(53399) <= 13121573;
srom_1(53400) <= 13584473;
srom_1(53401) <= 14023008;
srom_1(53402) <= 14435121;
srom_1(53403) <= 14818881;
srom_1(53404) <= 15172486;
srom_1(53405) <= 15494279;
srom_1(53406) <= 15782752;
srom_1(53407) <= 16036551;
srom_1(53408) <= 16254486;
srom_1(53409) <= 16435535;
srom_1(53410) <= 16578849;
srom_1(53411) <= 16683757;
srom_1(53412) <= 16749766;
srom_1(53413) <= 16776566;
srom_1(53414) <= 16764032;
srom_1(53415) <= 16712223;
srom_1(53416) <= 16621382;
srom_1(53417) <= 16491935;
srom_1(53418) <= 16324488;
srom_1(53419) <= 16119827;
srom_1(53420) <= 15878912;
srom_1(53421) <= 15602872;
srom_1(53422) <= 15293002;
srom_1(53423) <= 14950755;
srom_1(53424) <= 14577735;
srom_1(53425) <= 14175693;
srom_1(53426) <= 13746513;
srom_1(53427) <= 13292208;
srom_1(53428) <= 12814909;
srom_1(53429) <= 12316853;
srom_1(53430) <= 11800376;
srom_1(53431) <= 11267900;
srom_1(53432) <= 10721922;
srom_1(53433) <= 10165002;
srom_1(53434) <= 9599753;
srom_1(53435) <= 9028823;
srom_1(53436) <= 8454892;
srom_1(53437) <= 7880650;
srom_1(53438) <= 7308789;
srom_1(53439) <= 6741993;
srom_1(53440) <= 6182918;
srom_1(53441) <= 5634186;
srom_1(53442) <= 5098370;
srom_1(53443) <= 4577984;
srom_1(53444) <= 4075467;
srom_1(53445) <= 3593175;
srom_1(53446) <= 3133372;
srom_1(53447) <= 2698211;
srom_1(53448) <= 2289735;
srom_1(53449) <= 1909859;
srom_1(53450) <= 1560364;
srom_1(53451) <= 1242888;
srom_1(53452) <= 958922;
srom_1(53453) <= 709796;
srom_1(53454) <= 496678;
srom_1(53455) <= 320568;
srom_1(53456) <= 182292;
srom_1(53457) <= 82499;
srom_1(53458) <= 21655;
srom_1(53459) <= 47;
srom_1(53460) <= 17776;
srom_1(53461) <= 74759;
srom_1(53462) <= 170728;
srom_1(53463) <= 305233;
srom_1(53464) <= 477645;
srom_1(53465) <= 687153;
srom_1(53466) <= 932776;
srom_1(53467) <= 1213363;
srom_1(53468) <= 1527596;
srom_1(53469) <= 1874003;
srom_1(53470) <= 2250959;
srom_1(53471) <= 2656697;
srom_1(53472) <= 3089314;
srom_1(53473) <= 3546780;
srom_1(53474) <= 4026952;
srom_1(53475) <= 4527577;
srom_1(53476) <= 5046308;
srom_1(53477) <= 5580712;
srom_1(53478) <= 6128283;
srom_1(53479) <= 6686454;
srom_1(53480) <= 7252607;
srom_1(53481) <= 7824086;
srom_1(53482) <= 8398213;
srom_1(53483) <= 8972295;
srom_1(53484) <= 9543640;
srom_1(53485) <= 10109568;
srom_1(53486) <= 10667426;
srom_1(53487) <= 11214598;
srom_1(53488) <= 11748518;
srom_1(53489) <= 12266683;
srom_1(53490) <= 12766661;
srom_1(53491) <= 13246110;
srom_1(53492) <= 13702780;
srom_1(53493) <= 14134529;
srom_1(53494) <= 14539335;
srom_1(53495) <= 14915297;
srom_1(53496) <= 15260654;
srom_1(53497) <= 15573785;
srom_1(53498) <= 15853222;
srom_1(53499) <= 16097655;
srom_1(53500) <= 16305938;
srom_1(53501) <= 16477094;
srom_1(53502) <= 16610320;
srom_1(53503) <= 16704992;
srom_1(53504) <= 16760665;
srom_1(53505) <= 16777079;
srom_1(53506) <= 16754156;
srom_1(53507) <= 16692004;
srom_1(53508) <= 16590915;
srom_1(53509) <= 16451363;
srom_1(53510) <= 16274001;
srom_1(53511) <= 16059662;
srom_1(53512) <= 15809351;
srom_1(53513) <= 15524242;
srom_1(53514) <= 15205671;
srom_1(53515) <= 14855132;
srom_1(53516) <= 14474270;
srom_1(53517) <= 14064870;
srom_1(53518) <= 13628852;
srom_1(53519) <= 13168261;
srom_1(53520) <= 12685256;
srom_1(53521) <= 12182103;
srom_1(53522) <= 11661160;
srom_1(53523) <= 11124872;
srom_1(53524) <= 10575752;
srom_1(53525) <= 10016377;
srom_1(53526) <= 9449367;
srom_1(53527) <= 8877384;
srom_1(53528) <= 8303109;
srom_1(53529) <= 7729234;
srom_1(53530) <= 7158452;
srom_1(53531) <= 6593438;
srom_1(53532) <= 6036842;
srom_1(53533) <= 5491275;
srom_1(53534) <= 4959294;
srom_1(53535) <= 4443394;
srom_1(53536) <= 3945995;
srom_1(53537) <= 3469429;
srom_1(53538) <= 3015930;
srom_1(53539) <= 2587626;
srom_1(53540) <= 2186525;
srom_1(53541) <= 1814507;
srom_1(53542) <= 1473317;
srom_1(53543) <= 1164556;
srom_1(53544) <= 889671;
srom_1(53545) <= 649950;
srom_1(53546) <= 446519;
srom_1(53547) <= 280332;
srom_1(53548) <= 152166;
srom_1(53549) <= 62624;
srom_1(53550) <= 12126;
srom_1(53551) <= 908;
srom_1(53552) <= 29022;
srom_1(53553) <= 96338;
srom_1(53554) <= 202539;
srom_1(53555) <= 347127;
srom_1(53556) <= 529424;
srom_1(53557) <= 748576;
srom_1(53558) <= 1003554;
srom_1(53559) <= 1293164;
srom_1(53560) <= 1616046;
srom_1(53561) <= 1970688;
srom_1(53562) <= 2355425;
srom_1(53563) <= 2768454;
srom_1(53564) <= 3207838;
srom_1(53565) <= 3671516;
srom_1(53566) <= 4157314;
srom_1(53567) <= 4662954;
srom_1(53568) <= 5186065;
srom_1(53569) <= 5724194;
srom_1(53570) <= 6274817;
srom_1(53571) <= 6835352;
srom_1(53572) <= 7403171;
srom_1(53573) <= 7975612;
srom_1(53574) <= 8549989;
srom_1(53575) <= 9123609;
srom_1(53576) <= 9693782;
srom_1(53577) <= 10257835;
srom_1(53578) <= 10813123;
srom_1(53579) <= 11357041;
srom_1(53580) <= 11887039;
srom_1(53581) <= 12400632;
srom_1(53582) <= 12895411;
srom_1(53583) <= 13369056;
srom_1(53584) <= 13819346;
srom_1(53585) <= 14244170;
srom_1(53586) <= 14641534;
srom_1(53587) <= 15009577;
srom_1(53588) <= 15346572;
srom_1(53589) <= 15650938;
srom_1(53590) <= 15921249;
srom_1(53591) <= 16156236;
srom_1(53592) <= 16354799;
srom_1(53593) <= 16516005;
srom_1(53594) <= 16639099;
srom_1(53595) <= 16723504;
srom_1(53596) <= 16768823;
srom_1(53597) <= 16774845;
srom_1(53598) <= 16741541;
srom_1(53599) <= 16669067;
srom_1(53600) <= 16557763;
srom_1(53601) <= 16408151;
srom_1(53602) <= 16220933;
srom_1(53603) <= 15996986;
srom_1(53604) <= 15737361;
srom_1(53605) <= 15443276;
srom_1(53606) <= 15116108;
srom_1(53607) <= 14757393;
srom_1(53608) <= 14368812;
srom_1(53609) <= 13952188;
srom_1(53610) <= 13509475;
srom_1(53611) <= 13042748;
srom_1(53612) <= 12554196;
srom_1(53613) <= 12046111;
srom_1(53614) <= 11520874;
srom_1(53615) <= 10980948;
srom_1(53616) <= 10428867;
srom_1(53617) <= 9867218;
srom_1(53618) <= 9298635;
srom_1(53619) <= 8725785;
srom_1(53620) <= 8151353;
srom_1(53621) <= 7578035;
srom_1(53622) <= 7008517;
srom_1(53623) <= 6445471;
srom_1(53624) <= 5891537;
srom_1(53625) <= 5349312;
srom_1(53626) <= 4821340;
srom_1(53627) <= 4310096;
srom_1(53628) <= 3817978;
srom_1(53629) <= 3347293;
srom_1(53630) <= 2900248;
srom_1(53631) <= 2478940;
srom_1(53632) <= 2085344;
srom_1(53633) <= 1721307;
srom_1(53634) <= 1388535;
srom_1(53635) <= 1088589;
srom_1(53636) <= 822875;
srom_1(53637) <= 592639;
srom_1(53638) <= 398961;
srom_1(53639) <= 242750;
srom_1(53640) <= 124737;
srom_1(53641) <= 45476;
srom_1(53642) <= 5339;
srom_1(53643) <= 4514;
srom_1(53644) <= 43005;
srom_1(53645) <= 120632;
srom_1(53646) <= 237029;
srom_1(53647) <= 391653;
srom_1(53648) <= 583777;
srom_1(53649) <= 812500;
srom_1(53650) <= 1076750;
srom_1(53651) <= 1375288;
srom_1(53652) <= 1706714;
srom_1(53653) <= 2069474;
srom_1(53654) <= 2461866;
srom_1(53655) <= 2882051;
srom_1(53656) <= 3328058;
srom_1(53657) <= 3797795;
srom_1(53658) <= 4289061;
srom_1(53659) <= 4799550;
srom_1(53660) <= 5326870;
srom_1(53661) <= 5868548;
srom_1(53662) <= 6422042;
srom_1(53663) <= 6984759;
srom_1(53664) <= 7554059;
srom_1(53665) <= 8127272;
srom_1(53666) <= 8701711;
srom_1(53667) <= 9274682;
srom_1(53668) <= 9843497;
srom_1(53669) <= 10405490;
srom_1(53670) <= 10958025;
srom_1(53671) <= 11498512;
srom_1(53672) <= 12024415;
srom_1(53673) <= 12533268;
srom_1(53674) <= 13022685;
srom_1(53675) <= 13490372;
srom_1(53676) <= 13934135;
srom_1(53677) <= 14351893;
srom_1(53678) <= 14741687;
srom_1(53679) <= 15101689;
srom_1(53680) <= 15430212;
srom_1(53681) <= 15725713;
srom_1(53682) <= 15986809;
srom_1(53683) <= 16212274;
srom_1(53684) <= 16401051;
srom_1(53685) <= 16552255;
srom_1(53686) <= 16665177;
srom_1(53687) <= 16739287;
srom_1(53688) <= 16774238;
srom_1(53689) <= 16769866;
srom_1(53690) <= 16726191;
srom_1(53691) <= 16643419;
srom_1(53692) <= 16521937;
srom_1(53693) <= 16362314;
srom_1(53694) <= 16165301;
srom_1(53695) <= 15931820;
srom_1(53696) <= 15662966;
srom_1(53697) <= 15360000;
srom_1(53698) <= 15024343;
srom_1(53699) <= 14657568;
srom_1(53700) <= 14261397;
srom_1(53701) <= 13837685;
srom_1(53702) <= 13388422;
srom_1(53703) <= 12915712;
srom_1(53704) <= 12421773;
srom_1(53705) <= 11908921;
srom_1(53706) <= 11379562;
srom_1(53707) <= 10836176;
srom_1(53708) <= 10281313;
srom_1(53709) <= 9717575;
srom_1(53710) <= 9147605;
srom_1(53711) <= 8574075;
srom_1(53712) <= 7999676;
srom_1(53713) <= 7427100;
srom_1(53714) <= 6859034;
srom_1(53715) <= 6298140;
srom_1(53716) <= 5747049;
srom_1(53717) <= 5208345;
srom_1(53718) <= 4684554;
srom_1(53719) <= 4178133;
srom_1(53720) <= 3691457;
srom_1(53721) <= 3226807;
srom_1(53722) <= 2786362;
srom_1(53723) <= 2372188;
srom_1(53724) <= 1986228;
srom_1(53725) <= 1630290;
srom_1(53726) <= 1306044;
srom_1(53727) <= 1015011;
srom_1(53728) <= 758556;
srom_1(53729) <= 537880;
srom_1(53730) <= 354019;
srom_1(53731) <= 207834;
srom_1(53732) <= 100013;
srom_1(53733) <= 31059;
srom_1(53734) <= 1297;
srom_1(53735) <= 10866;
srom_1(53736) <= 59721;
srom_1(53737) <= 147632;
srom_1(53738) <= 274189;
srom_1(53739) <= 438797;
srom_1(53740) <= 640684;
srom_1(53741) <= 878904;
srom_1(53742) <= 1152340;
srom_1(53743) <= 1459709;
srom_1(53744) <= 1799570;
srom_1(53745) <= 2170329;
srom_1(53746) <= 2570247;
srom_1(53747) <= 2997451;
srom_1(53748) <= 3449935;
srom_1(53749) <= 3925578;
srom_1(53750) <= 4422150;
srom_1(53751) <= 4937321;
srom_1(53752) <= 5468678;
srom_1(53753) <= 6013726;
srom_1(53754) <= 6569912;
srom_1(53755) <= 7134626;
srom_1(53756) <= 7705220;
srom_1(53757) <= 8279019;
srom_1(53758) <= 8853331;
srom_1(53759) <= 9425465;
srom_1(53760) <= 9992736;
srom_1(53761) <= 10552485;
srom_1(53762) <= 11102087;
srom_1(53763) <= 11638964;
srom_1(53764) <= 12160600;
srom_1(53765) <= 12664547;
srom_1(53766) <= 13148443;
srom_1(53767) <= 13610018;
srom_1(53768) <= 14047108;
srom_1(53769) <= 14457664;
srom_1(53770) <= 14839759;
srom_1(53771) <= 15191604;
srom_1(53772) <= 15511546;
srom_1(53773) <= 15798087;
srom_1(53774) <= 16049882;
srom_1(53775) <= 16265750;
srom_1(53776) <= 16444680;
srom_1(53777) <= 16585832;
srom_1(53778) <= 16688545;
srom_1(53779) <= 16752337;
srom_1(53780) <= 16776908;
srom_1(53781) <= 16762143;
srom_1(53782) <= 16708112;
srom_1(53783) <= 16615068;
srom_1(53784) <= 16483447;
srom_1(53785) <= 16313867;
srom_1(53786) <= 16107122;
srom_1(53787) <= 15864183;
srom_1(53788) <= 15586188;
srom_1(53789) <= 15274442;
srom_1(53790) <= 14930405;
srom_1(53791) <= 14555691;
srom_1(53792) <= 14152058;
srom_1(53793) <= 13721398;
srom_1(53794) <= 13265731;
srom_1(53795) <= 12787193;
srom_1(53796) <= 12288029;
srom_1(53797) <= 11770579;
srom_1(53798) <= 11237270;
srom_1(53799) <= 10690603;
srom_1(53800) <= 10133140;
srom_1(53801) <= 9567497;
srom_1(53802) <= 8996326;
srom_1(53803) <= 8422305;
srom_1(53804) <= 7848125;
srom_1(53805) <= 7276481;
srom_1(53806) <= 6710051;
srom_1(53807) <= 6151493;
srom_1(53808) <= 5603426;
srom_1(53809) <= 5068419;
srom_1(53810) <= 4548981;
srom_1(53811) <= 4047549;
srom_1(53812) <= 3566474;
srom_1(53813) <= 3108011;
srom_1(53814) <= 2674311;
srom_1(53815) <= 2267407;
srom_1(53816) <= 1889207;
srom_1(53817) <= 1541486;
srom_1(53818) <= 1225873;
srom_1(53819) <= 943848;
srom_1(53820) <= 696734;
srom_1(53821) <= 485691;
srom_1(53822) <= 311706;
srom_1(53823) <= 175598;
srom_1(53824) <= 78002;
srom_1(53825) <= 19378;
srom_1(53826) <= 1;
srom_1(53827) <= 19960;
srom_1(53828) <= 79163;
srom_1(53829) <= 177331;
srom_1(53830) <= 314005;
srom_1(53831) <= 488544;
srom_1(53832) <= 700129;
srom_1(53833) <= 947767;
srom_1(53834) <= 1230299;
srom_1(53835) <= 1546398;
srom_1(53836) <= 1894582;
srom_1(53837) <= 2273219;
srom_1(53838) <= 2680534;
srom_1(53839) <= 3114615;
srom_1(53840) <= 3573428;
srom_1(53841) <= 4054821;
srom_1(53842) <= 4556537;
srom_1(53843) <= 5076223;
srom_1(53844) <= 5611441;
srom_1(53845) <= 6159683;
srom_1(53846) <= 6718377;
srom_1(53847) <= 7284903;
srom_1(53848) <= 7856604;
srom_1(53849) <= 8430801;
srom_1(53850) <= 9004799;
srom_1(53851) <= 9575908;
srom_1(53852) <= 10141450;
srom_1(53853) <= 10698771;
srom_1(53854) <= 11245260;
srom_1(53855) <= 11778353;
srom_1(53856) <= 12295550;
srom_1(53857) <= 12794426;
srom_1(53858) <= 13272641;
srom_1(53859) <= 13727954;
srom_1(53860) <= 14158229;
srom_1(53861) <= 14561448;
srom_1(53862) <= 14935720;
srom_1(53863) <= 15279291;
srom_1(53864) <= 15590549;
srom_1(53865) <= 15868034;
srom_1(53866) <= 16110446;
srom_1(53867) <= 16316648;
srom_1(53868) <= 16485672;
srom_1(53869) <= 16616726;
srom_1(53870) <= 16709196;
srom_1(53871) <= 16762648;
srom_1(53872) <= 16776831;
srom_1(53873) <= 16751678;
srom_1(53874) <= 16687309;
srom_1(53875) <= 16584024;
srom_1(53876) <= 16442308;
srom_1(53877) <= 16262825;
srom_1(53878) <= 16046417;
srom_1(53879) <= 15794099;
srom_1(53880) <= 15507055;
srom_1(53881) <= 15186629;
srom_1(53882) <= 14834325;
srom_1(53883) <= 14451795;
srom_1(53884) <= 14040833;
srom_1(53885) <= 13603365;
srom_1(53886) <= 13141444;
srom_1(53887) <= 12657235;
srom_1(53888) <= 12153009;
srom_1(53889) <= 11631130;
srom_1(53890) <= 11094046;
srom_1(53891) <= 10544275;
srom_1(53892) <= 9984396;
srom_1(53893) <= 9417033;
srom_1(53894) <= 8844848;
srom_1(53895) <= 8270523;
srom_1(53896) <= 7696752;
srom_1(53897) <= 7126226;
srom_1(53898) <= 6561619;
srom_1(53899) <= 6005579;
srom_1(53900) <= 5460714;
srom_1(53901) <= 4929579;
srom_1(53902) <= 4414665;
srom_1(53903) <= 3918386;
srom_1(53904) <= 3443069;
srom_1(53905) <= 2990944;
srom_1(53906) <= 2564130;
srom_1(53907) <= 2164629;
srom_1(53908) <= 1794315;
srom_1(53909) <= 1454923;
srom_1(53910) <= 1148046;
srom_1(53911) <= 875122;
srom_1(53912) <= 637432;
srom_1(53913) <= 436089;
srom_1(53914) <= 272039;
srom_1(53915) <= 146050;
srom_1(53916) <= 58713;
srom_1(53917) <= 10438;
srom_1(53918) <= 1451;
srom_1(53919) <= 31794;
srom_1(53920) <= 101325;
srom_1(53921) <= 209718;
srom_1(53922) <= 356465;
srom_1(53923) <= 540877;
srom_1(53924) <= 762090;
srom_1(53925) <= 1019066;
srom_1(53926) <= 1310601;
srom_1(53927) <= 1635327;
srom_1(53928) <= 1991721;
srom_1(53929) <= 2378112;
srom_1(53930) <= 2792689;
srom_1(53931) <= 3233507;
srom_1(53932) <= 3698499;
srom_1(53933) <= 4185484;
srom_1(53934) <= 4692179;
srom_1(53935) <= 5216208;
srom_1(53936) <= 5755114;
srom_1(53937) <= 6306369;
srom_1(53938) <= 6867388;
srom_1(53939) <= 7435541;
srom_1(53940) <= 8008163;
srom_1(53941) <= 8582569;
srom_1(53942) <= 9156066;
srom_1(53943) <= 9725963;
srom_1(53944) <= 10289590;
srom_1(53945) <= 10844301;
srom_1(53946) <= 11387498;
srom_1(53947) <= 11916631;
srom_1(53948) <= 12429221;
srom_1(53949) <= 12922862;
srom_1(53950) <= 13395241;
srom_1(53951) <= 13844142;
srom_1(53952) <= 14267460;
srom_1(53953) <= 14663211;
srom_1(53954) <= 15029537;
srom_1(53955) <= 15364722;
srom_1(53956) <= 15667193;
srom_1(53957) <= 15935533;
srom_1(53958) <= 16168482;
srom_1(53959) <= 16364949;
srom_1(53960) <= 16524012;
srom_1(53961) <= 16644926;
srom_1(53962) <= 16727123;
srom_1(53963) <= 16770217;
srom_1(53964) <= 16774008;
srom_1(53965) <= 16738476;
srom_1(53966) <= 16663789;
srom_1(53967) <= 16550296;
srom_1(53968) <= 16398531;
srom_1(53969) <= 16209205;
srom_1(53970) <= 15983205;
srom_1(53971) <= 15721591;
srom_1(53972) <= 15425590;
srom_1(53973) <= 15096591;
srom_1(53974) <= 14736136;
srom_1(53975) <= 14345914;
srom_1(53976) <= 13927757;
srom_1(53977) <= 13483625;
srom_1(53978) <= 13015601;
srom_1(53979) <= 12525879;
srom_1(53980) <= 12016756;
srom_1(53981) <= 11490619;
srom_1(53982) <= 10949936;
srom_1(53983) <= 10397242;
srom_1(53984) <= 9835129;
srom_1(53985) <= 9266233;
srom_1(53986) <= 8693221;
srom_1(53987) <= 8118780;
srom_1(53988) <= 7545605;
srom_1(53989) <= 6976383;
srom_1(53990) <= 6413784;
srom_1(53991) <= 5860445;
srom_1(53992) <= 5318962;
srom_1(53993) <= 4791873;
srom_1(53994) <= 4281650;
srom_1(53995) <= 3790687;
srom_1(53996) <= 3321284;
srom_1(53997) <= 2875644;
srom_1(53998) <= 2455856;
srom_1(53999) <= 2063889;
srom_1(54000) <= 1701581;
srom_1(54001) <= 1370630;
srom_1(54002) <= 1072590;
srom_1(54003) <= 808856;
srom_1(54004) <= 580666;
srom_1(54005) <= 389091;
srom_1(54006) <= 235028;
srom_1(54007) <= 119200;
srom_1(54008) <= 42150;
srom_1(54009) <= 4240;
srom_1(54010) <= 5647;
srom_1(54011) <= 46364;
srom_1(54012) <= 126201;
srom_1(54013) <= 244783;
srom_1(54014) <= 401554;
srom_1(54015) <= 595780;
srom_1(54016) <= 826548;
srom_1(54017) <= 1092778;
srom_1(54018) <= 1393220;
srom_1(54019) <= 1726467;
srom_1(54020) <= 2090954;
srom_1(54021) <= 2484973;
srom_1(54022) <= 2906676;
srom_1(54023) <= 3354086;
srom_1(54024) <= 3825104;
srom_1(54025) <= 4317523;
srom_1(54026) <= 4829032;
srom_1(54027) <= 5357233;
srom_1(54028) <= 5899649;
srom_1(54029) <= 6453737;
srom_1(54030) <= 7016898;
srom_1(54031) <= 7586491;
srom_1(54032) <= 8159846;
srom_1(54033) <= 8734274;
srom_1(54034) <= 9307081;
srom_1(54035) <= 9875580;
srom_1(54036) <= 10437107;
srom_1(54037) <= 10989028;
srom_1(54038) <= 11528754;
srom_1(54039) <= 12053755;
srom_1(54040) <= 12561569;
srom_1(54041) <= 13049814;
srom_1(54042) <= 13516202;
srom_1(54043) <= 13958544;
srom_1(54044) <= 14374767;
srom_1(54045) <= 14762919;
srom_1(54046) <= 15121180;
srom_1(54047) <= 15447869;
srom_1(54048) <= 15741455;
srom_1(54049) <= 16000561;
srom_1(54050) <= 16223972;
srom_1(54051) <= 16410640;
srom_1(54052) <= 16559690;
srom_1(54053) <= 16670423;
srom_1(54054) <= 16742319;
srom_1(54055) <= 16775043;
srom_1(54056) <= 16768439;
srom_1(54057) <= 16722540;
srom_1(54058) <= 16637559;
srom_1(54059) <= 16513897;
srom_1(54060) <= 16352132;
srom_1(54061) <= 16153024;
srom_1(54062) <= 15917506;
srom_1(54063) <= 15646682;
srom_1(54064) <= 15341822;
srom_1(54065) <= 15004357;
srom_1(54066) <= 14635868;
srom_1(54067) <= 14238083;
srom_1(54068) <= 13812868;
srom_1(54069) <= 13362217;
srom_1(54070) <= 12888243;
srom_1(54071) <= 12393168;
srom_1(54072) <= 11879315;
srom_1(54073) <= 11349093;
srom_1(54074) <= 10804988;
srom_1(54075) <= 10249552;
srom_1(54076) <= 9685389;
srom_1(54077) <= 9115145;
srom_1(54078) <= 8541494;
srom_1(54079) <= 7967126;
srom_1(54080) <= 7394735;
srom_1(54081) <= 6827004;
srom_1(54082) <= 6266596;
srom_1(54083) <= 5716139;
srom_1(54084) <= 5178214;
srom_1(54085) <= 4655343;
srom_1(54086) <= 4149980;
srom_1(54087) <= 3664492;
srom_1(54088) <= 3201158;
srom_1(54089) <= 2762149;
srom_1(54090) <= 2349525;
srom_1(54091) <= 1965220;
srom_1(54092) <= 1611037;
srom_1(54093) <= 1288635;
srom_1(54094) <= 999528;
srom_1(54095) <= 745071;
srom_1(54096) <= 526458;
srom_1(54097) <= 344712;
srom_1(54098) <= 200687;
srom_1(54099) <= 95058;
srom_1(54100) <= 28320;
srom_1(54101) <= 787;
srom_1(54102) <= 12587;
srom_1(54103) <= 63665;
srom_1(54104) <= 153781;
srom_1(54105) <= 282514;
srom_1(54106) <= 449259;
srom_1(54107) <= 653234;
srom_1(54108) <= 893482;
srom_1(54109) <= 1168878;
srom_1(54110) <= 1478130;
srom_1(54111) <= 1819788;
srom_1(54112) <= 2192248;
srom_1(54113) <= 2593766;
srom_1(54114) <= 3022458;
srom_1(54115) <= 3476313;
srom_1(54116) <= 3953204;
srom_1(54117) <= 4450894;
srom_1(54118) <= 4967049;
srom_1(54119) <= 5499250;
srom_1(54120) <= 6044999;
srom_1(54121) <= 6601738;
srom_1(54122) <= 7166857;
srom_1(54123) <= 7737704;
srom_1(54124) <= 8311604;
srom_1(54125) <= 8885866;
srom_1(54126) <= 9457795;
srom_1(54127) <= 10024710;
srom_1(54128) <= 10583954;
srom_1(54129) <= 11132902;
srom_1(54130) <= 11668982;
srom_1(54131) <= 12189679;
srom_1(54132) <= 12692551;
srom_1(54133) <= 13175240;
srom_1(54134) <= 13635484;
srom_1(54135) <= 14071123;
srom_1(54136) <= 14480114;
srom_1(54137) <= 14860541;
srom_1(54138) <= 15210618;
srom_1(54139) <= 15528705;
srom_1(54140) <= 15813309;
srom_1(54141) <= 16063097;
srom_1(54142) <= 16276896;
srom_1(54143) <= 16453704;
srom_1(54144) <= 16592692;
srom_1(54145) <= 16693208;
srom_1(54146) <= 16754781;
srom_1(54147) <= 16777123;
srom_1(54148) <= 16760127;
srom_1(54149) <= 16703875;
srom_1(54150) <= 16608630;
srom_1(54151) <= 16474838;
srom_1(54152) <= 16303127;
srom_1(54153) <= 16094302;
srom_1(54154) <= 15849342;
srom_1(54155) <= 15569396;
srom_1(54156) <= 15255778;
srom_1(54157) <= 14909956;
srom_1(54158) <= 14533554;
srom_1(54159) <= 14128336;
srom_1(54160) <= 13696203;
srom_1(54161) <= 13239180;
srom_1(54162) <= 12759412;
srom_1(54163) <= 12259147;
srom_1(54164) <= 11740732;
srom_1(54165) <= 11206597;
srom_1(54166) <= 10659249;
srom_1(54167) <= 10101252;
srom_1(54168) <= 9535224;
srom_1(54169) <= 8963819;
srom_1(54170) <= 8389717;
srom_1(54171) <= 7815610;
srom_1(54172) <= 7244189;
srom_1(54173) <= 6678135;
srom_1(54174) <= 6120102;
srom_1(54175) <= 5572707;
srom_1(54176) <= 5038517;
srom_1(54177) <= 4520037;
srom_1(54178) <= 4019697;
srom_1(54179) <= 3539845;
srom_1(54180) <= 3082730;
srom_1(54181) <= 2650496;
srom_1(54182) <= 2245171;
srom_1(54183) <= 1868654;
srom_1(54184) <= 1522711;
srom_1(54185) <= 1208965;
srom_1(54186) <= 928887;
srom_1(54187) <= 683789;
srom_1(54188) <= 474823;
srom_1(54189) <= 302967;
srom_1(54190) <= 169027;
srom_1(54191) <= 73631;
srom_1(54192) <= 17228;
srom_1(54193) <= 80;
srom_1(54194) <= 22270;
srom_1(54195) <= 83692;
srom_1(54196) <= 184058;
srom_1(54197) <= 322899;
srom_1(54198) <= 499562;
srom_1(54199) <= 713220;
srom_1(54200) <= 962870;
srom_1(54201) <= 1247342;
srom_1(54202) <= 1565302;
srom_1(54203) <= 1915259;
srom_1(54204) <= 2295572;
srom_1(54205) <= 2704457;
srom_1(54206) <= 3139997;
srom_1(54207) <= 3600149;
srom_1(54208) <= 4082756;
srom_1(54209) <= 4585555;
srom_1(54210) <= 5106187;
srom_1(54211) <= 5642212;
srom_1(54212) <= 6191116;
srom_1(54213) <= 6750324;
srom_1(54214) <= 7317215;
srom_1(54215) <= 7889131;
srom_1(54216) <= 8463388;
srom_1(54217) <= 9037294;
srom_1(54218) <= 9608159;
srom_1(54219) <= 10173305;
srom_1(54220) <= 10730082;
srom_1(54221) <= 11275878;
srom_1(54222) <= 11808136;
srom_1(54223) <= 12324358;
srom_1(54224) <= 12822124;
srom_1(54225) <= 13299099;
srom_1(54226) <= 13753048;
srom_1(54227) <= 14181841;
srom_1(54228) <= 14583467;
srom_1(54229) <= 14956044;
srom_1(54230) <= 15297824;
srom_1(54231) <= 15607204;
srom_1(54232) <= 15882733;
srom_1(54233) <= 16123120;
srom_1(54234) <= 16327237;
srom_1(54235) <= 16494127;
srom_1(54236) <= 16623008;
srom_1(54237) <= 16713275;
srom_1(54238) <= 16764504;
srom_1(54239) <= 16776456;
srom_1(54240) <= 16749075;
srom_1(54241) <= 16682488;
srom_1(54242) <= 16577008;
srom_1(54243) <= 16433131;
srom_1(54244) <= 16251529;
srom_1(54245) <= 16033056;
srom_1(54246) <= 15778736;
srom_1(54247) <= 15489760;
srom_1(54248) <= 15167485;
srom_1(54249) <= 14813421;
srom_1(54250) <= 14429229;
srom_1(54251) <= 14016711;
srom_1(54252) <= 13577800;
srom_1(54253) <= 13114556;
srom_1(54254) <= 12629150;
srom_1(54255) <= 12123858;
srom_1(54256) <= 11601051;
srom_1(54257) <= 11063179;
srom_1(54258) <= 10512766;
srom_1(54259) <= 9952391;
srom_1(54260) <= 9384684;
srom_1(54261) <= 8812305;
srom_1(54262) <= 8237940;
srom_1(54263) <= 7664281;
srom_1(54264) <= 7094018;
srom_1(54265) <= 6529827;
srom_1(54266) <= 5974352;
srom_1(54267) <= 5430198;
srom_1(54268) <= 4899917;
srom_1(54269) <= 4385996;
srom_1(54270) <= 3890845;
srom_1(54271) <= 3416785;
srom_1(54272) <= 2966039;
srom_1(54273) <= 2540722;
srom_1(54274) <= 2142828;
srom_1(54275) <= 1774222;
srom_1(54276) <= 1436633;
srom_1(54277) <= 1131645;
srom_1(54278) <= 860687;
srom_1(54279) <= 625030;
srom_1(54280) <= 425779;
srom_1(54281) <= 263868;
srom_1(54282) <= 140057;
srom_1(54283) <= 54927;
srom_1(54284) <= 8876;
srom_1(54285) <= 2120;
srom_1(54286) <= 34691;
srom_1(54287) <= 106437;
srom_1(54288) <= 217021;
srom_1(54289) <= 365924;
srom_1(54290) <= 552448;
srom_1(54291) <= 775719;
srom_1(54292) <= 1034689;
srom_1(54293) <= 1328145;
srom_1(54294) <= 1654709;
srom_1(54295) <= 2012850;
srom_1(54296) <= 2400890;
srom_1(54297) <= 2817008;
srom_1(54298) <= 3259254;
srom_1(54299) <= 3725552;
srom_1(54300) <= 4213718;
srom_1(54301) <= 4721461;
srom_1(54302) <= 5246400;
srom_1(54303) <= 5786074;
srom_1(54304) <= 6337953;
srom_1(54305) <= 6899447;
srom_1(54306) <= 7467925;
srom_1(54307) <= 8040720;
srom_1(54308) <= 8615147;
srom_1(54309) <= 9188511;
srom_1(54310) <= 9758124;
srom_1(54311) <= 10321315;
srom_1(54312) <= 10875443;
srom_1(54313) <= 11417909;
srom_1(54314) <= 11946170;
srom_1(54315) <= 12457748;
srom_1(54316) <= 12950245;
srom_1(54317) <= 13421351;
srom_1(54318) <= 13868856;
srom_1(54319) <= 14290662;
srom_1(54320) <= 14684792;
srom_1(54321) <= 15049397;
srom_1(54322) <= 15382767;
srom_1(54323) <= 15683339;
srom_1(54324) <= 15949703;
srom_1(54325) <= 16180611;
srom_1(54326) <= 16374980;
srom_1(54327) <= 16531897;
srom_1(54328) <= 16650628;
srom_1(54329) <= 16730616;
srom_1(54330) <= 16771485;
srom_1(54331) <= 16773043;
srom_1(54332) <= 16735285;
srom_1(54333) <= 16658386;
srom_1(54334) <= 16542707;
srom_1(54335) <= 16388790;
srom_1(54336) <= 16197358;
srom_1(54337) <= 15969308;
srom_1(54338) <= 15705710;
srom_1(54339) <= 15407799;
srom_1(54340) <= 15076973;
srom_1(54341) <= 14714782;
srom_1(54342) <= 14322926;
srom_1(54343) <= 13903243;
srom_1(54344) <= 13457699;
srom_1(54345) <= 12988384;
srom_1(54346) <= 12497499;
srom_1(54347) <= 11987347;
srom_1(54348) <= 11460318;
srom_1(54349) <= 10918885;
srom_1(54350) <= 10365587;
srom_1(54351) <= 9803019;
srom_1(54352) <= 9233817;
srom_1(54353) <= 8660652;
srom_1(54354) <= 8086212;
srom_1(54355) <= 7513189;
srom_1(54356) <= 6944271;
srom_1(54357) <= 6382127;
srom_1(54358) <= 5829392;
srom_1(54359) <= 5288657;
srom_1(54360) <= 4762460;
srom_1(54361) <= 4253266;
srom_1(54362) <= 3763465;
srom_1(54363) <= 3295352;
srom_1(54364) <= 2851124;
srom_1(54365) <= 2432862;
srom_1(54366) <= 2042530;
srom_1(54367) <= 1681956;
srom_1(54368) <= 1352832;
srom_1(54369) <= 1056701;
srom_1(54370) <= 794952;
srom_1(54371) <= 568812;
srom_1(54372) <= 379342;
srom_1(54373) <= 227430;
srom_1(54374) <= 113788;
srom_1(54375) <= 38951;
srom_1(54376) <= 3267;
srom_1(54377) <= 6905;
srom_1(54378) <= 49848;
srom_1(54379) <= 131894;
srom_1(54380) <= 252659;
srom_1(54381) <= 411576;
srom_1(54382) <= 607900;
srom_1(54383) <= 840711;
srom_1(54384) <= 1108916;
srom_1(54385) <= 1411258;
srom_1(54386) <= 1746319;
srom_1(54387) <= 2112529;
srom_1(54388) <= 2508169;
srom_1(54389) <= 2931384;
srom_1(54390) <= 3380190;
srom_1(54391) <= 3852482;
srom_1(54392) <= 4346046;
srom_1(54393) <= 4858567;
srom_1(54394) <= 5387641;
srom_1(54395) <= 5930788;
srom_1(54396) <= 6485460;
srom_1(54397) <= 7049057;
srom_1(54398) <= 7618936;
srom_1(54399) <= 8192424;
srom_1(54400) <= 8766831;
srom_1(54401) <= 9339466;
srom_1(54402) <= 9907641;
srom_1(54403) <= 10468693;
srom_1(54404) <= 11019990;
srom_1(54405) <= 11558949;
srom_1(54406) <= 12083040;
srom_1(54407) <= 12589807;
srom_1(54408) <= 13076873;
srom_1(54409) <= 13541954;
srom_1(54410) <= 13982869;
srom_1(54411) <= 14397551;
srom_1(54412) <= 14784055;
srom_1(54413) <= 15140569;
srom_1(54414) <= 15465420;
srom_1(54415) <= 15757086;
srom_1(54416) <= 16014198;
srom_1(54417) <= 16235551;
srom_1(54418) <= 16420107;
srom_1(54419) <= 16567001;
srom_1(54420) <= 16675544;
srom_1(54421) <= 16745226;
srom_1(54422) <= 16775721;
srom_1(54423) <= 16766886;
srom_1(54424) <= 16718762;
srom_1(54425) <= 16631576;
srom_1(54426) <= 16505735;
srom_1(54427) <= 16341830;
srom_1(54428) <= 16140630;
srom_1(54429) <= 15903078;
srom_1(54430) <= 15630288;
srom_1(54431) <= 15323540;
srom_1(54432) <= 14984271;
srom_1(54433) <= 14614073;
srom_1(54434) <= 14214681;
srom_1(54435) <= 13787969;
srom_1(54436) <= 13335937;
srom_1(54437) <= 12860706;
srom_1(54438) <= 12364504;
srom_1(54439) <= 11849657;
srom_1(54440) <= 11318580;
srom_1(54441) <= 10773763;
srom_1(54442) <= 10217762;
srom_1(54443) <= 9653183;
srom_1(54444) <= 9082674;
srom_1(54445) <= 8508910;
srom_1(54446) <= 7934583;
srom_1(54447) <= 7362384;
srom_1(54448) <= 6794997;
srom_1(54449) <= 6235084;
srom_1(54450) <= 5685269;
srom_1(54451) <= 5148131;
srom_1(54452) <= 4626189;
srom_1(54453) <= 4121890;
srom_1(54454) <= 3637599;
srom_1(54455) <= 3175587;
srom_1(54456) <= 2738021;
srom_1(54457) <= 2326953;
srom_1(54458) <= 1944309;
srom_1(54459) <= 1591885;
srom_1(54460) <= 1271334;
srom_1(54461) <= 984157;
srom_1(54462) <= 731703;
srom_1(54463) <= 515154;
srom_1(54464) <= 335527;
srom_1(54465) <= 193663;
srom_1(54466) <= 90229;
srom_1(54467) <= 25708;
srom_1(54468) <= 404;
srom_1(54469) <= 14435;
srom_1(54470) <= 67735;
srom_1(54471) <= 160055;
srom_1(54472) <= 290961;
srom_1(54473) <= 459840;
srom_1(54474) <= 665900;
srom_1(54475) <= 908174;
srom_1(54476) <= 1185526;
srom_1(54477) <= 1496656;
srom_1(54478) <= 1840105;
srom_1(54479) <= 2214262;
srom_1(54480) <= 2617372;
srom_1(54481) <= 3047546;
srom_1(54482) <= 3502766;
srom_1(54483) <= 3980898;
srom_1(54484) <= 4479698;
srom_1(54485) <= 4996829;
srom_1(54486) <= 5529865;
srom_1(54487) <= 6076307;
srom_1(54488) <= 6633591;
srom_1(54489) <= 7199106;
srom_1(54490) <= 7770199;
srom_1(54491) <= 8344191;
srom_1(54492) <= 8918392;
srom_1(54493) <= 9490109;
srom_1(54494) <= 10056660;
srom_1(54495) <= 10615389;
srom_1(54496) <= 11163676;
srom_1(54497) <= 11698950;
srom_1(54498) <= 12218700;
srom_1(54499) <= 12720490;
srom_1(54500) <= 13201966;
srom_1(54501) <= 13660871;
srom_1(54502) <= 14095052;
srom_1(54503) <= 14502473;
srom_1(54504) <= 14881225;
srom_1(54505) <= 15229530;
srom_1(54506) <= 15545756;
srom_1(54507) <= 15828420;
srom_1(54508) <= 16076196;
srom_1(54509) <= 16287922;
srom_1(54510) <= 16462606;
srom_1(54511) <= 16599427;
srom_1(54512) <= 16697746;
srom_1(54513) <= 16757100;
srom_1(54514) <= 16777211;
srom_1(54515) <= 16757985;
srom_1(54516) <= 16699513;
srom_1(54517) <= 16602067;
srom_1(54518) <= 16466106;
srom_1(54519) <= 16292267;
srom_1(54520) <= 16081364;
srom_1(54521) <= 15834388;
srom_1(54522) <= 15552496;
srom_1(54523) <= 15237010;
srom_1(54524) <= 14889410;
srom_1(54525) <= 14511324;
srom_1(54526) <= 14104528;
srom_1(54527) <= 13670927;
srom_1(54528) <= 13212556;
srom_1(54529) <= 12731564;
srom_1(54530) <= 12230206;
srom_1(54531) <= 11710834;
srom_1(54532) <= 11175882;
srom_1(54533) <= 10627860;
srom_1(54534) <= 10069338;
srom_1(54535) <= 9502933;
srom_1(54536) <= 8931304;
srom_1(54537) <= 8357129;
srom_1(54538) <= 7783102;
srom_1(54539) <= 7211915;
srom_1(54540) <= 6646245;
srom_1(54541) <= 6088746;
srom_1(54542) <= 5542032;
srom_1(54543) <= 5008666;
srom_1(54544) <= 4491150;
srom_1(54545) <= 3991911;
srom_1(54546) <= 3513289;
srom_1(54547) <= 3057529;
srom_1(54548) <= 2626769;
srom_1(54549) <= 2223027;
srom_1(54550) <= 1848199;
srom_1(54551) <= 1504040;
srom_1(54552) <= 1192165;
srom_1(54553) <= 914038;
srom_1(54554) <= 670961;
srom_1(54555) <= 464074;
srom_1(54556) <= 294349;
srom_1(54557) <= 162580;
srom_1(54558) <= 69386;
srom_1(54559) <= 15203;
srom_1(54560) <= 287;
srom_1(54561) <= 24706;
srom_1(54562) <= 88346;
srom_1(54563) <= 190909;
srom_1(54564) <= 331914;
srom_1(54565) <= 510699;
srom_1(54566) <= 726427;
srom_1(54567) <= 978085;
srom_1(54568) <= 1264494;
srom_1(54569) <= 1584310;
srom_1(54570) <= 1936034;
srom_1(54571) <= 2318016;
srom_1(54572) <= 2728466;
srom_1(54573) <= 3165457;
srom_1(54574) <= 3626942;
srom_1(54575) <= 4110756;
srom_1(54576) <= 4614630;
srom_1(54577) <= 5136202;
srom_1(54578) <= 5673025;
srom_1(54579) <= 6222582;
srom_1(54580) <= 6782297;
srom_1(54581) <= 7349544;
srom_1(54582) <= 7921664;
srom_1(54583) <= 8495974;
srom_1(54584) <= 9069780;
srom_1(54585) <= 9640391;
srom_1(54586) <= 10205133;
srom_1(54587) <= 10761357;
srom_1(54588) <= 11306453;
srom_1(54589) <= 11837867;
srom_1(54590) <= 12353106;
srom_1(54591) <= 12849755;
srom_1(54592) <= 13325483;
srom_1(54593) <= 13778061;
srom_1(54594) <= 14205366;
srom_1(54595) <= 14605393;
srom_1(54596) <= 14976269;
srom_1(54597) <= 15316252;
srom_1(54598) <= 15623750;
srom_1(54599) <= 15897319;
srom_1(54600) <= 16135677;
srom_1(54601) <= 16337707;
srom_1(54602) <= 16502461;
srom_1(54603) <= 16629166;
srom_1(54604) <= 16717228;
srom_1(54605) <= 16766234;
srom_1(54606) <= 16775955;
srom_1(54607) <= 16746345;
srom_1(54608) <= 16677542;
srom_1(54609) <= 16569870;
srom_1(54610) <= 16423832;
srom_1(54611) <= 16240115;
srom_1(54612) <= 16019580;
srom_1(54613) <= 15763260;
srom_1(54614) <= 15472358;
srom_1(54615) <= 15148238;
srom_1(54616) <= 14792420;
srom_1(54617) <= 14406572;
srom_1(54618) <= 13992504;
srom_1(54619) <= 13552157;
srom_1(54620) <= 13087596;
srom_1(54621) <= 12601000;
srom_1(54622) <= 12094651;
srom_1(54623) <= 11570923;
srom_1(54624) <= 11032272;
srom_1(54625) <= 10481224;
srom_1(54626) <= 9920363;
srom_1(54627) <= 9352319;
srom_1(54628) <= 8779756;
srom_1(54629) <= 8205358;
srom_1(54630) <= 7631820;
srom_1(54631) <= 7061831;
srom_1(54632) <= 6498063;
srom_1(54633) <= 5943161;
srom_1(54634) <= 5399726;
srom_1(54635) <= 4870308;
srom_1(54636) <= 4357387;
srom_1(54637) <= 3863371;
srom_1(54638) <= 3390575;
srom_1(54639) <= 2941216;
srom_1(54640) <= 2517402;
srom_1(54641) <= 2121121;
srom_1(54642) <= 1754229;
srom_1(54643) <= 1418449;
srom_1(54644) <= 1115354;
srom_1(54645) <= 846365;
srom_1(54646) <= 612745;
srom_1(54647) <= 415589;
srom_1(54648) <= 255820;
srom_1(54649) <= 134190;
srom_1(54650) <= 51267;
srom_1(54651) <= 7440;
srom_1(54652) <= 2916;
srom_1(54653) <= 37715;
srom_1(54654) <= 111675;
srom_1(54655) <= 224447;
srom_1(54656) <= 375505;
srom_1(54657) <= 564138;
srom_1(54658) <= 789463;
srom_1(54659) <= 1050423;
srom_1(54660) <= 1345795;
srom_1(54661) <= 1674192;
srom_1(54662) <= 2034076;
srom_1(54663) <= 2423758;
srom_1(54664) <= 2841412;
srom_1(54665) <= 3285078;
srom_1(54666) <= 3752677;
srom_1(54667) <= 4242014;
srom_1(54668) <= 4750797;
srom_1(54669) <= 5276639;
srom_1(54670) <= 5817074;
srom_1(54671) <= 6369567;
srom_1(54672) <= 6931529;
srom_1(54673) <= 7500323;
srom_1(54674) <= 8073282;
srom_1(54675) <= 8647721;
srom_1(54676) <= 9220944;
srom_1(54677) <= 9790264;
srom_1(54678) <= 10353012;
srom_1(54679) <= 10906547;
srom_1(54680) <= 11448275;
srom_1(54681) <= 11975655;
srom_1(54682) <= 12486215;
srom_1(54683) <= 12977559;
srom_1(54684) <= 13447384;
srom_1(54685) <= 13893487;
srom_1(54686) <= 14313775;
srom_1(54687) <= 14706278;
srom_1(54688) <= 15069156;
srom_1(54689) <= 15400706;
srom_1(54690) <= 15699374;
srom_1(54691) <= 15963759;
srom_1(54692) <= 16192622;
srom_1(54693) <= 16384889;
srom_1(54694) <= 16539659;
srom_1(54695) <= 16656206;
srom_1(54696) <= 16733983;
srom_1(54697) <= 16772626;
srom_1(54698) <= 16771953;
srom_1(54699) <= 16731968;
srom_1(54700) <= 16652858;
srom_1(54701) <= 16534994;
srom_1(54702) <= 16378928;
srom_1(54703) <= 16185394;
srom_1(54704) <= 15955297;
srom_1(54705) <= 15689718;
srom_1(54706) <= 15389902;
srom_1(54707) <= 15057253;
srom_1(54708) <= 14693334;
srom_1(54709) <= 14299849;
srom_1(54710) <= 13878645;
srom_1(54711) <= 13431695;
srom_1(54712) <= 12961097;
srom_1(54713) <= 12469057;
srom_1(54714) <= 11957883;
srom_1(54715) <= 11429971;
srom_1(54716) <= 10887796;
srom_1(54717) <= 10333903;
srom_1(54718) <= 9770887;
srom_1(54719) <= 9201389;
srom_1(54720) <= 8628080;
srom_1(54721) <= 8053647;
srom_1(54722) <= 7480786;
srom_1(54723) <= 6912181;
srom_1(54724) <= 6350500;
srom_1(54725) <= 5798377;
srom_1(54726) <= 5258400;
srom_1(54727) <= 4733101;
srom_1(54728) <= 4224944;
srom_1(54729) <= 3736313;
srom_1(54730) <= 3269497;
srom_1(54731) <= 2826687;
srom_1(54732) <= 2409958;
srom_1(54733) <= 2021266;
srom_1(54734) <= 1662432;
srom_1(54735) <= 1335139;
srom_1(54736) <= 1040923;
srom_1(54737) <= 781162;
srom_1(54738) <= 557075;
srom_1(54739) <= 369713;
srom_1(54740) <= 219955;
srom_1(54741) <= 108502;
srom_1(54742) <= 35877;
srom_1(54743) <= 2421;
srom_1(54744) <= 8291;
srom_1(54745) <= 53459;
srom_1(54746) <= 137713;
srom_1(54747) <= 260658;
srom_1(54748) <= 421719;
srom_1(54749) <= 620139;
srom_1(54750) <= 854987;
srom_1(54751) <= 1125164;
srom_1(54752) <= 1429401;
srom_1(54753) <= 1766273;
srom_1(54754) <= 2134198;
srom_1(54755) <= 2531453;
srom_1(54756) <= 2956174;
srom_1(54757) <= 3406370;
srom_1(54758) <= 3879929;
srom_1(54759) <= 4374631;
srom_1(54760) <= 4888155;
srom_1(54761) <= 5418095;
srom_1(54762) <= 5961964;
srom_1(54763) <= 6517213;
srom_1(54764) <= 7081237;
srom_1(54765) <= 7651392;
srom_1(54766) <= 8225004;
srom_1(54767) <= 8799383;
srom_1(54768) <= 9371836;
srom_1(54769) <= 9939678;
srom_1(54770) <= 10500247;
srom_1(54771) <= 11050913;
srom_1(54772) <= 11589095;
srom_1(54773) <= 12112269;
srom_1(54774) <= 12617982;
srom_1(54775) <= 13103861;
srom_1(54776) <= 13567629;
srom_1(54777) <= 14007110;
srom_1(54778) <= 14420245;
srom_1(54779) <= 14805095;
srom_1(54780) <= 15159856;
srom_1(54781) <= 15482864;
srom_1(54782) <= 15772605;
srom_1(54783) <= 16027720;
srom_1(54784) <= 16247012;
srom_1(54785) <= 16429454;
srom_1(54786) <= 16574189;
srom_1(54787) <= 16680539;
srom_1(54788) <= 16748006;
srom_1(54789) <= 16776272;
srom_1(54790) <= 16765206;
srom_1(54791) <= 16714859;
srom_1(54792) <= 16625467;
srom_1(54793) <= 16497450;
srom_1(54794) <= 16331408;
srom_1(54795) <= 16128119;
srom_1(54796) <= 15888537;
srom_1(54797) <= 15613786;
srom_1(54798) <= 15305153;
srom_1(54799) <= 14964085;
srom_1(54800) <= 14592184;
srom_1(54801) <= 14191191;
srom_1(54802) <= 13762988;
srom_1(54803) <= 13309583;
srom_1(54804) <= 12833102;
srom_1(54805) <= 12335779;
srom_1(54806) <= 11819946;
srom_1(54807) <= 11288022;
srom_1(54808) <= 10742503;
srom_1(54809) <= 10185944;
srom_1(54810) <= 9620958;
srom_1(54811) <= 9050193;
srom_1(54812) <= 8476325;
srom_1(54813) <= 7902046;
srom_1(54814) <= 7330049;
srom_1(54815) <= 6763015;
srom_1(54816) <= 6203605;
srom_1(54817) <= 5654440;
srom_1(54818) <= 5118098;
srom_1(54819) <= 4597091;
srom_1(54820) <= 4093865;
srom_1(54821) <= 3610778;
srom_1(54822) <= 3150095;
srom_1(54823) <= 2713978;
srom_1(54824) <= 2304472;
srom_1(54825) <= 1923496;
srom_1(54826) <= 1572837;
srom_1(54827) <= 1254139;
srom_1(54828) <= 968898;
srom_1(54829) <= 718450;
srom_1(54830) <= 503970;
srom_1(54831) <= 326463;
srom_1(54832) <= 186763;
srom_1(54833) <= 85525;
srom_1(54834) <= 23222;
srom_1(54835) <= 147;
srom_1(54836) <= 16409;
srom_1(54837) <= 71931;
srom_1(54838) <= 166452;
srom_1(54839) <= 299531;
srom_1(54840) <= 470541;
srom_1(54841) <= 678682;
srom_1(54842) <= 922978;
srom_1(54843) <= 1202282;
srom_1(54844) <= 1515286;
srom_1(54845) <= 1860521;
srom_1(54846) <= 2236368;
srom_1(54847) <= 2641066;
srom_1(54848) <= 3072715;
srom_1(54849) <= 3529293;
srom_1(54850) <= 4008658;
srom_1(54851) <= 4508561;
srom_1(54852) <= 5026660;
srom_1(54853) <= 5560524;
srom_1(54854) <= 6107649;
srom_1(54855) <= 6665471;
srom_1(54856) <= 7231374;
srom_1(54857) <= 7802703;
srom_1(54858) <= 8376779;
srom_1(54859) <= 8950911;
srom_1(54860) <= 9522406;
srom_1(54861) <= 10088584;
srom_1(54862) <= 10646791;
srom_1(54863) <= 11194408;
srom_1(54864) <= 11728868;
srom_1(54865) <= 12247664;
srom_1(54866) <= 12748364;
srom_1(54867) <= 13228619;
srom_1(54868) <= 13686178;
srom_1(54869) <= 14118894;
srom_1(54870) <= 14524740;
srom_1(54871) <= 14901811;
srom_1(54872) <= 15248339;
srom_1(54873) <= 15562700;
srom_1(54874) <= 15843419;
srom_1(54875) <= 16089179;
srom_1(54876) <= 16298829;
srom_1(54877) <= 16471386;
srom_1(54878) <= 16606039;
srom_1(54879) <= 16702158;
srom_1(54880) <= 16759292;
srom_1(54881) <= 16777173;
srom_1(54882) <= 16755717;
srom_1(54883) <= 16695025;
srom_1(54884) <= 16595381;
srom_1(54885) <= 16457252;
srom_1(54886) <= 16281288;
srom_1(54887) <= 16068311;
srom_1(54888) <= 15819322;
srom_1(54889) <= 15535488;
srom_1(54890) <= 15218139;
srom_1(54891) <= 14868765;
srom_1(54892) <= 14489002;
srom_1(54893) <= 14080633;
srom_1(54894) <= 13645572;
srom_1(54895) <= 13185860;
srom_1(54896) <= 12703651;
srom_1(54897) <= 12201207;
srom_1(54898) <= 11680885;
srom_1(54899) <= 11145125;
srom_1(54900) <= 10596438;
srom_1(54901) <= 10037398;
srom_1(54902) <= 9470626;
srom_1(54903) <= 8898780;
srom_1(54904) <= 8324542;
srom_1(54905) <= 7750604;
srom_1(54906) <= 7179658;
srom_1(54907) <= 6614381;
srom_1(54908) <= 6057424;
srom_1(54909) <= 5511399;
srom_1(54910) <= 4978866;
srom_1(54911) <= 4462323;
srom_1(54912) <= 3964191;
srom_1(54913) <= 3486807;
srom_1(54914) <= 3032409;
srom_1(54915) <= 2603128;
srom_1(54916) <= 2200977;
srom_1(54917) <= 1827842;
srom_1(54918) <= 1485473;
srom_1(54919) <= 1175475;
srom_1(54920) <= 899301;
srom_1(54921) <= 658248;
srom_1(54922) <= 453445;
srom_1(54923) <= 285853;
srom_1(54924) <= 156257;
srom_1(54925) <= 65266;
srom_1(54926) <= 13305;
srom_1(54927) <= 620;
srom_1(54928) <= 27268;
srom_1(54929) <= 93126;
srom_1(54930) <= 197884;
srom_1(54931) <= 341051;
srom_1(54932) <= 521956;
srom_1(54933) <= 739750;
srom_1(54934) <= 993412;
srom_1(54935) <= 1281753;
srom_1(54936) <= 1603421;
srom_1(54937) <= 1956906;
srom_1(54938) <= 2340552;
srom_1(54939) <= 2752560;
srom_1(54940) <= 3190997;
srom_1(54941) <= 3653807;
srom_1(54942) <= 4138820;
srom_1(54943) <= 4643762;
srom_1(54944) <= 5166265;
srom_1(54945) <= 5703878;
srom_1(54946) <= 6254081;
srom_1(54947) <= 6814294;
srom_1(54948) <= 7381889;
srom_1(54949) <= 7954205;
srom_1(54950) <= 8528558;
srom_1(54951) <= 9102255;
srom_1(54952) <= 9672605;
srom_1(54953) <= 10236934;
srom_1(54954) <= 10792596;
srom_1(54955) <= 11336984;
srom_1(54956) <= 11867547;
srom_1(54957) <= 12381795;
srom_1(54958) <= 12877318;
srom_1(54959) <= 13351792;
srom_1(54960) <= 13802992;
srom_1(54961) <= 14228802;
srom_1(54962) <= 14627226;
srom_1(54963) <= 14996394;
srom_1(54964) <= 15334576;
srom_1(54965) <= 15640186;
srom_1(54966) <= 15911791;
srom_1(54967) <= 16148118;
srom_1(54968) <= 16348057;
srom_1(54969) <= 16510671;
srom_1(54970) <= 16635199;
srom_1(54971) <= 16721055;
srom_1(54972) <= 16767838;
srom_1(54973) <= 16775327;
srom_1(54974) <= 16743488;
srom_1(54975) <= 16672471;
srom_1(54976) <= 16562607;
srom_1(54977) <= 16414413;
srom_1(54978) <= 16228583;
srom_1(54979) <= 16005989;
srom_1(54980) <= 15747674;
srom_1(54981) <= 15454850;
srom_1(54982) <= 15128890;
srom_1(54983) <= 14771322;
srom_1(54984) <= 14383824;
srom_1(54985) <= 13968212;
srom_1(54986) <= 13526435;
srom_1(54987) <= 13060565;
srom_1(54988) <= 12572787;
srom_1(54989) <= 12065388;
srom_1(54990) <= 11540747;
srom_1(54991) <= 11001325;
srom_1(54992) <= 10449651;
srom_1(54993) <= 9888311;
srom_1(54994) <= 9319940;
srom_1(54995) <= 8747200;
srom_1(54996) <= 8172780;
srom_1(54997) <= 7599371;
srom_1(54998) <= 7029663;
srom_1(54999) <= 6466328;
srom_1(55000) <= 5912007;
srom_1(55001) <= 5369300;
srom_1(55002) <= 4840751;
srom_1(55003) <= 4328840;
srom_1(55004) <= 3835966;
srom_1(55005) <= 3364441;
srom_1(55006) <= 2916476;
srom_1(55007) <= 2494171;
srom_1(55008) <= 2099508;
srom_1(55009) <= 1734336;
srom_1(55010) <= 1400369;
srom_1(55011) <= 1099172;
srom_1(55012) <= 832157;
srom_1(55013) <= 600578;
srom_1(55014) <= 405519;
srom_1(55015) <= 247895;
srom_1(55016) <= 128446;
srom_1(55017) <= 47732;
srom_1(55018) <= 6131;
srom_1(55019) <= 3839;
srom_1(55020) <= 40865;
srom_1(55021) <= 117037;
srom_1(55022) <= 231997;
srom_1(55023) <= 385206;
srom_1(55024) <= 575946;
srom_1(55025) <= 803322;
srom_1(55026) <= 1066268;
srom_1(55027) <= 1363551;
srom_1(55028) <= 1693777;
srom_1(55029) <= 2055398;
srom_1(55030) <= 2446717;
srom_1(55031) <= 2865899;
srom_1(55032) <= 3310980;
srom_1(55033) <= 3779871;
srom_1(55034) <= 4270374;
srom_1(55035) <= 4780189;
srom_1(55036) <= 5306925;
srom_1(55037) <= 5848112;
srom_1(55038) <= 6401212;
srom_1(55039) <= 6963632;
srom_1(55040) <= 7532734;
srom_1(55041) <= 8105850;
srom_1(55042) <= 8680291;
srom_1(55043) <= 9253365;
srom_1(55044) <= 9822383;
srom_1(55045) <= 10384678;
srom_1(55046) <= 10937613;
srom_1(55047) <= 11478595;
srom_1(55048) <= 12005086;
srom_1(55049) <= 12514619;
srom_1(55050) <= 13004804;
srom_1(55051) <= 13473341;
srom_1(55052) <= 13918035;
srom_1(55053) <= 14336799;
srom_1(55054) <= 14727669;
srom_1(55055) <= 15088814;
srom_1(55056) <= 15418540;
srom_1(55057) <= 15715299;
srom_1(55058) <= 15977701;
srom_1(55059) <= 16204516;
srom_1(55060) <= 16394678;
srom_1(55061) <= 16547298;
srom_1(55062) <= 16661659;
srom_1(55063) <= 16737224;
srom_1(55064) <= 16773640;
srom_1(55065) <= 16770736;
srom_1(55066) <= 16728525;
srom_1(55067) <= 16647205;
srom_1(55068) <= 16527158;
srom_1(55069) <= 16368946;
srom_1(55070) <= 16173312;
srom_1(55071) <= 15941172;
srom_1(55072) <= 15673616;
srom_1(55073) <= 15371899;
srom_1(55074) <= 15037434;
srom_1(55075) <= 14671790;
srom_1(55076) <= 14276683;
srom_1(55077) <= 13853964;
srom_1(55078) <= 13405616;
srom_1(55079) <= 12933742;
srom_1(55080) <= 12440554;
srom_1(55081) <= 11928365;
srom_1(55082) <= 11399577;
srom_1(55083) <= 10856670;
srom_1(55084) <= 10302189;
srom_1(55085) <= 9738734;
srom_1(55086) <= 9168948;
srom_1(55087) <= 8595503;
srom_1(55088) <= 8021088;
srom_1(55089) <= 7448396;
srom_1(55090) <= 6880113;
srom_1(55091) <= 6318904;
srom_1(55092) <= 5767401;
srom_1(55093) <= 5228189;
srom_1(55094) <= 4703798;
srom_1(55095) <= 4196686;
srom_1(55096) <= 3709231;
srom_1(55097) <= 3243719;
srom_1(55098) <= 2802334;
srom_1(55099) <= 2387145;
srom_1(55100) <= 2000098;
srom_1(55101) <= 1643009;
srom_1(55102) <= 1317553;
srom_1(55103) <= 1025256;
srom_1(55104) <= 767487;
srom_1(55105) <= 545457;
srom_1(55106) <= 360206;
srom_1(55107) <= 212603;
srom_1(55108) <= 103340;
srom_1(55109) <= 32929;
srom_1(55110) <= 1701;
srom_1(55111) <= 9802;
srom_1(55112) <= 57195;
srom_1(55113) <= 143656;
srom_1(55114) <= 268780;
srom_1(55115) <= 431981;
srom_1(55116) <= 632494;
srom_1(55117) <= 869377;
srom_1(55118) <= 1141521;
srom_1(55119) <= 1447649;
srom_1(55120) <= 1786326;
srom_1(55121) <= 2155962;
srom_1(55122) <= 2554826;
srom_1(55123) <= 2981047;
srom_1(55124) <= 3432625;
srom_1(55125) <= 3907444;
srom_1(55126) <= 4403276;
srom_1(55127) <= 4917797;
srom_1(55128) <= 5448594;
srom_1(55129) <= 5993177;
srom_1(55130) <= 6548993;
srom_1(55131) <= 7113436;
srom_1(55132) <= 7683859;
srom_1(55133) <= 8257587;
srom_1(55134) <= 8831929;
srom_1(55135) <= 9404192;
srom_1(55136) <= 9971692;
srom_1(55137) <= 10531769;
srom_1(55138) <= 11081796;
srom_1(55139) <= 11619194;
srom_1(55140) <= 12141442;
srom_1(55141) <= 12646092;
srom_1(55142) <= 13130778;
srom_1(55143) <= 13593225;
srom_1(55144) <= 14031266;
srom_1(55145) <= 14442847;
srom_1(55146) <= 14826038;
srom_1(55147) <= 15179041;
srom_1(55148) <= 15500201;
srom_1(55149) <= 15788013;
srom_1(55150) <= 16041126;
srom_1(55151) <= 16258355;
srom_1(55152) <= 16438679;
srom_1(55153) <= 16581253;
srom_1(55154) <= 16685410;
srom_1(55155) <= 16750660;
srom_1(55156) <= 16776697;
srom_1(55157) <= 16763400;
srom_1(55158) <= 16710830;
srom_1(55159) <= 16619235;
srom_1(55160) <= 16489043;
srom_1(55161) <= 16320866;
srom_1(55162) <= 16115492;
srom_1(55163) <= 15873883;
srom_1(55164) <= 15597174;
srom_1(55165) <= 15286661;
srom_1(55166) <= 14943801;
srom_1(55167) <= 14570201;
srom_1(55168) <= 14167614;
srom_1(55169) <= 13737926;
srom_1(55170) <= 13283154;
srom_1(55171) <= 12805430;
srom_1(55172) <= 12306994;
srom_1(55173) <= 11790183;
srom_1(55174) <= 11257421;
srom_1(55175) <= 10711206;
srom_1(55176) <= 10154100;
srom_1(55177) <= 9588715;
srom_1(55178) <= 9017702;
srom_1(55179) <= 8443738;
srom_1(55180) <= 7869517;
srom_1(55181) <= 7297729;
srom_1(55182) <= 6731057;
srom_1(55183) <= 6172158;
srom_1(55184) <= 5623653;
srom_1(55185) <= 5088113;
srom_1(55186) <= 4568051;
srom_1(55187) <= 4065904;
srom_1(55188) <= 3584028;
srom_1(55189) <= 3124683;
srom_1(55190) <= 2690021;
srom_1(55191) <= 2282083;
srom_1(55192) <= 1902780;
srom_1(55193) <= 1553891;
srom_1(55194) <= 1237052;
srom_1(55195) <= 953750;
srom_1(55196) <= 705312;
srom_1(55197) <= 492904;
srom_1(55198) <= 317521;
srom_1(55199) <= 179987;
srom_1(55200) <= 80946;
srom_1(55201) <= 20862;
srom_1(55202) <= 17;
srom_1(55203) <= 18509;
srom_1(55204) <= 76252;
srom_1(55205) <= 172974;
srom_1(55206) <= 308222;
srom_1(55207) <= 481362;
srom_1(55208) <= 691581;
srom_1(55209) <= 937895;
srom_1(55210) <= 1219147;
srom_1(55211) <= 1534019;
srom_1(55212) <= 1881035;
srom_1(55213) <= 2258568;
srom_1(55214) <= 2664846;
srom_1(55215) <= 3097964;
srom_1(55216) <= 3555893;
srom_1(55217) <= 4036484;
srom_1(55218) <= 4537483;
srom_1(55219) <= 5056541;
srom_1(55220) <= 5591225;
srom_1(55221) <= 6139027;
srom_1(55222) <= 6697377;
srom_1(55223) <= 7263659;
srom_1(55224) <= 7835215;
srom_1(55225) <= 8409367;
srom_1(55226) <= 8983421;
srom_1(55227) <= 9554686;
srom_1(55228) <= 10120483;
srom_1(55229) <= 10678159;
srom_1(55230) <= 11225098;
srom_1(55231) <= 11758735;
srom_1(55232) <= 12276570;
srom_1(55233) <= 12776172;
srom_1(55234) <= 13255199;
srom_1(55235) <= 13711405;
srom_1(55236) <= 14142651;
srom_1(55237) <= 14546914;
srom_1(55238) <= 14922298;
srom_1(55239) <= 15267044;
srom_1(55240) <= 15579535;
srom_1(55241) <= 15858305;
srom_1(55242) <= 16102046;
srom_1(55243) <= 16309617;
srom_1(55244) <= 16480044;
srom_1(55245) <= 16612527;
srom_1(55246) <= 16706445;
srom_1(55247) <= 16761358;
srom_1(55248) <= 16777008;
srom_1(55249) <= 16753322;
srom_1(55250) <= 16690411;
srom_1(55251) <= 16588571;
srom_1(55252) <= 16448277;
srom_1(55253) <= 16270189;
srom_1(55254) <= 16055142;
srom_1(55255) <= 15804144;
srom_1(55256) <= 15518371;
srom_1(55257) <= 15199165;
srom_1(55258) <= 14848022;
srom_1(55259) <= 14466588;
srom_1(55260) <= 14056653;
srom_1(55261) <= 13620138;
srom_1(55262) <= 13159090;
srom_1(55263) <= 12675673;
srom_1(55264) <= 12172151;
srom_1(55265) <= 11650888;
srom_1(55266) <= 11114326;
srom_1(55267) <= 10564983;
srom_1(55268) <= 10005433;
srom_1(55269) <= 9438302;
srom_1(55270) <= 8866249;
srom_1(55271) <= 8291956;
srom_1(55272) <= 7718116;
srom_1(55273) <= 7147420;
srom_1(55274) <= 6582544;
srom_1(55275) <= 6026138;
srom_1(55276) <= 5480810;
srom_1(55277) <= 4949118;
srom_1(55278) <= 4433554;
srom_1(55279) <= 3936538;
srom_1(55280) <= 3460398;
srom_1(55281) <= 3007369;
srom_1(55282) <= 2579574;
srom_1(55283) <= 2179020;
srom_1(55284) <= 1807585;
srom_1(55285) <= 1467010;
srom_1(55286) <= 1158893;
srom_1(55287) <= 884678;
srom_1(55288) <= 645653;
srom_1(55289) <= 442936;
srom_1(55290) <= 277479;
srom_1(55291) <= 150059;
srom_1(55292) <= 61271;
srom_1(55293) <= 11534;
srom_1(55294) <= 1079;
srom_1(55295) <= 29957;
srom_1(55296) <= 98031;
srom_1(55297) <= 204982;
srom_1(55298) <= 350309;
srom_1(55299) <= 533331;
srom_1(55300) <= 753188;
srom_1(55301) <= 1008851;
srom_1(55302) <= 1299120;
srom_1(55303) <= 1622634;
srom_1(55304) <= 1977876;
srom_1(55305) <= 2363180;
srom_1(55306) <= 2776739;
srom_1(55307) <= 3216614;
srom_1(55308) <= 3680743;
srom_1(55309) <= 4166948;
srom_1(55310) <= 4672950;
srom_1(55311) <= 5196377;
srom_1(55312) <= 5734772;
srom_1(55313) <= 6285613;
srom_1(55314) <= 6846315;
srom_1(55315) <= 7414249;
srom_1(55316) <= 7986752;
srom_1(55317) <= 8561140;
srom_1(55318) <= 9134719;
srom_1(55319) <= 9704799;
srom_1(55320) <= 10268707;
srom_1(55321) <= 10823798;
srom_1(55322) <= 11367470;
srom_1(55323) <= 11897174;
srom_1(55324) <= 12410424;
srom_1(55325) <= 12904814;
srom_1(55326) <= 13378027;
srom_1(55327) <= 13827842;
srom_1(55328) <= 14252151;
srom_1(55329) <= 14648964;
srom_1(55330) <= 15016420;
srom_1(55331) <= 15352796;
srom_1(55332) <= 15656514;
srom_1(55333) <= 15926150;
srom_1(55334) <= 16160441;
srom_1(55335) <= 16358286;
srom_1(55336) <= 16518760;
srom_1(55337) <= 16641107;
srom_1(55338) <= 16724757;
srom_1(55339) <= 16769315;
srom_1(55340) <= 16774573;
srom_1(55341) <= 16740506;
srom_1(55342) <= 16667275;
srom_1(55343) <= 16555222;
srom_1(55344) <= 16404872;
srom_1(55345) <= 16216932;
srom_1(55346) <= 15992282;
srom_1(55347) <= 15731976;
srom_1(55348) <= 15437235;
srom_1(55349) <= 15109439;
srom_1(55350) <= 14750128;
srom_1(55351) <= 14360985;
srom_1(55352) <= 13943836;
srom_1(55353) <= 13500636;
srom_1(55354) <= 13033464;
srom_1(55355) <= 12544511;
srom_1(55356) <= 12036070;
srom_1(55357) <= 11510524;
srom_1(55358) <= 10970338;
srom_1(55359) <= 10418046;
srom_1(55360) <= 9856237;
srom_1(55361) <= 9287546;
srom_1(55362) <= 8714640;
srom_1(55363) <= 8140204;
srom_1(55364) <= 7566934;
srom_1(55365) <= 6997516;
srom_1(55366) <= 6434622;
srom_1(55367) <= 5880891;
srom_1(55368) <= 5338919;
srom_1(55369) <= 4811248;
srom_1(55370) <= 4300353;
srom_1(55371) <= 3808629;
srom_1(55372) <= 3338382;
srom_1(55373) <= 2891817;
srom_1(55374) <= 2471029;
srom_1(55375) <= 2077990;
srom_1(55376) <= 1714544;
srom_1(55377) <= 1382395;
srom_1(55378) <= 1083100;
srom_1(55379) <= 818064;
srom_1(55380) <= 588528;
srom_1(55381) <= 395569;
srom_1(55382) <= 240093;
srom_1(55383) <= 122828;
srom_1(55384) <= 44324;
srom_1(55385) <= 4949;
srom_1(55386) <= 4888;
srom_1(55387) <= 44141;
srom_1(55388) <= 122524;
srom_1(55389) <= 239669;
srom_1(55390) <= 395028;
srom_1(55391) <= 587872;
srom_1(55392) <= 817295;
srom_1(55393) <= 1082224;
srom_1(55394) <= 1381414;
srom_1(55395) <= 1713463;
srom_1(55396) <= 2076815;
srom_1(55397) <= 2469765;
srom_1(55398) <= 2890470;
srom_1(55399) <= 3336958;
srom_1(55400) <= 3807134;
srom_1(55401) <= 4298795;
srom_1(55402) <= 4809635;
srom_1(55403) <= 5337257;
srom_1(55404) <= 5879188;
srom_1(55405) <= 6432887;
srom_1(55406) <= 6995757;
srom_1(55407) <= 7565158;
srom_1(55408) <= 8138421;
srom_1(55409) <= 8712857;
srom_1(55410) <= 9285772;
srom_1(55411) <= 9854481;
srom_1(55412) <= 10416315;
srom_1(55413) <= 10968641;
srom_1(55414) <= 11508868;
srom_1(55415) <= 12034463;
srom_1(55416) <= 12542961;
srom_1(55417) <= 13031979;
srom_1(55418) <= 13499221;
srom_1(55419) <= 13942499;
srom_1(55420) <= 14359732;
srom_1(55421) <= 14748965;
srom_1(55422) <= 15108372;
srom_1(55423) <= 15436267;
srom_1(55424) <= 15731114;
srom_1(55425) <= 15991529;
srom_1(55426) <= 16216291;
srom_1(55427) <= 16404347;
srom_1(55428) <= 16554814;
srom_1(55429) <= 16666986;
srom_1(55430) <= 16740339;
srom_1(55431) <= 16774528;
srom_1(55432) <= 16769392;
srom_1(55433) <= 16724956;
srom_1(55434) <= 16641427;
srom_1(55435) <= 16519199;
srom_1(55436) <= 16358843;
srom_1(55437) <= 16161112;
srom_1(55438) <= 15926933;
srom_1(55439) <= 15657405;
srom_1(55440) <= 15353790;
srom_1(55441) <= 15017513;
srom_1(55442) <= 14650152;
srom_1(55443) <= 14253427;
srom_1(55444) <= 13829200;
srom_1(55445) <= 13379461;
srom_1(55446) <= 12906318;
srom_1(55447) <= 12411989;
srom_1(55448) <= 11898794;
srom_1(55449) <= 11369138;
srom_1(55450) <= 10825506;
srom_1(55451) <= 10270446;
srom_1(55452) <= 9706561;
srom_1(55453) <= 9136496;
srom_1(55454) <= 8562924;
srom_1(55455) <= 7988534;
srom_1(55456) <= 7416021;
srom_1(55457) <= 6848068;
srom_1(55458) <= 6287340;
srom_1(55459) <= 5736465;
srom_1(55460) <= 5198027;
srom_1(55461) <= 4674550;
srom_1(55462) <= 4168490;
srom_1(55463) <= 3682220;
srom_1(55464) <= 3218019;
srom_1(55465) <= 2778065;
srom_1(55466) <= 2364421;
srom_1(55467) <= 1979027;
srom_1(55468) <= 1623689;
srom_1(55469) <= 1300074;
srom_1(55470) <= 1009699;
srom_1(55471) <= 753927;
srom_1(55472) <= 533957;
srom_1(55473) <= 350820;
srom_1(55474) <= 205374;
srom_1(55475) <= 98303;
srom_1(55476) <= 30108;
srom_1(55477) <= 1108;
srom_1(55478) <= 11441;
srom_1(55479) <= 61056;
srom_1(55480) <= 149723;
srom_1(55481) <= 277025;
srom_1(55482) <= 442364;
srom_1(55483) <= 644966;
srom_1(55484) <= 883881;
srom_1(55485) <= 1157988;
srom_1(55486) <= 1466002;
srom_1(55487) <= 1806478;
srom_1(55488) <= 2177821;
srom_1(55489) <= 2578287;
srom_1(55490) <= 3006001;
srom_1(55491) <= 3458955;
srom_1(55492) <= 3935026;
srom_1(55493) <= 4431981;
srom_1(55494) <= 4947491;
srom_1(55495) <= 5479136;
srom_1(55496) <= 6024426;
srom_1(55497) <= 6580802;
srom_1(55498) <= 7145655;
srom_1(55499) <= 7716337;
srom_1(55500) <= 8290172;
srom_1(55501) <= 8864468;
srom_1(55502) <= 9436532;
srom_1(55503) <= 10003683;
srom_1(55504) <= 10563259;
srom_1(55505) <= 11112639;
srom_1(55506) <= 11649244;
srom_1(55507) <= 12170559;
srom_1(55508) <= 12674139;
srom_1(55509) <= 13157623;
srom_1(55510) <= 13618743;
srom_1(55511) <= 14055337;
srom_1(55512) <= 14465358;
srom_1(55513) <= 14846883;
srom_1(55514) <= 15198123;
srom_1(55515) <= 15517431;
srom_1(55516) <= 15803309;
srom_1(55517) <= 16054418;
srom_1(55518) <= 16269578;
srom_1(55519) <= 16447782;
srom_1(55520) <= 16588194;
srom_1(55521) <= 16690155;
srom_1(55522) <= 16753188;
srom_1(55523) <= 16776995;
srom_1(55524) <= 16761467;
srom_1(55525) <= 16706676;
srom_1(55526) <= 16612878;
srom_1(55527) <= 16480514;
srom_1(55528) <= 16310204;
srom_1(55529) <= 16102747;
srom_1(55530) <= 15859116;
srom_1(55531) <= 15580453;
srom_1(55532) <= 15268065;
srom_1(55533) <= 14923417;
srom_1(55534) <= 14548125;
srom_1(55535) <= 14143949;
srom_1(55536) <= 13712784;
srom_1(55537) <= 13256652;
srom_1(55538) <= 12777692;
srom_1(55539) <= 12278150;
srom_1(55540) <= 11760369;
srom_1(55541) <= 11226777;
srom_1(55542) <= 10679875;
srom_1(55543) <= 10122229;
srom_1(55544) <= 9556453;
srom_1(55545) <= 8985201;
srom_1(55546) <= 8411151;
srom_1(55547) <= 7836995;
srom_1(55548) <= 7265427;
srom_1(55549) <= 6699125;
srom_1(55550) <= 6140745;
srom_1(55551) <= 5592907;
srom_1(55552) <= 5058179;
srom_1(55553) <= 4539068;
srom_1(55554) <= 4038009;
srom_1(55555) <= 3557351;
srom_1(55556) <= 3099349;
srom_1(55557) <= 2666150;
srom_1(55558) <= 2259786;
srom_1(55559) <= 1882161;
srom_1(55560) <= 1535048;
srom_1(55561) <= 1220073;
srom_1(55562) <= 938715;
srom_1(55563) <= 692291;
srom_1(55564) <= 481958;
srom_1(55565) <= 308701;
srom_1(55566) <= 173335;
srom_1(55567) <= 76492;
srom_1(55568) <= 18628;
srom_1(55569) <= 14;
srom_1(55570) <= 20736;
srom_1(55571) <= 80699;
srom_1(55572) <= 179620;
srom_1(55573) <= 317035;
srom_1(55574) <= 492302;
srom_1(55575) <= 704596;
srom_1(55576) <= 952924;
srom_1(55577) <= 1236120;
srom_1(55578) <= 1552856;
srom_1(55579) <= 1901648;
srom_1(55580) <= 2280860;
srom_1(55581) <= 2688712;
srom_1(55582) <= 3123294;
srom_1(55583) <= 3582566;
srom_1(55584) <= 4064375;
srom_1(55585) <= 4566462;
srom_1(55586) <= 5086473;
srom_1(55587) <= 5621968;
srom_1(55588) <= 6170438;
srom_1(55589) <= 6729308;
srom_1(55590) <= 7295960;
srom_1(55591) <= 7867736;
srom_1(55592) <= 8441954;
srom_1(55593) <= 9015922;
srom_1(55594) <= 9586949;
srom_1(55595) <= 10152356;
srom_1(55596) <= 10709492;
srom_1(55597) <= 11255745;
srom_1(55598) <= 11788552;
srom_1(55599) <= 12305416;
srom_1(55600) <= 12803913;
srom_1(55601) <= 13281705;
srom_1(55602) <= 13736552;
srom_1(55603) <= 14166320;
srom_1(55604) <= 14568995;
srom_1(55605) <= 14942687;
srom_1(55606) <= 15285646;
srom_1(55607) <= 15596261;
srom_1(55608) <= 15873078;
srom_1(55609) <= 16114797;
srom_1(55610) <= 16320285;
srom_1(55611) <= 16488580;
srom_1(55612) <= 16618890;
srom_1(55613) <= 16710606;
srom_1(55614) <= 16763297;
srom_1(55615) <= 16776717;
srom_1(55616) <= 16750801;
srom_1(55617) <= 16685673;
srom_1(55618) <= 16581637;
srom_1(55619) <= 16439180;
srom_1(55620) <= 16258972;
srom_1(55621) <= 16041857;
srom_1(55622) <= 15788853;
srom_1(55623) <= 15501147;
srom_1(55624) <= 15180088;
srom_1(55625) <= 14827181;
srom_1(55626) <= 14444082;
srom_1(55627) <= 14032586;
srom_1(55628) <= 13594624;
srom_1(55629) <= 13132249;
srom_1(55630) <= 12647630;
srom_1(55631) <= 12143038;
srom_1(55632) <= 11620840;
srom_1(55633) <= 11083486;
srom_1(55634) <= 10533494;
srom_1(55635) <= 9973444;
srom_1(55636) <= 9405963;
srom_1(55637) <= 8833710;
srom_1(55638) <= 8259371;
srom_1(55639) <= 7685637;
srom_1(55640) <= 7115200;
srom_1(55641) <= 6550734;
srom_1(55642) <= 5994887;
srom_1(55643) <= 5450265;
srom_1(55644) <= 4919421;
srom_1(55645) <= 4404846;
srom_1(55646) <= 3908952;
srom_1(55647) <= 3434065;
srom_1(55648) <= 2982411;
srom_1(55649) <= 2556108;
srom_1(55650) <= 2157157;
srom_1(55651) <= 1787426;
srom_1(55652) <= 1448651;
srom_1(55653) <= 1142420;
srom_1(55654) <= 870169;
srom_1(55655) <= 633174;
srom_1(55656) <= 432547;
srom_1(55657) <= 269228;
srom_1(55658) <= 143985;
srom_1(55659) <= 57403;
srom_1(55660) <= 9889;
srom_1(55661) <= 1665;
srom_1(55662) <= 32771;
srom_1(55663) <= 103061;
srom_1(55664) <= 212204;
srom_1(55665) <= 359689;
srom_1(55666) <= 544824;
srom_1(55667) <= 766742;
srom_1(55668) <= 1024401;
srom_1(55669) <= 1316593;
srom_1(55670) <= 1641949;
srom_1(55671) <= 1998942;
srom_1(55672) <= 2385898;
srom_1(55673) <= 2801003;
srom_1(55674) <= 3242310;
srom_1(55675) <= 3707750;
srom_1(55676) <= 4195140;
srom_1(55677) <= 4702195;
srom_1(55678) <= 5226537;
srom_1(55679) <= 5765706;
srom_1(55680) <= 6317175;
srom_1(55681) <= 6878358;
srom_1(55682) <= 7446623;
srom_1(55683) <= 8019306;
srom_1(55684) <= 8593720;
srom_1(55685) <= 9167172;
srom_1(55686) <= 9736973;
srom_1(55687) <= 10300451;
srom_1(55688) <= 10854964;
srom_1(55689) <= 11397912;
srom_1(55690) <= 11926748;
srom_1(55691) <= 12438992;
srom_1(55692) <= 12932242;
srom_1(55693) <= 13404186;
srom_1(55694) <= 13852610;
srom_1(55695) <= 14275412;
srom_1(55696) <= 14670608;
srom_1(55697) <= 15036346;
srom_1(55698) <= 15370910;
srom_1(55699) <= 15672732;
srom_1(55700) <= 15940396;
srom_1(55701) <= 16172647;
srom_1(55702) <= 16368396;
srom_1(55703) <= 16526725;
srom_1(55704) <= 16646892;
srom_1(55705) <= 16728332;
srom_1(55706) <= 16770665;
srom_1(55707) <= 16773692;
srom_1(55708) <= 16737398;
srom_1(55709) <= 16661953;
srom_1(55710) <= 16547713;
srom_1(55711) <= 16395211;
srom_1(55712) <= 16205163;
srom_1(55713) <= 15978461;
srom_1(55714) <= 15716168;
srom_1(55715) <= 15419513;
srom_1(55716) <= 15089888;
srom_1(55717) <= 14728838;
srom_1(55718) <= 14338056;
srom_1(55719) <= 13919376;
srom_1(55720) <= 13474760;
srom_1(55721) <= 13006293;
srom_1(55722) <= 12516173;
srom_1(55723) <= 12006696;
srom_1(55724) <= 11480253;
srom_1(55725) <= 10939313;
srom_1(55726) <= 10386411;
srom_1(55727) <= 9824141;
srom_1(55728) <= 9255139;
srom_1(55729) <= 8682074;
srom_1(55730) <= 8107633;
srom_1(55731) <= 7534509;
srom_1(55732) <= 6965390;
srom_1(55733) <= 6402945;
srom_1(55734) <= 5849812;
srom_1(55735) <= 5308584;
srom_1(55736) <= 4781799;
srom_1(55737) <= 4271928;
srom_1(55738) <= 3781362;
srom_1(55739) <= 3312400;
srom_1(55740) <= 2867242;
srom_1(55741) <= 2447976;
srom_1(55742) <= 2056568;
srom_1(55743) <= 1694853;
srom_1(55744) <= 1364527;
srom_1(55745) <= 1067139;
srom_1(55746) <= 804084;
srom_1(55747) <= 576596;
srom_1(55748) <= 385741;
srom_1(55749) <= 232414;
srom_1(55750) <= 117334;
srom_1(55751) <= 41041;
srom_1(55752) <= 3893;
srom_1(55753) <= 6063;
srom_1(55754) <= 47542;
srom_1(55755) <= 128135;
srom_1(55756) <= 247465;
srom_1(55757) <= 404971;
srom_1(55758) <= 599915;
srom_1(55759) <= 831383;
srom_1(55760) <= 1098289;
srom_1(55761) <= 1399382;
srom_1(55762) <= 1733250;
srom_1(55763) <= 2098327;
srom_1(55764) <= 2492902;
srom_1(55765) <= 2915123;
srom_1(55766) <= 3363012;
srom_1(55767) <= 3834467;
srom_1(55768) <= 4327278;
srom_1(55769) <= 4839135;
srom_1(55770) <= 5367635;
srom_1(55771) <= 5910303;
srom_1(55772) <= 6464592;
srom_1(55773) <= 7027903;
srom_1(55774) <= 7597595;
srom_1(55775) <= 8170996;
srom_1(55776) <= 8745418;
srom_1(55777) <= 9318166;
srom_1(55778) <= 9886556;
srom_1(55779) <= 10447921;
srom_1(55780) <= 10999629;
srom_1(55781) <= 11539094;
srom_1(55782) <= 12063784;
srom_1(55783) <= 12571241;
srom_1(55784) <= 13059084;
srom_1(55785) <= 13525025;
srom_1(55786) <= 13966879;
srom_1(55787) <= 14382576;
srom_1(55788) <= 14770164;
srom_1(55789) <= 15127827;
srom_1(55790) <= 15453888;
srom_1(55791) <= 15746817;
srom_1(55792) <= 16005241;
srom_1(55793) <= 16227948;
srom_1(55794) <= 16413894;
srom_1(55795) <= 16562206;
srom_1(55796) <= 16672189;
srom_1(55797) <= 16743328;
srom_1(55798) <= 16775289;
srom_1(55799) <= 16767922;
srom_1(55800) <= 16721261;
srom_1(55801) <= 16635525;
srom_1(55802) <= 16511117;
srom_1(55803) <= 16348620;
srom_1(55804) <= 16148795;
srom_1(55805) <= 15912581;
srom_1(55806) <= 15641083;
srom_1(55807) <= 15335577;
srom_1(55808) <= 14997493;
srom_1(55809) <= 14628418;
srom_1(55810) <= 14230083;
srom_1(55811) <= 13804355;
srom_1(55812) <= 13353231;
srom_1(55813) <= 12878826;
srom_1(55814) <= 12383364;
srom_1(55815) <= 11869170;
srom_1(55816) <= 11338654;
srom_1(55817) <= 10794305;
srom_1(55818) <= 10238674;
srom_1(55819) <= 9674368;
srom_1(55820) <= 9104032;
srom_1(55821) <= 8530342;
srom_1(55822) <= 7955987;
srom_1(55823) <= 7383660;
srom_1(55824) <= 6816046;
srom_1(55825) <= 6255807;
srom_1(55826) <= 5705569;
srom_1(55827) <= 5167912;
srom_1(55828) <= 4645359;
srom_1(55829) <= 4140358;
srom_1(55830) <= 3655280;
srom_1(55831) <= 3192397;
srom_1(55832) <= 2753881;
srom_1(55833) <= 2341789;
srom_1(55834) <= 1958052;
srom_1(55835) <= 1604470;
srom_1(55836) <= 1282701;
srom_1(55837) <= 994255;
srom_1(55838) <= 740483;
srom_1(55839) <= 522575;
srom_1(55840) <= 341555;
srom_1(55841) <= 198269;
srom_1(55842) <= 93391;
srom_1(55843) <= 27412;
srom_1(55844) <= 642;
srom_1(55845) <= 13205;
srom_1(55846) <= 65044;
srom_1(55847) <= 155915;
srom_1(55848) <= 285391;
srom_1(55849) <= 452867;
srom_1(55850) <= 657556;
srom_1(55851) <= 898498;
srom_1(55852) <= 1174564;
srom_1(55853) <= 1484459;
srom_1(55854) <= 1826730;
srom_1(55855) <= 2199772;
srom_1(55856) <= 2601836;
srom_1(55857) <= 3031036;
srom_1(55858) <= 3485359;
srom_1(55859) <= 3962675;
srom_1(55860) <= 4460746;
srom_1(55861) <= 4977236;
srom_1(55862) <= 5509723;
srom_1(55863) <= 6055711;
srom_1(55864) <= 6612637;
srom_1(55865) <= 7177893;
srom_1(55866) <= 7748825;
srom_1(55867) <= 8322758;
srom_1(55868) <= 8896999;
srom_1(55869) <= 9468857;
srom_1(55870) <= 10035648;
srom_1(55871) <= 10594717;
srom_1(55872) <= 11143440;
srom_1(55873) <= 11679244;
srom_1(55874) <= 12199618;
srom_1(55875) <= 12702121;
srom_1(55876) <= 13184396;
srom_1(55877) <= 13644182;
srom_1(55878) <= 14079322;
srom_1(55879) <= 14487778;
srom_1(55880) <= 14867631;
srom_1(55881) <= 15217103;
srom_1(55882) <= 15534553;
srom_1(55883) <= 15818494;
srom_1(55884) <= 16067593;
srom_1(55885) <= 16280683;
srom_1(55886) <= 16456764;
srom_1(55887) <= 16595011;
srom_1(55888) <= 16694775;
srom_1(55889) <= 16755589;
srom_1(55890) <= 16777167;
srom_1(55891) <= 16759408;
srom_1(55892) <= 16702396;
srom_1(55893) <= 16606397;
srom_1(55894) <= 16471863;
srom_1(55895) <= 16299423;
srom_1(55896) <= 16089887;
srom_1(55897) <= 15844236;
srom_1(55898) <= 15563624;
srom_1(55899) <= 15249366;
srom_1(55900) <= 14902935;
srom_1(55901) <= 14525956;
srom_1(55902) <= 14120197;
srom_1(55903) <= 13687561;
srom_1(55904) <= 13230076;
srom_1(55905) <= 12749888;
srom_1(55906) <= 12249248;
srom_1(55907) <= 11730504;
srom_1(55908) <= 11196089;
srom_1(55909) <= 10648509;
srom_1(55910) <= 10090331;
srom_1(55911) <= 9524174;
srom_1(55912) <= 8952691;
srom_1(55913) <= 8378563;
srom_1(55914) <= 7804482;
srom_1(55915) <= 7233141;
srom_1(55916) <= 6667217;
srom_1(55917) <= 6109366;
srom_1(55918) <= 5562203;
srom_1(55919) <= 5028294;
srom_1(55920) <= 4510143;
srom_1(55921) <= 4010179;
srom_1(55922) <= 3530747;
srom_1(55923) <= 3074096;
srom_1(55924) <= 2642365;
srom_1(55925) <= 2237581;
srom_1(55926) <= 1861641;
srom_1(55927) <= 1516309;
srom_1(55928) <= 1203203;
srom_1(55929) <= 923792;
srom_1(55930) <= 679385;
srom_1(55931) <= 471130;
srom_1(55932) <= 300003;
srom_1(55933) <= 166806;
srom_1(55934) <= 72164;
srom_1(55935) <= 16521;
srom_1(55936) <= 137;
srom_1(55937) <= 23089;
srom_1(55938) <= 85271;
srom_1(55939) <= 186389;
srom_1(55940) <= 325971;
srom_1(55941) <= 503361;
srom_1(55942) <= 717727;
srom_1(55943) <= 968065;
srom_1(55944) <= 1253201;
srom_1(55945) <= 1571797;
srom_1(55946) <= 1922359;
srom_1(55947) <= 2303244;
srom_1(55948) <= 2712665;
srom_1(55949) <= 3148702;
srom_1(55950) <= 3609311;
srom_1(55951) <= 4092332;
srom_1(55952) <= 4595500;
srom_1(55953) <= 5116455;
srom_1(55954) <= 5652754;
srom_1(55955) <= 6201882;
srom_1(55956) <= 6761265;
srom_1(55957) <= 7328279;
srom_1(55958) <= 7900265;
srom_1(55959) <= 8474541;
srom_1(55960) <= 9048414;
srom_1(55961) <= 9619193;
srom_1(55962) <= 10184202;
srom_1(55963) <= 10740790;
srom_1(55964) <= 11286348;
srom_1(55965) <= 11818318;
srom_1(55966) <= 12334204;
srom_1(55967) <= 12831588;
srom_1(55968) <= 13308138;
srom_1(55969) <= 13761618;
srom_1(55970) <= 14189902;
srom_1(55971) <= 14590982;
srom_1(55972) <= 14962977;
srom_1(55973) <= 15304143;
srom_1(55974) <= 15612879;
srom_1(55975) <= 15887738;
srom_1(55976) <= 16127431;
srom_1(55977) <= 16330834;
srom_1(55978) <= 16496993;
srom_1(55979) <= 16625129;
srom_1(55980) <= 16714642;
srom_1(55981) <= 16765110;
srom_1(55982) <= 16776299;
srom_1(55983) <= 16748154;
srom_1(55984) <= 16680809;
srom_1(55985) <= 16574579;
srom_1(55986) <= 16429962;
srom_1(55987) <= 16247636;
srom_1(55988) <= 16028457;
srom_1(55989) <= 15773452;
srom_1(55990) <= 15483816;
srom_1(55991) <= 15160909;
srom_1(55992) <= 14806244;
srom_1(55993) <= 14421485;
srom_1(55994) <= 14008435;
srom_1(55995) <= 13569032;
srom_1(55996) <= 13105336;
srom_1(55997) <= 12619522;
srom_1(55998) <= 12113868;
srom_1(55999) <= 11590745;
srom_1(56000) <= 11052605;
srom_1(56001) <= 10501974;
srom_1(56002) <= 9941432;
srom_1(56003) <= 9373608;
srom_1(56004) <= 8801165;
srom_1(56005) <= 8226788;
srom_1(56006) <= 7653169;
srom_1(56007) <= 7082999;
srom_1(56008) <= 6518952;
srom_1(56009) <= 5963672;
srom_1(56010) <= 5419764;
srom_1(56011) <= 4889777;
srom_1(56012) <= 4376197;
srom_1(56013) <= 3881434;
srom_1(56014) <= 3407805;
srom_1(56015) <= 2957534;
srom_1(56016) <= 2532731;
srom_1(56017) <= 2135387;
srom_1(56018) <= 1767368;
srom_1(56019) <= 1430397;
srom_1(56020) <= 1126057;
srom_1(56021) <= 855772;
srom_1(56022) <= 620812;
srom_1(56023) <= 422277;
srom_1(56024) <= 261100;
srom_1(56025) <= 138035;
srom_1(56026) <= 53660;
srom_1(56027) <= 8370;
srom_1(56028) <= 2378;
srom_1(56029) <= 35712;
srom_1(56030) <= 108216;
srom_1(56031) <= 219549;
srom_1(56032) <= 369190;
srom_1(56033) <= 556436;
srom_1(56034) <= 780410;
srom_1(56035) <= 1040062;
srom_1(56036) <= 1334174;
srom_1(56037) <= 1661366;
srom_1(56038) <= 2020104;
srom_1(56039) <= 2408707;
srom_1(56040) <= 2825351;
srom_1(56041) <= 3268084;
srom_1(56042) <= 3734828;
srom_1(56043) <= 4223396;
srom_1(56044) <= 4731495;
srom_1(56045) <= 5256744;
srom_1(56046) <= 5796680;
srom_1(56047) <= 6348770;
srom_1(56048) <= 6910425;
srom_1(56049) <= 7479012;
srom_1(56050) <= 8051865;
srom_1(56051) <= 8626296;
srom_1(56052) <= 9199613;
srom_1(56053) <= 9769127;
srom_1(56054) <= 10332167;
srom_1(56055) <= 10886093;
srom_1(56056) <= 11428308;
srom_1(56057) <= 11956268;
srom_1(56058) <= 12467498;
srom_1(56059) <= 12959601;
srom_1(56060) <= 13430269;
srom_1(56061) <= 13877295;
srom_1(56062) <= 14298583;
srom_1(56063) <= 14692157;
srom_1(56064) <= 15056171;
srom_1(56065) <= 15388919;
srom_1(56066) <= 15688839;
srom_1(56067) <= 15954527;
srom_1(56068) <= 16184735;
srom_1(56069) <= 16378385;
srom_1(56070) <= 16534568;
srom_1(56071) <= 16652551;
srom_1(56072) <= 16731782;
srom_1(56073) <= 16771889;
srom_1(56074) <= 16772684;
srom_1(56075) <= 16734164;
srom_1(56076) <= 16656508;
srom_1(56077) <= 16540080;
srom_1(56078) <= 16385428;
srom_1(56079) <= 16193276;
srom_1(56080) <= 15964526;
srom_1(56081) <= 15700249;
srom_1(56082) <= 15401685;
srom_1(56083) <= 15070235;
srom_1(56084) <= 14707452;
srom_1(56085) <= 14315038;
srom_1(56086) <= 13894833;
srom_1(56087) <= 13448807;
srom_1(56088) <= 12979052;
srom_1(56089) <= 12487771;
srom_1(56090) <= 11977268;
srom_1(56091) <= 11449936;
srom_1(56092) <= 10908249;
srom_1(56093) <= 10354746;
srom_1(56094) <= 9792023;
srom_1(56095) <= 9222719;
srom_1(56096) <= 8649504;
srom_1(56097) <= 8075065;
srom_1(56098) <= 7502097;
srom_1(56099) <= 6933286;
srom_1(56100) <= 6371299;
srom_1(56101) <= 5818772;
srom_1(56102) <= 5278296;
srom_1(56103) <= 4752405;
srom_1(56104) <= 4243566;
srom_1(56105) <= 3754164;
srom_1(56106) <= 3286494;
srom_1(56107) <= 2842750;
srom_1(56108) <= 2425013;
srom_1(56109) <= 2035241;
srom_1(56110) <= 1675262;
srom_1(56111) <= 1346764;
srom_1(56112) <= 1051288;
srom_1(56113) <= 790219;
srom_1(56114) <= 564782;
srom_1(56115) <= 376033;
srom_1(56116) <= 224857;
srom_1(56117) <= 111965;
srom_1(56118) <= 37884;
srom_1(56119) <= 2963;
srom_1(56120) <= 7365;
srom_1(56121) <= 51070;
srom_1(56122) <= 133872;
srom_1(56123) <= 255383;
srom_1(56124) <= 415034;
srom_1(56125) <= 612076;
srom_1(56126) <= 845584;
srom_1(56127) <= 1114465;
srom_1(56128) <= 1417456;
srom_1(56129) <= 1753137;
srom_1(56130) <= 2119935;
srom_1(56131) <= 2516128;
srom_1(56132) <= 2939860;
srom_1(56133) <= 3389142;
srom_1(56134) <= 3861869;
srom_1(56135) <= 4355823;
srom_1(56136) <= 4868688;
srom_1(56137) <= 5398059;
srom_1(56138) <= 5941454;
srom_1(56139) <= 6496325;
srom_1(56140) <= 7060069;
srom_1(56141) <= 7630043;
srom_1(56142) <= 8203575;
srom_1(56143) <= 8777973;
srom_1(56144) <= 9350546;
srom_1(56145) <= 9918609;
srom_1(56146) <= 10479496;
srom_1(56147) <= 11030579;
srom_1(56148) <= 11569272;
srom_1(56149) <= 12093050;
srom_1(56150) <= 12599457;
srom_1(56151) <= 13086118;
srom_1(56152) <= 13550750;
srom_1(56153) <= 13991176;
srom_1(56154) <= 14405329;
srom_1(56155) <= 14791267;
srom_1(56156) <= 15147182;
srom_1(56157) <= 15471403;
srom_1(56158) <= 15762410;
srom_1(56159) <= 16018839;
srom_1(56160) <= 16239487;
srom_1(56161) <= 16423320;
srom_1(56162) <= 16569475;
srom_1(56163) <= 16677267;
srom_1(56164) <= 16746191;
srom_1(56165) <= 16775924;
srom_1(56166) <= 16766325;
srom_1(56167) <= 16717440;
srom_1(56168) <= 16629499;
srom_1(56169) <= 16502913;
srom_1(56170) <= 16338277;
srom_1(56171) <= 16136361;
srom_1(56172) <= 15898114;
srom_1(56173) <= 15624652;
srom_1(56174) <= 15317258;
srom_1(56175) <= 14977373;
srom_1(56176) <= 14606591;
srom_1(56177) <= 14206651;
srom_1(56178) <= 13779428;
srom_1(56179) <= 13326925;
srom_1(56180) <= 12851266;
srom_1(56181) <= 12354679;
srom_1(56182) <= 11839494;
srom_1(56183) <= 11308126;
srom_1(56184) <= 10763068;
srom_1(56185) <= 10206875;
srom_1(56186) <= 9642156;
srom_1(56187) <= 9071558;
srom_1(56188) <= 8497758;
srom_1(56189) <= 7923446;
srom_1(56190) <= 7351315;
srom_1(56191) <= 6784048;
srom_1(56192) <= 6224306;
srom_1(56193) <= 5674713;
srom_1(56194) <= 5137846;
srom_1(56195) <= 4616223;
srom_1(56196) <= 4112291;
srom_1(56197) <= 3628411;
srom_1(56198) <= 3166853;
srom_1(56199) <= 2729783;
srom_1(56200) <= 2319248;
srom_1(56201) <= 1937174;
srom_1(56202) <= 1585354;
srom_1(56203) <= 1265436;
srom_1(56204) <= 978922;
srom_1(56205) <= 727154;
srom_1(56206) <= 511313;
srom_1(56207) <= 332411;
srom_1(56208) <= 191288;
srom_1(56209) <= 88605;
srom_1(56210) <= 24843;
srom_1(56211) <= 302;
srom_1(56212) <= 15096;
srom_1(56213) <= 69157;
srom_1(56214) <= 162231;
srom_1(56215) <= 293880;
srom_1(56216) <= 463489;
srom_1(56217) <= 670262;
srom_1(56218) <= 913228;
srom_1(56219) <= 1191249;
srom_1(56220) <= 1503021;
srom_1(56221) <= 1847081;
srom_1(56222) <= 2221818;
srom_1(56223) <= 2625472;
srom_1(56224) <= 3056152;
srom_1(56225) <= 3511837;
srom_1(56226) <= 3990391;
srom_1(56227) <= 4489570;
srom_1(56228) <= 5007033;
srom_1(56229) <= 5540354;
srom_1(56230) <= 6087030;
srom_1(56231) <= 6644500;
srom_1(56232) <= 7210148;
srom_1(56233) <= 7781323;
srom_1(56234) <= 8355345;
srom_1(56235) <= 8929523;
srom_1(56236) <= 9501165;
srom_1(56237) <= 10067589;
srom_1(56238) <= 10626141;
srom_1(56239) <= 11174199;
srom_1(56240) <= 11709195;
srom_1(56241) <= 12228620;
srom_1(56242) <= 12730038;
srom_1(56243) <= 13211097;
srom_1(56244) <= 13669541;
srom_1(56245) <= 14103222;
srom_1(56246) <= 14510105;
srom_1(56247) <= 14888282;
srom_1(56248) <= 15235980;
srom_1(56249) <= 15551568;
srom_1(56250) <= 15833566;
srom_1(56251) <= 16080653;
srom_1(56252) <= 16291669;
srom_1(56253) <= 16465624;
srom_1(56254) <= 16601704;
srom_1(56255) <= 16699270;
srom_1(56256) <= 16757864;
srom_1(56257) <= 16777212;
srom_1(56258) <= 16757223;
srom_1(56259) <= 16697991;
srom_1(56260) <= 16599793;
srom_1(56261) <= 16463089;
srom_1(56262) <= 16288522;
srom_1(56263) <= 16076910;
srom_1(56264) <= 15829244;
srom_1(56265) <= 15546687;
srom_1(56266) <= 15230563;
srom_1(56267) <= 14882354;
srom_1(56268) <= 14503695;
srom_1(56269) <= 14096359;
srom_1(56270) <= 13662258;
srom_1(56271) <= 13203427;
srom_1(56272) <= 12722018;
srom_1(56273) <= 12220287;
srom_1(56274) <= 11700589;
srom_1(56275) <= 11165360;
srom_1(56276) <= 10617109;
srom_1(56277) <= 10058408;
srom_1(56278) <= 9491877;
srom_1(56279) <= 8920173;
srom_1(56280) <= 8345976;
srom_1(56281) <= 7771978;
srom_1(56282) <= 7200872;
srom_1(56283) <= 6635336;
srom_1(56284) <= 6078022;
srom_1(56285) <= 5531542;
srom_1(56286) <= 4998461;
srom_1(56287) <= 4481277;
srom_1(56288) <= 3982416;
srom_1(56289) <= 3504217;
srom_1(56290) <= 3048922;
srom_1(56291) <= 2618667;
srom_1(56292) <= 2215470;
srom_1(56293) <= 1841220;
srom_1(56294) <= 1497673;
srom_1(56295) <= 1186441;
srom_1(56296) <= 908981;
srom_1(56297) <= 666596;
srom_1(56298) <= 460423;
srom_1(56299) <= 291427;
srom_1(56300) <= 160402;
srom_1(56301) <= 67962;
srom_1(56302) <= 14540;
srom_1(56303) <= 386;
srom_1(56304) <= 25569;
srom_1(56305) <= 89968;
srom_1(56306) <= 193282;
srom_1(56307) <= 335028;
srom_1(56308) <= 514539;
srom_1(56309) <= 730974;
srom_1(56310) <= 983319;
srom_1(56311) <= 1270389;
srom_1(56312) <= 1590840;
srom_1(56313) <= 1943167;
srom_1(56314) <= 2325719;
srom_1(56315) <= 2736703;
srom_1(56316) <= 3174190;
srom_1(56317) <= 3636129;
srom_1(56318) <= 4120354;
srom_1(56319) <= 4624594;
srom_1(56320) <= 5146486;
srom_1(56321) <= 5683580;
srom_1(56322) <= 6233360;
srom_1(56323) <= 6793246;
srom_1(56324) <= 7360613;
srom_1(56325) <= 7932801;
srom_1(56326) <= 8507126;
srom_1(56327) <= 9080896;
srom_1(56328) <= 9651419;
srom_1(56329) <= 10216021;
srom_1(56330) <= 10772053;
srom_1(56331) <= 11316908;
srom_1(56332) <= 11848031;
srom_1(56333) <= 12362932;
srom_1(56334) <= 12859196;
srom_1(56335) <= 13334496;
srom_1(56336) <= 13786603;
srom_1(56337) <= 14213397;
srom_1(56338) <= 14612877;
srom_1(56339) <= 14983168;
srom_1(56340) <= 15322536;
srom_1(56341) <= 15629388;
srom_1(56342) <= 15902285;
srom_1(56343) <= 16139948;
srom_1(56344) <= 16341263;
srom_1(56345) <= 16505285;
srom_1(56346) <= 16631244;
srom_1(56347) <= 16718552;
srom_1(56348) <= 16766797;
srom_1(56349) <= 16775754;
srom_1(56350) <= 16745381;
srom_1(56351) <= 16675820;
srom_1(56352) <= 16567398;
srom_1(56353) <= 16420622;
srom_1(56354) <= 16236182;
srom_1(56355) <= 16014941;
srom_1(56356) <= 15757938;
srom_1(56357) <= 15466378;
srom_1(56358) <= 15141627;
srom_1(56359) <= 14785210;
srom_1(56360) <= 14398796;
srom_1(56361) <= 13984199;
srom_1(56362) <= 13543362;
srom_1(56363) <= 13078352;
srom_1(56364) <= 12591351;
srom_1(56365) <= 12084642;
srom_1(56366) <= 11560600;
srom_1(56367) <= 11021684;
srom_1(56368) <= 10470421;
srom_1(56369) <= 9909395;
srom_1(56370) <= 9341238;
srom_1(56371) <= 8768614;
srom_1(56372) <= 8194207;
srom_1(56373) <= 7620713;
srom_1(56374) <= 7050819;
srom_1(56375) <= 6487198;
srom_1(56376) <= 5932494;
srom_1(56377) <= 5389307;
srom_1(56378) <= 4860186;
srom_1(56379) <= 4347610;
srom_1(56380) <= 3853983;
srom_1(56381) <= 3381621;
srom_1(56382) <= 2932739;
srom_1(56383) <= 2509441;
srom_1(56384) <= 2113713;
srom_1(56385) <= 1747409;
srom_1(56386) <= 1412249;
srom_1(56387) <= 1109803;
srom_1(56388) <= 841490;
srom_1(56389) <= 608567;
srom_1(56390) <= 412128;
srom_1(56391) <= 253094;
srom_1(56392) <= 132210;
srom_1(56393) <= 50043;
srom_1(56394) <= 6978;
srom_1(56395) <= 3218;
srom_1(56396) <= 38779;
srom_1(56397) <= 113496;
srom_1(56398) <= 227017;
srom_1(56399) <= 378812;
srom_1(56400) <= 568166;
srom_1(56401) <= 794194;
srom_1(56402) <= 1055834;
srom_1(56403) <= 1351860;
srom_1(56404) <= 1680884;
srom_1(56405) <= 2041363;
srom_1(56406) <= 2431606;
srom_1(56407) <= 2849784;
srom_1(56408) <= 3293935;
srom_1(56409) <= 3761976;
srom_1(56410) <= 4251714;
srom_1(56411) <= 4760851;
srom_1(56412) <= 5286999;
srom_1(56413) <= 5827693;
srom_1(56414) <= 6380395;
srom_1(56415) <= 6942514;
srom_1(56416) <= 7511415;
srom_1(56417) <= 8084429;
srom_1(56418) <= 8658869;
srom_1(56419) <= 9232042;
srom_1(56420) <= 9801260;
srom_1(56421) <= 10363853;
srom_1(56422) <= 10917184;
srom_1(56423) <= 11458658;
srom_1(56424) <= 11985735;
srom_1(56425) <= 12495944;
srom_1(56426) <= 12986892;
srom_1(56427) <= 13456277;
srom_1(56428) <= 13901898;
srom_1(56429) <= 14321665;
srom_1(56430) <= 14713611;
srom_1(56431) <= 15075896;
srom_1(56432) <= 15406822;
srom_1(56433) <= 15704837;
srom_1(56434) <= 15968544;
srom_1(56435) <= 16196706;
srom_1(56436) <= 16388253;
srom_1(56437) <= 16542287;
srom_1(56438) <= 16658086;
srom_1(56439) <= 16735106;
srom_1(56440) <= 16772987;
srom_1(56441) <= 16771550;
srom_1(56442) <= 16730803;
srom_1(56443) <= 16650937;
srom_1(56444) <= 16532325;
srom_1(56445) <= 16375525;
srom_1(56446) <= 16181272;
srom_1(56447) <= 15950476;
srom_1(56448) <= 15684219;
srom_1(56449) <= 15383752;
srom_1(56450) <= 15050481;
srom_1(56451) <= 14685971;
srom_1(56452) <= 14291930;
srom_1(56453) <= 13870206;
srom_1(56454) <= 13422778;
srom_1(56455) <= 12951742;
srom_1(56456) <= 12459309;
srom_1(56457) <= 11947786;
srom_1(56458) <= 11419573;
srom_1(56459) <= 10877147;
srom_1(56460) <= 10323051;
srom_1(56461) <= 9759884;
srom_1(56462) <= 9190287;
srom_1(56463) <= 8616930;
srom_1(56464) <= 8042503;
srom_1(56465) <= 7469698;
srom_1(56466) <= 6901203;
srom_1(56467) <= 6339683;
srom_1(56468) <= 5787770;
srom_1(56469) <= 5248054;
srom_1(56470) <= 4723065;
srom_1(56471) <= 4215265;
srom_1(56472) <= 3727036;
srom_1(56473) <= 3260666;
srom_1(56474) <= 2818342;
srom_1(56475) <= 2402140;
srom_1(56476) <= 2014010;
srom_1(56477) <= 1655773;
srom_1(56478) <= 1329108;
srom_1(56479) <= 1035548;
srom_1(56480) <= 776469;
srom_1(56481) <= 553085;
srom_1(56482) <= 366446;
srom_1(56483) <= 217424;
srom_1(56484) <= 106721;
srom_1(56485) <= 34854;
srom_1(56486) <= 2160;
srom_1(56487) <= 8794;
srom_1(56488) <= 54723;
srom_1(56489) <= 139733;
srom_1(56490) <= 263424;
srom_1(56491) <= 425218;
srom_1(56492) <= 624354;
srom_1(56493) <= 859900;
srom_1(56494) <= 1130750;
srom_1(56495) <= 1435635;
srom_1(56496) <= 1773125;
srom_1(56497) <= 2141637;
srom_1(56498) <= 2539443;
srom_1(56499) <= 2964678;
srom_1(56500) <= 3415348;
srom_1(56501) <= 3889339;
srom_1(56502) <= 4384428;
srom_1(56503) <= 4898295;
srom_1(56504) <= 5428529;
srom_1(56505) <= 5972643;
srom_1(56506) <= 6528087;
srom_1(56507) <= 7092256;
srom_1(56508) <= 7662503;
srom_1(56509) <= 8236156;
srom_1(56510) <= 8810523;
srom_1(56511) <= 9382912;
srom_1(56512) <= 9950638;
srom_1(56513) <= 10511040;
srom_1(56514) <= 11061488;
srom_1(56515) <= 11599403;
srom_1(56516) <= 12122261;
srom_1(56517) <= 12627610;
srom_1(56518) <= 13113082;
srom_1(56519) <= 13576398;
srom_1(56520) <= 14015388;
srom_1(56521) <= 14427991;
srom_1(56522) <= 14812274;
srom_1(56523) <= 15166434;
srom_1(56524) <= 15488810;
srom_1(56525) <= 15777891;
srom_1(56526) <= 16032321;
srom_1(56527) <= 16250908;
srom_1(56528) <= 16432625;
srom_1(56529) <= 16576621;
srom_1(56530) <= 16682220;
srom_1(56531) <= 16748928;
srom_1(56532) <= 16776432;
srom_1(56533) <= 16764602;
srom_1(56534) <= 16713494;
srom_1(56535) <= 16623348;
srom_1(56536) <= 16494587;
srom_1(56537) <= 16327813;
srom_1(56538) <= 16123810;
srom_1(56539) <= 15883535;
srom_1(56540) <= 15608112;
srom_1(56541) <= 15298835;
srom_1(56542) <= 14957154;
srom_1(56543) <= 14584670;
srom_1(56544) <= 14183131;
srom_1(56545) <= 13754419;
srom_1(56546) <= 13300546;
srom_1(56547) <= 12823638;
srom_1(56548) <= 12325933;
srom_1(56549) <= 11809765;
srom_1(56550) <= 11277553;
srom_1(56551) <= 10731795;
srom_1(56552) <= 10175048;
srom_1(56553) <= 9609924;
srom_1(56554) <= 9039073;
srom_1(56555) <= 8465172;
srom_1(56556) <= 7890912;
srom_1(56557) <= 7318985;
srom_1(56558) <= 6752074;
srom_1(56559) <= 6192838;
srom_1(56560) <= 5643898;
srom_1(56561) <= 5107829;
srom_1(56562) <= 4587145;
srom_1(56563) <= 4084287;
srom_1(56564) <= 3601614;
srom_1(56565) <= 3141389;
srom_1(56566) <= 2705769;
srom_1(56567) <= 2296798;
srom_1(56568) <= 1916394;
srom_1(56569) <= 1566340;
srom_1(56570) <= 1248279;
srom_1(56571) <= 963700;
srom_1(56572) <= 713940;
srom_1(56573) <= 500169;
srom_1(56574) <= 323389;
srom_1(56575) <= 184430;
srom_1(56576) <= 83943;
srom_1(56577) <= 22400;
srom_1(56578) <= 88;
srom_1(56579) <= 17114;
srom_1(56580) <= 73396;
srom_1(56581) <= 168671;
srom_1(56582) <= 302492;
srom_1(56583) <= 474231;
srom_1(56584) <= 683084;
srom_1(56585) <= 928071;
srom_1(56586) <= 1208042;
srom_1(56587) <= 1521686;
srom_1(56588) <= 1867531;
srom_1(56589) <= 2243956;
srom_1(56590) <= 2649195;
srom_1(56591) <= 3081348;
srom_1(56592) <= 3538389;
srom_1(56593) <= 4018174;
srom_1(56594) <= 4518454;
srom_1(56595) <= 5036882;
srom_1(56596) <= 5571027;
srom_1(56597) <= 6118385;
srom_1(56598) <= 6676389;
srom_1(56599) <= 7242422;
srom_1(56600) <= 7813830;
srom_1(56601) <= 8387933;
srom_1(56602) <= 8962039;
srom_1(56603) <= 9533456;
srom_1(56604) <= 10099505;
srom_1(56605) <= 10657531;
srom_1(56606) <= 11204917;
srom_1(56607) <= 11739096;
srom_1(56608) <= 12257564;
srom_1(56609) <= 12757889;
srom_1(56610) <= 13237725;
srom_1(56611) <= 13694821;
srom_1(56612) <= 14127035;
srom_1(56613) <= 14532340;
srom_1(56614) <= 14908834;
srom_1(56615) <= 15254753;
srom_1(56616) <= 15568474;
srom_1(56617) <= 15848526;
srom_1(56618) <= 16093596;
srom_1(56619) <= 16302535;
srom_1(56620) <= 16474363;
srom_1(56621) <= 16608273;
srom_1(56622) <= 16703639;
srom_1(56623) <= 16760013;
srom_1(56624) <= 16777131;
srom_1(56625) <= 16754911;
srom_1(56626) <= 16693460;
srom_1(56627) <= 16593064;
srom_1(56628) <= 16454194;
srom_1(56629) <= 16277502;
srom_1(56630) <= 16063817;
srom_1(56631) <= 15814140;
srom_1(56632) <= 15529641;
srom_1(56633) <= 15211657;
srom_1(56634) <= 14861676;
srom_1(56635) <= 14481341;
srom_1(56636) <= 14072435;
srom_1(56637) <= 13636876;
srom_1(56638) <= 13176705;
srom_1(56639) <= 12694082;
srom_1(56640) <= 12191269;
srom_1(56641) <= 11670624;
srom_1(56642) <= 11134588;
srom_1(56643) <= 10585676;
srom_1(56644) <= 10026460;
srom_1(56645) <= 9459564;
srom_1(56646) <= 8887647;
srom_1(56647) <= 8313389;
srom_1(56648) <= 7739483;
srom_1(56649) <= 7168622;
srom_1(56650) <= 6603481;
srom_1(56651) <= 6046712;
srom_1(56652) <= 5500925;
srom_1(56653) <= 4968679;
srom_1(56654) <= 4452470;
srom_1(56655) <= 3954719;
srom_1(56656) <= 3477760;
srom_1(56657) <= 3023829;
srom_1(56658) <= 2595056;
srom_1(56659) <= 2193451;
srom_1(56660) <= 1820897;
srom_1(56661) <= 1479142;
srom_1(56662) <= 1169787;
srom_1(56663) <= 894284;
srom_1(56664) <= 653924;
srom_1(56665) <= 449835;
srom_1(56666) <= 282973;
srom_1(56667) <= 154122;
srom_1(56668) <= 63885;
srom_1(56669) <= 12685;
srom_1(56670) <= 763;
srom_1(56671) <= 28174;
srom_1(56672) <= 94791;
srom_1(56673) <= 200299;
srom_1(56674) <= 344206;
srom_1(56675) <= 525836;
srom_1(56676) <= 744337;
srom_1(56677) <= 998684;
srom_1(56678) <= 1287685;
srom_1(56679) <= 1609985;
srom_1(56680) <= 1964073;
srom_1(56681) <= 2348287;
srom_1(56682) <= 2760826;
srom_1(56683) <= 3199756;
srom_1(56684) <= 3663018;
srom_1(56685) <= 4148440;
srom_1(56686) <= 4653746;
srom_1(56687) <= 5176566;
srom_1(56688) <= 5714448;
srom_1(56689) <= 6264870;
srom_1(56690) <= 6825251;
srom_1(56691) <= 7392963;
srom_1(56692) <= 7965344;
srom_1(56693) <= 8539710;
srom_1(56694) <= 9113367;
srom_1(56695) <= 9683626;
srom_1(56696) <= 10247812;
srom_1(56697) <= 10803279;
srom_1(56698) <= 11347424;
srom_1(56699) <= 11877693;
srom_1(56700) <= 12391601;
srom_1(56701) <= 12886737;
srom_1(56702) <= 13360780;
srom_1(56703) <= 13811507;
srom_1(56704) <= 14236804;
srom_1(56705) <= 14634677;
srom_1(56706) <= 15003260;
srom_1(56707) <= 15340824;
srom_1(56708) <= 15645787;
srom_1(56709) <= 15916719;
srom_1(56710) <= 16152349;
srom_1(56711) <= 16351572;
srom_1(56712) <= 16513453;
srom_1(56713) <= 16637235;
srom_1(56714) <= 16722336;
srom_1(56715) <= 16768357;
srom_1(56716) <= 16775083;
srom_1(56717) <= 16742482;
srom_1(56718) <= 16670706;
srom_1(56719) <= 16560093;
srom_1(56720) <= 16411161;
srom_1(56721) <= 16224609;
srom_1(56722) <= 16001310;
srom_1(56723) <= 15742314;
srom_1(56724) <= 15448833;
srom_1(56725) <= 15122244;
srom_1(56726) <= 14764079;
srom_1(56727) <= 14376017;
srom_1(56728) <= 13959878;
srom_1(56729) <= 13517614;
srom_1(56730) <= 13051298;
srom_1(56731) <= 12563116;
srom_1(56732) <= 12055360;
srom_1(56733) <= 11530408;
srom_1(56734) <= 10990724;
srom_1(56735) <= 10438837;
srom_1(56736) <= 9877336;
srom_1(56737) <= 9308854;
srom_1(56738) <= 8736057;
srom_1(56739) <= 8161630;
srom_1(56740) <= 7588267;
srom_1(56741) <= 7018658;
srom_1(56742) <= 6455473;
srom_1(56743) <= 5901353;
srom_1(56744) <= 5358896;
srom_1(56745) <= 4830647;
srom_1(56746) <= 4319083;
srom_1(56747) <= 3826602;
srom_1(56748) <= 3355513;
srom_1(56749) <= 2908027;
srom_1(56750) <= 2486240;
srom_1(56751) <= 2092132;
srom_1(56752) <= 1727551;
srom_1(56753) <= 1394205;
srom_1(56754) <= 1093659;
srom_1(56755) <= 827321;
srom_1(56756) <= 596440;
srom_1(56757) <= 402100;
srom_1(56758) <= 245211;
srom_1(56759) <= 126509;
srom_1(56760) <= 46551;
srom_1(56761) <= 5712;
srom_1(56762) <= 4183;
srom_1(56763) <= 41972;
srom_1(56764) <= 118901;
srom_1(56765) <= 234609;
srom_1(56766) <= 388554;
srom_1(56767) <= 580014;
srom_1(56768) <= 808092;
srom_1(56769) <= 1071717;
srom_1(56770) <= 1369653;
srom_1(56771) <= 1700504;
srom_1(56772) <= 2062717;
srom_1(56773) <= 2454595;
srom_1(56774) <= 2874300;
srom_1(56775) <= 3319862;
srom_1(56776) <= 3789194;
srom_1(56777) <= 4280095;
srom_1(56778) <= 4790261;
srom_1(56779) <= 5317301;
srom_1(56780) <= 5858744;
srom_1(56781) <= 6412050;
srom_1(56782) <= 6974625;
srom_1(56783) <= 7543830;
srom_1(56784) <= 8116997;
srom_1(56785) <= 8691438;
srom_1(56786) <= 9264458;
srom_1(56787) <= 9833372;
srom_1(56788) <= 10395510;
srom_1(56789) <= 10948237;
srom_1(56790) <= 11488962;
srom_1(56791) <= 12015147;
srom_1(56792) <= 12524327;
srom_1(56793) <= 13014113;
srom_1(56794) <= 13482208;
srom_1(56795) <= 13926417;
srom_1(56796) <= 14344658;
srom_1(56797) <= 14734969;
srom_1(56798) <= 15095520;
srom_1(56799) <= 15424619;
srom_1(56800) <= 15720724;
srom_1(56801) <= 15982447;
srom_1(56802) <= 16208559;
srom_1(56803) <= 16398001;
srom_1(56804) <= 16549884;
srom_1(56805) <= 16663496;
srom_1(56806) <= 16738304;
srom_1(56807) <= 16773958;
srom_1(56808) <= 16770290;
srom_1(56809) <= 16727317;
srom_1(56810) <= 16645241;
srom_1(56811) <= 16524447;
srom_1(56812) <= 16365502;
srom_1(56813) <= 16169149;
srom_1(56814) <= 15936312;
srom_1(56815) <= 15668080;
srom_1(56816) <= 15365712;
srom_1(56817) <= 15030627;
srom_1(56818) <= 14664395;
srom_1(56819) <= 14268733;
srom_1(56820) <= 13845497;
srom_1(56821) <= 13396673;
srom_1(56822) <= 12924363;
srom_1(56823) <= 12430784;
srom_1(56824) <= 11918250;
srom_1(56825) <= 11389164;
srom_1(56826) <= 10846007;
srom_1(56827) <= 10291327;
srom_1(56828) <= 9727725;
srom_1(56829) <= 9157842;
srom_1(56830) <= 8584353;
srom_1(56831) <= 8009945;
srom_1(56832) <= 7437314;
srom_1(56833) <= 6869143;
srom_1(56834) <= 6308097;
srom_1(56835) <= 5756808;
srom_1(56836) <= 5217860;
srom_1(56837) <= 4693781;
srom_1(56838) <= 4187028;
srom_1(56839) <= 3699978;
srom_1(56840) <= 3234914;
srom_1(56841) <= 2794018;
srom_1(56842) <= 2379357;
srom_1(56843) <= 1992875;
srom_1(56844) <= 1636385;
srom_1(56845) <= 1311559;
srom_1(56846) <= 1019919;
srom_1(56847) <= 762833;
srom_1(56848) <= 541508;
srom_1(56849) <= 356980;
srom_1(56850) <= 210115;
srom_1(56851) <= 101602;
srom_1(56852) <= 31949;
srom_1(56853) <= 1484;
srom_1(56854) <= 10349;
srom_1(56855) <= 58502;
srom_1(56856) <= 145718;
srom_1(56857) <= 271588;
srom_1(56858) <= 435522;
srom_1(56859) <= 636750;
srom_1(56860) <= 874329;
srom_1(56861) <= 1147145;
srom_1(56862) <= 1453919;
srom_1(56863) <= 1793212;
srom_1(56864) <= 2163433;
srom_1(56865) <= 2562846;
srom_1(56866) <= 2989578;
srom_1(56867) <= 3441628;
srom_1(56868) <= 3916876;
srom_1(56869) <= 4413094;
srom_1(56870) <= 4927954;
srom_1(56871) <= 5459042;
srom_1(56872) <= 6003868;
srom_1(56873) <= 6559877;
srom_1(56874) <= 7124462;
srom_1(56875) <= 7694974;
srom_1(56876) <= 8268739;
srom_1(56877) <= 8843066;
srom_1(56878) <= 9415263;
srom_1(56879) <= 9982644;
srom_1(56880) <= 10542551;
srom_1(56881) <= 11092357;
srom_1(56882) <= 11629485;
srom_1(56883) <= 12151414;
srom_1(56884) <= 12655699;
srom_1(56885) <= 13139974;
srom_1(56886) <= 13601968;
srom_1(56887) <= 14039515;
srom_1(56888) <= 14450562;
srom_1(56889) <= 14833183;
srom_1(56890) <= 15185584;
srom_1(56891) <= 15506111;
srom_1(56892) <= 15793261;
srom_1(56893) <= 16045689;
srom_1(56894) <= 16262209;
srom_1(56895) <= 16441808;
srom_1(56896) <= 16583643;
srom_1(56897) <= 16687048;
srom_1(56898) <= 16751539;
srom_1(56899) <= 16776813;
srom_1(56900) <= 16762753;
srom_1(56901) <= 16709423;
srom_1(56902) <= 16617073;
srom_1(56903) <= 16486138;
srom_1(56904) <= 16317230;
srom_1(56905) <= 16111143;
srom_1(56906) <= 15868842;
srom_1(56907) <= 15591463;
srom_1(56908) <= 15280308;
srom_1(56909) <= 14936835;
srom_1(56910) <= 14562656;
srom_1(56911) <= 14159524;
srom_1(56912) <= 13729330;
srom_1(56913) <= 13274092;
srom_1(56914) <= 12795944;
srom_1(56915) <= 12297128;
srom_1(56916) <= 11779985;
srom_1(56917) <= 11246937;
srom_1(56918) <= 10700487;
srom_1(56919) <= 10143195;
srom_1(56920) <= 9577675;
srom_1(56921) <= 9006579;
srom_1(56922) <= 8432585;
srom_1(56923) <= 7858385;
srom_1(56924) <= 7286671;
srom_1(56925) <= 6720125;
srom_1(56926) <= 6161403;
srom_1(56927) <= 5613125;
srom_1(56928) <= 5077862;
srom_1(56929) <= 4558124;
srom_1(56930) <= 4056349;
srom_1(56931) <= 3574889;
srom_1(56932) <= 3116003;
srom_1(56933) <= 2681841;
srom_1(56934) <= 2274441;
srom_1(56935) <= 1895712;
srom_1(56936) <= 1547430;
srom_1(56937) <= 1231229;
srom_1(56938) <= 948591;
srom_1(56939) <= 700842;
srom_1(56940) <= 489144;
srom_1(56941) <= 314489;
srom_1(56942) <= 177696;
srom_1(56943) <= 79407;
srom_1(56944) <= 20083;
srom_1(56945) <= 2;
srom_1(56946) <= 19257;
srom_1(56947) <= 77760;
srom_1(56948) <= 175235;
srom_1(56949) <= 311225;
srom_1(56950) <= 485093;
srom_1(56951) <= 696023;
srom_1(56952) <= 943026;
srom_1(56953) <= 1224944;
srom_1(56954) <= 1540455;
srom_1(56955) <= 1888079;
srom_1(56956) <= 2266187;
srom_1(56957) <= 2673005;
srom_1(56958) <= 3106625;
srom_1(56959) <= 3565014;
srom_1(56960) <= 4046023;
srom_1(56961) <= 4547395;
srom_1(56962) <= 5066780;
srom_1(56963) <= 5601743;
srom_1(56964) <= 6149774;
srom_1(56965) <= 6708303;
srom_1(56966) <= 7274712;
srom_1(56967) <= 7846345;
srom_1(56968) <= 8420521;
srom_1(56969) <= 8994546;
srom_1(56970) <= 9565731;
srom_1(56971) <= 10131395;
srom_1(56972) <= 10688887;
srom_1(56973) <= 11235592;
srom_1(56974) <= 11768946;
srom_1(56975) <= 12286449;
srom_1(56976) <= 12785674;
srom_1(56977) <= 13264279;
srom_1(56978) <= 13720021;
srom_1(56979) <= 14150762;
srom_1(56980) <= 14554482;
srom_1(56981) <= 14929288;
srom_1(56982) <= 15273423;
srom_1(56983) <= 15585272;
srom_1(56984) <= 15863374;
srom_1(56985) <= 16106424;
srom_1(56986) <= 16313282;
srom_1(56987) <= 16482979;
srom_1(56988) <= 16614719;
srom_1(56989) <= 16707883;
srom_1(56990) <= 16762036;
srom_1(56991) <= 16776923;
srom_1(56992) <= 16752474;
srom_1(56993) <= 16688804;
srom_1(56994) <= 16586211;
srom_1(56995) <= 16445177;
srom_1(56996) <= 16266363;
srom_1(56997) <= 16050608;
srom_1(56998) <= 15798923;
srom_1(56999) <= 15512488;
srom_1(57000) <= 15192647;
srom_1(57001) <= 14840900;
srom_1(57002) <= 14458895;
srom_1(57003) <= 14048425;
srom_1(57004) <= 13611414;
srom_1(57005) <= 13149912;
srom_1(57006) <= 12666082;
srom_1(57007) <= 12162193;
srom_1(57008) <= 11640609;
srom_1(57009) <= 11103775;
srom_1(57010) <= 10554209;
srom_1(57011) <= 9994487;
srom_1(57012) <= 9427235;
srom_1(57013) <= 8855113;
srom_1(57014) <= 8280803;
srom_1(57015) <= 7706998;
srom_1(57016) <= 7136390;
srom_1(57017) <= 6571654;
srom_1(57018) <= 6015438;
srom_1(57019) <= 5470350;
srom_1(57020) <= 4938948;
srom_1(57021) <= 4423722;
srom_1(57022) <= 3927089;
srom_1(57023) <= 3451377;
srom_1(57024) <= 2998818;
srom_1(57025) <= 2571533;
srom_1(57026) <= 2171526;
srom_1(57027) <= 1800674;
srom_1(57028) <= 1460715;
srom_1(57029) <= 1153242;
srom_1(57030) <= 879699;
srom_1(57031) <= 641368;
srom_1(57032) <= 439367;
srom_1(57033) <= 274642;
srom_1(57034) <= 147966;
srom_1(57035) <= 59933;
srom_1(57036) <= 10957;
srom_1(57037) <= 1266;
srom_1(57038) <= 30906;
srom_1(57039) <= 99738;
srom_1(57040) <= 207440;
srom_1(57041) <= 353506;
srom_1(57042) <= 537251;
srom_1(57043) <= 757814;
srom_1(57044) <= 1014161;
srom_1(57045) <= 1305088;
srom_1(57046) <= 1629233;
srom_1(57047) <= 1985075;
srom_1(57048) <= 2370945;
srom_1(57049) <= 2785034;
srom_1(57050) <= 3225401;
srom_1(57051) <= 3689979;
srom_1(57052) <= 4176590;
srom_1(57053) <= 4682954;
srom_1(57054) <= 5206694;
srom_1(57055) <= 5745355;
srom_1(57056) <= 6296412;
srom_1(57057) <= 6857279;
srom_1(57058) <= 7425328;
srom_1(57059) <= 7997894;
srom_1(57060) <= 8572291;
srom_1(57061) <= 9145828;
srom_1(57062) <= 9715813;
srom_1(57063) <= 10279575;
srom_1(57064) <= 10834470;
srom_1(57065) <= 11377895;
srom_1(57066) <= 11907302;
srom_1(57067) <= 12420208;
srom_1(57068) <= 12914210;
srom_1(57069) <= 13386989;
srom_1(57070) <= 13836329;
srom_1(57071) <= 14260122;
srom_1(57072) <= 14656383;
srom_1(57073) <= 15023251;
srom_1(57074) <= 15359007;
srom_1(57075) <= 15662077;
srom_1(57076) <= 15931039;
srom_1(57077) <= 16164632;
srom_1(57078) <= 16361760;
srom_1(57079) <= 16521500;
srom_1(57080) <= 16643101;
srom_1(57081) <= 16725995;
srom_1(57082) <= 16769791;
srom_1(57083) <= 16774285;
srom_1(57084) <= 16739456;
srom_1(57085) <= 16665467;
srom_1(57086) <= 16552665;
srom_1(57087) <= 16401579;
srom_1(57088) <= 16212917;
srom_1(57089) <= 15987565;
srom_1(57090) <= 15726578;
srom_1(57091) <= 15431181;
srom_1(57092) <= 15102759;
srom_1(57093) <= 14742852;
srom_1(57094) <= 14353148;
srom_1(57095) <= 13935474;
srom_1(57096) <= 13491788;
srom_1(57097) <= 13024172;
srom_1(57098) <= 12534819;
srom_1(57099) <= 12026022;
srom_1(57100) <= 11500169;
srom_1(57101) <= 10959724;
srom_1(57102) <= 10407222;
srom_1(57103) <= 9845254;
srom_1(57104) <= 9276456;
srom_1(57105) <= 8703494;
srom_1(57106) <= 8129056;
srom_1(57107) <= 7555834;
srom_1(57108) <= 6986518;
srom_1(57109) <= 6423777;
srom_1(57110) <= 5870249;
srom_1(57111) <= 5328531;
srom_1(57112) <= 4801163;
srom_1(57113) <= 4290617;
srom_1(57114) <= 3799289;
srom_1(57115) <= 3329481;
srom_1(57116) <= 2883397;
srom_1(57117) <= 2463129;
srom_1(57118) <= 2070647;
srom_1(57119) <= 1707793;
srom_1(57120) <= 1376267;
srom_1(57121) <= 1077625;
srom_1(57122) <= 813266;
srom_1(57123) <= 584431;
srom_1(57124) <= 392192;
srom_1(57125) <= 237451;
srom_1(57126) <= 120933;
srom_1(57127) <= 43186;
srom_1(57128) <= 4573;
srom_1(57129) <= 5276;
srom_1(57130) <= 45291;
srom_1(57131) <= 124430;
srom_1(57132) <= 242324;
srom_1(57133) <= 398418;
srom_1(57134) <= 591980;
srom_1(57135) <= 822104;
srom_1(57136) <= 1087710;
srom_1(57137) <= 1387552;
srom_1(57138) <= 1720224;
srom_1(57139) <= 2084167;
srom_1(57140) <= 2477674;
srom_1(57141) <= 2898899;
srom_1(57142) <= 3345867;
srom_1(57143) <= 3816482;
srom_1(57144) <= 4308537;
srom_1(57145) <= 4819725;
srom_1(57146) <= 5347649;
srom_1(57147) <= 5889833;
srom_1(57148) <= 6443735;
srom_1(57149) <= 7006757;
srom_1(57150) <= 7576259;
srom_1(57151) <= 8149570;
srom_1(57152) <= 8724002;
srom_1(57153) <= 9296861;
srom_1(57154) <= 9865462;
srom_1(57155) <= 10427136;
srom_1(57156) <= 10979252;
srom_1(57157) <= 11519219;
srom_1(57158) <= 12044505;
srom_1(57159) <= 12552648;
srom_1(57160) <= 13041264;
srom_1(57161) <= 13508062;
srom_1(57162) <= 13950853;
srom_1(57163) <= 14367561;
srom_1(57164) <= 14756232;
srom_1(57165) <= 15115042;
srom_1(57166) <= 15442310;
srom_1(57167) <= 15736501;
srom_1(57168) <= 15996235;
srom_1(57169) <= 16220294;
srom_1(57170) <= 16407628;
srom_1(57171) <= 16557358;
srom_1(57172) <= 16668781;
srom_1(57173) <= 16741376;
srom_1(57174) <= 16774803;
srom_1(57175) <= 16768903;
srom_1(57176) <= 16723705;
srom_1(57177) <= 16639421;
srom_1(57178) <= 16516447;
srom_1(57179) <= 16355358;
srom_1(57180) <= 16156910;
srom_1(57181) <= 15922034;
srom_1(57182) <= 15651831;
srom_1(57183) <= 15347568;
srom_1(57184) <= 15010672;
srom_1(57185) <= 14642724;
srom_1(57186) <= 14245447;
srom_1(57187) <= 13820706;
srom_1(57188) <= 13370492;
srom_1(57189) <= 12896916;
srom_1(57190) <= 12402199;
srom_1(57191) <= 11888661;
srom_1(57192) <= 11358710;
srom_1(57193) <= 10814831;
srom_1(57194) <= 10259574;
srom_1(57195) <= 9695545;
srom_1(57196) <= 9125386;
srom_1(57197) <= 8551772;
srom_1(57198) <= 7977394;
srom_1(57199) <= 7404943;
srom_1(57200) <= 6837106;
srom_1(57201) <= 6276543;
srom_1(57202) <= 5725886;
srom_1(57203) <= 5187714;
srom_1(57204) <= 4664552;
srom_1(57205) <= 4158854;
srom_1(57206) <= 3672991;
srom_1(57207) <= 3209241;
srom_1(57208) <= 2769778;
srom_1(57209) <= 2356665;
srom_1(57210) <= 1971837;
srom_1(57211) <= 1617099;
srom_1(57212) <= 1294116;
srom_1(57213) <= 1004401;
srom_1(57214) <= 749313;
srom_1(57215) <= 530048;
srom_1(57216) <= 347635;
srom_1(57217) <= 202929;
srom_1(57218) <= 96608;
srom_1(57219) <= 29171;
srom_1(57220) <= 934;
srom_1(57221) <= 12030;
srom_1(57222) <= 62407;
srom_1(57223) <= 151828;
srom_1(57224) <= 279874;
srom_1(57225) <= 445945;
srom_1(57226) <= 649262;
srom_1(57227) <= 888871;
srom_1(57228) <= 1163649;
srom_1(57229) <= 1472308;
srom_1(57230) <= 1813399;
srom_1(57231) <= 2185323;
srom_1(57232) <= 2586337;
srom_1(57233) <= 3014560;
srom_1(57234) <= 3467984;
srom_1(57235) <= 3944482;
srom_1(57236) <= 4441820;
srom_1(57237) <= 4957666;
srom_1(57238) <= 5489600;
srom_1(57239) <= 6035130;
srom_1(57240) <= 6591695;
srom_1(57241) <= 7156687;
srom_1(57242) <= 7727456;
srom_1(57243) <= 8301325;
srom_1(57244) <= 8875603;
srom_1(57245) <= 9447598;
srom_1(57246) <= 10014626;
srom_1(57247) <= 10574030;
srom_1(57248) <= 11123185;
srom_1(57249) <= 11659518;
srom_1(57250) <= 12180511;
srom_1(57251) <= 12683723;
srom_1(57252) <= 13166794;
srom_1(57253) <= 13627459;
srom_1(57254) <= 14063556;
srom_1(57255) <= 14473042;
srom_1(57256) <= 14853996;
srom_1(57257) <= 15204631;
srom_1(57258) <= 15523304;
srom_1(57259) <= 15808519;
srom_1(57260) <= 16058940;
srom_1(57261) <= 16273392;
srom_1(57262) <= 16450870;
srom_1(57263) <= 16590541;
srom_1(57264) <= 16691751;
srom_1(57265) <= 16754024;
srom_1(57266) <= 16777068;
srom_1(57267) <= 16760777;
srom_1(57268) <= 16705225;
srom_1(57269) <= 16610674;
srom_1(57270) <= 16477567;
srom_1(57271) <= 16306528;
srom_1(57272) <= 16098359;
srom_1(57273) <= 15854036;
srom_1(57274) <= 15574705;
srom_1(57275) <= 15261677;
srom_1(57276) <= 14916418;
srom_1(57277) <= 14540548;
srom_1(57278) <= 14135829;
srom_1(57279) <= 13704160;
srom_1(57280) <= 13247564;
srom_1(57281) <= 12768183;
srom_1(57282) <= 12268265;
srom_1(57283) <= 11750153;
srom_1(57284) <= 11216278;
srom_1(57285) <= 10669143;
srom_1(57286) <= 10111314;
srom_1(57287) <= 9545407;
srom_1(57288) <= 8974075;
srom_1(57289) <= 8399997;
srom_1(57290) <= 7825866;
srom_1(57291) <= 7254374;
srom_1(57292) <= 6688201;
srom_1(57293) <= 6130002;
srom_1(57294) <= 5582393;
srom_1(57295) <= 5047945;
srom_1(57296) <= 4529161;
srom_1(57297) <= 4028476;
srom_1(57298) <= 3548237;
srom_1(57299) <= 3090697;
srom_1(57300) <= 2658000;
srom_1(57301) <= 2252175;
srom_1(57302) <= 1875127;
srom_1(57303) <= 1528623;
srom_1(57304) <= 1214287;
srom_1(57305) <= 933594;
srom_1(57306) <= 687861;
srom_1(57307) <= 478238;
srom_1(57308) <= 305711;
srom_1(57309) <= 171086;
srom_1(57310) <= 74997;
srom_1(57311) <= 17893;
srom_1(57312) <= 42;
srom_1(57313) <= 21527;
srom_1(57314) <= 82249;
srom_1(57315) <= 181923;
srom_1(57316) <= 320080;
srom_1(57317) <= 496073;
srom_1(57318) <= 709078;
srom_1(57319) <= 958094;
srom_1(57320) <= 1241954;
srom_1(57321) <= 1559327;
srom_1(57322) <= 1908726;
srom_1(57323) <= 2288510;
srom_1(57324) <= 2696901;
srom_1(57325) <= 3131981;
srom_1(57326) <= 3591712;
srom_1(57327) <= 4073937;
srom_1(57328) <= 4576394;
srom_1(57329) <= 5096729;
srom_1(57330) <= 5632501;
srom_1(57331) <= 6181196;
srom_1(57332) <= 6740243;
srom_1(57333) <= 7307020;
srom_1(57334) <= 7878869;
srom_1(57335) <= 8453108;
srom_1(57336) <= 9027044;
srom_1(57337) <= 9597987;
srom_1(57338) <= 10163259;
srom_1(57339) <= 10720208;
srom_1(57340) <= 11266224;
srom_1(57341) <= 11798746;
srom_1(57342) <= 12315276;
srom_1(57343) <= 12813393;
srom_1(57344) <= 13290761;
srom_1(57345) <= 13745140;
srom_1(57346) <= 14174401;
srom_1(57347) <= 14576531;
srom_1(57348) <= 14949643;
srom_1(57349) <= 15291988;
srom_1(57350) <= 15601961;
srom_1(57351) <= 15878108;
srom_1(57352) <= 16119134;
srom_1(57353) <= 16323909;
srom_1(57354) <= 16491473;
srom_1(57355) <= 16621040;
srom_1(57356) <= 16712002;
srom_1(57357) <= 16763932;
srom_1(57358) <= 16776588;
srom_1(57359) <= 16749910;
srom_1(57360) <= 16684022;
srom_1(57361) <= 16579235;
srom_1(57362) <= 16436039;
srom_1(57363) <= 16255106;
srom_1(57364) <= 16037284;
srom_1(57365) <= 15783594;
srom_1(57366) <= 15495228;
srom_1(57367) <= 15173535;
srom_1(57368) <= 14820026;
srom_1(57369) <= 14436358;
srom_1(57370) <= 14024330;
srom_1(57371) <= 13585874;
srom_1(57372) <= 13123046;
srom_1(57373) <= 12638017;
srom_1(57374) <= 12133060;
srom_1(57375) <= 11610545;
srom_1(57376) <= 11072921;
srom_1(57377) <= 10522709;
srom_1(57378) <= 9962490;
srom_1(57379) <= 9394890;
srom_1(57380) <= 8822572;
srom_1(57381) <= 8248218;
srom_1(57382) <= 7674523;
srom_1(57383) <= 7104177;
srom_1(57384) <= 6539853;
srom_1(57385) <= 5984199;
srom_1(57386) <= 5439820;
srom_1(57387) <= 4909269;
srom_1(57388) <= 4395034;
srom_1(57389) <= 3899526;
srom_1(57390) <= 3425069;
srom_1(57391) <= 2973887;
srom_1(57392) <= 2548097;
srom_1(57393) <= 2149695;
srom_1(57394) <= 1780550;
srom_1(57395) <= 1442392;
srom_1(57396) <= 1136807;
srom_1(57397) <= 865228;
srom_1(57398) <= 628929;
srom_1(57399) <= 429018;
srom_1(57400) <= 266433;
srom_1(57401) <= 141934;
srom_1(57402) <= 56108;
srom_1(57403) <= 9355;
srom_1(57404) <= 1895;
srom_1(57405) <= 33764;
srom_1(57406) <= 104811;
srom_1(57407) <= 214704;
srom_1(57408) <= 362927;
srom_1(57409) <= 548785;
srom_1(57410) <= 771407;
srom_1(57411) <= 1029749;
srom_1(57412) <= 1322599;
srom_1(57413) <= 1648583;
srom_1(57414) <= 2006174;
srom_1(57415) <= 2393695;
srom_1(57416) <= 2809327;
srom_1(57417) <= 3251123;
srom_1(57418) <= 3717010;
srom_1(57419) <= 4204804;
srom_1(57420) <= 4712217;
srom_1(57421) <= 5236870;
srom_1(57422) <= 5776303;
srom_1(57423) <= 6327986;
srom_1(57424) <= 6889331;
srom_1(57425) <= 7457707;
srom_1(57426) <= 8030449;
srom_1(57427) <= 8604870;
srom_1(57428) <= 9178277;
srom_1(57429) <= 9747981;
srom_1(57430) <= 10311310;
srom_1(57431) <= 10865623;
srom_1(57432) <= 11408320;
srom_1(57433) <= 11936857;
srom_1(57434) <= 12448755;
srom_1(57435) <= 12941614;
srom_1(57436) <= 13413122;
srom_1(57437) <= 13861068;
srom_1(57438) <= 14283352;
srom_1(57439) <= 14677994;
srom_1(57440) <= 15043142;
srom_1(57441) <= 15377086;
srom_1(57442) <= 15678257;
srom_1(57443) <= 15945245;
srom_1(57444) <= 16176798;
srom_1(57445) <= 16371828;
srom_1(57446) <= 16529423;
srom_1(57447) <= 16648843;
srom_1(57448) <= 16729527;
srom_1(57449) <= 16771099;
srom_1(57450) <= 16773361;
srom_1(57451) <= 16736305;
srom_1(57452) <= 16660104;
srom_1(57453) <= 16545114;
srom_1(57454) <= 16391876;
srom_1(57455) <= 16201108;
srom_1(57456) <= 15973704;
srom_1(57457) <= 15710732;
srom_1(57458) <= 15413423;
srom_1(57459) <= 15083173;
srom_1(57460) <= 14721529;
srom_1(57461) <= 14330188;
srom_1(57462) <= 13910985;
srom_1(57463) <= 13465886;
srom_1(57464) <= 12996977;
srom_1(57465) <= 12506459;
srom_1(57466) <= 11996630;
srom_1(57467) <= 11469882;
srom_1(57468) <= 10928685;
srom_1(57469) <= 10375577;
srom_1(57470) <= 9813151;
srom_1(57471) <= 9244045;
srom_1(57472) <= 8670927;
srom_1(57473) <= 8096486;
srom_1(57474) <= 7523414;
srom_1(57475) <= 6954399;
srom_1(57476) <= 6392110;
srom_1(57477) <= 5839184;
srom_1(57478) <= 5298212;
srom_1(57479) <= 4771733;
srom_1(57480) <= 4262214;
srom_1(57481) <= 3772045;
srom_1(57482) <= 3303525;
srom_1(57483) <= 2858850;
srom_1(57484) <= 2440107;
srom_1(57485) <= 2049258;
srom_1(57486) <= 1688136;
srom_1(57487) <= 1358435;
srom_1(57488) <= 1061701;
srom_1(57489) <= 799326;
srom_1(57490) <= 572539;
srom_1(57491) <= 382404;
srom_1(57492) <= 229814;
srom_1(57493) <= 115482;
srom_1(57494) <= 39946;
srom_1(57495) <= 3560;
srom_1(57496) <= 6495;
srom_1(57497) <= 48735;
srom_1(57498) <= 130085;
srom_1(57499) <= 250161;
srom_1(57500) <= 408402;
srom_1(57501) <= 604064;
srom_1(57502) <= 836231;
srom_1(57503) <= 1103813;
srom_1(57504) <= 1405556;
srom_1(57505) <= 1740046;
srom_1(57506) <= 2105712;
srom_1(57507) <= 2500842;
srom_1(57508) <= 2923581;
srom_1(57509) <= 3371947;
srom_1(57510) <= 3843838;
srom_1(57511) <= 4337041;
srom_1(57512) <= 4849244;
srom_1(57513) <= 5378043;
srom_1(57514) <= 5920961;
srom_1(57515) <= 6475450;
srom_1(57516) <= 7038910;
srom_1(57517) <= 7608699;
srom_1(57518) <= 8182146;
srom_1(57519) <= 8756561;
srom_1(57520) <= 9329251;
srom_1(57521) <= 9897529;
srom_1(57522) <= 10458732;
srom_1(57523) <= 11010227;
srom_1(57524) <= 11549428;
srom_1(57525) <= 12073807;
srom_1(57526) <= 12580906;
srom_1(57527) <= 13068344;
srom_1(57528) <= 13533838;
srom_1(57529) <= 13975205;
srom_1(57530) <= 14390374;
srom_1(57531) <= 14777398;
srom_1(57532) <= 15134463;
srom_1(57533) <= 15459895;
srom_1(57534) <= 15752167;
srom_1(57535) <= 16009908;
srom_1(57536) <= 16231911;
srom_1(57537) <= 16417134;
srom_1(57538) <= 16564708;
srom_1(57539) <= 16673942;
srom_1(57540) <= 16744322;
srom_1(57541) <= 16775521;
srom_1(57542) <= 16767389;
srom_1(57543) <= 16719967;
srom_1(57544) <= 16633477;
srom_1(57545) <= 16508323;
srom_1(57546) <= 16345093;
srom_1(57547) <= 16144553;
srom_1(57548) <= 15907642;
srom_1(57549) <= 15635472;
srom_1(57550) <= 15329319;
srom_1(57551) <= 14990618;
srom_1(57552) <= 14620958;
srom_1(57553) <= 14222073;
srom_1(57554) <= 13795833;
srom_1(57555) <= 13344236;
srom_1(57556) <= 12869400;
srom_1(57557) <= 12373553;
srom_1(57558) <= 11859019;
srom_1(57559) <= 11328210;
srom_1(57560) <= 10783618;
srom_1(57561) <= 10227794;
srom_1(57562) <= 9663345;
srom_1(57563) <= 9092919;
srom_1(57564) <= 8519190;
srom_1(57565) <= 7944848;
srom_1(57566) <= 7372588;
srom_1(57567) <= 6805092;
srom_1(57568) <= 6245021;
srom_1(57569) <= 5695003;
srom_1(57570) <= 5157616;
srom_1(57571) <= 4635380;
srom_1(57572) <= 4130744;
srom_1(57573) <= 3646075;
srom_1(57574) <= 3183646;
srom_1(57575) <= 2745624;
srom_1(57576) <= 2334064;
srom_1(57577) <= 1950895;
srom_1(57578) <= 1597916;
srom_1(57579) <= 1276780;
srom_1(57580) <= 988994;
srom_1(57581) <= 735908;
srom_1(57582) <= 518707;
srom_1(57583) <= 338411;
srom_1(57584) <= 195866;
srom_1(57585) <= 91739;
srom_1(57586) <= 26519;
srom_1(57587) <= 511;
srom_1(57588) <= 13838;
srom_1(57589) <= 66438;
srom_1(57590) <= 158062;
srom_1(57591) <= 288283;
srom_1(57592) <= 456489;
srom_1(57593) <= 661891;
srom_1(57594) <= 903527;
srom_1(57595) <= 1180262;
srom_1(57596) <= 1490801;
srom_1(57597) <= 1833685;
srom_1(57598) <= 2207307;
srom_1(57599) <= 2609916;
srom_1(57600) <= 3039623;
srom_1(57601) <= 3494413;
srom_1(57602) <= 3972154;
srom_1(57603) <= 4470605;
srom_1(57604) <= 4987429;
srom_1(57605) <= 5520202;
srom_1(57606) <= 6066426;
srom_1(57607) <= 6623540;
srom_1(57608) <= 7188931;
srom_1(57609) <= 7759947;
srom_1(57610) <= 8333911;
srom_1(57611) <= 8908132;
srom_1(57612) <= 9479917;
srom_1(57613) <= 10046584;
srom_1(57614) <= 10605476;
srom_1(57615) <= 11153972;
srom_1(57616) <= 11689501;
srom_1(57617) <= 12209551;
srom_1(57618) <= 12711683;
srom_1(57619) <= 13193543;
srom_1(57620) <= 13652870;
srom_1(57621) <= 14087512;
srom_1(57622) <= 14495430;
srom_1(57623) <= 14874710;
srom_1(57624) <= 15223575;
srom_1(57625) <= 15540389;
srom_1(57626) <= 15823665;
srom_1(57627) <= 16072076;
srom_1(57628) <= 16284456;
srom_1(57629) <= 16459811;
srom_1(57630) <= 16597316;
srom_1(57631) <= 16696328;
srom_1(57632) <= 16756382;
srom_1(57633) <= 16777197;
srom_1(57634) <= 16758675;
srom_1(57635) <= 16700902;
srom_1(57636) <= 16604151;
srom_1(57637) <= 16468874;
srom_1(57638) <= 16295706;
srom_1(57639) <= 16085458;
srom_1(57640) <= 15839118;
srom_1(57641) <= 15557839;
srom_1(57642) <= 15242942;
srom_1(57643) <= 14895902;
srom_1(57644) <= 14518347;
srom_1(57645) <= 14112048;
srom_1(57646) <= 13678910;
srom_1(57647) <= 13220963;
srom_1(57648) <= 12740356;
srom_1(57649) <= 12239342;
srom_1(57650) <= 11720271;
srom_1(57651) <= 11185576;
srom_1(57652) <= 10637766;
srom_1(57653) <= 10079408;
srom_1(57654) <= 9513122;
srom_1(57655) <= 8941562;
srom_1(57656) <= 8367409;
srom_1(57657) <= 7793356;
srom_1(57658) <= 7222094;
srom_1(57659) <= 6656303;
srom_1(57660) <= 6098634;
srom_1(57661) <= 5551704;
srom_1(57662) <= 5018078;
srom_1(57663) <= 4500257;
srom_1(57664) <= 4000669;
srom_1(57665) <= 3521658;
srom_1(57666) <= 3065471;
srom_1(57667) <= 2634245;
srom_1(57668) <= 2230003;
srom_1(57669) <= 1854641;
srom_1(57670) <= 1509919;
srom_1(57671) <= 1197453;
srom_1(57672) <= 918710;
srom_1(57673) <= 674995;
srom_1(57674) <= 467452;
srom_1(57675) <= 297054;
srom_1(57676) <= 164600;
srom_1(57677) <= 70712;
srom_1(57678) <= 15828;
srom_1(57679) <= 208;
srom_1(57680) <= 23924;
srom_1(57681) <= 86864;
srom_1(57682) <= 188735;
srom_1(57683) <= 329057;
srom_1(57684) <= 507173;
srom_1(57685) <= 722248;
srom_1(57686) <= 973273;
srom_1(57687) <= 1259072;
srom_1(57688) <= 1578303;
srom_1(57689) <= 1929470;
srom_1(57690) <= 2310926;
srom_1(57691) <= 2720882;
srom_1(57692) <= 3157417;
srom_1(57693) <= 3618482;
srom_1(57694) <= 4101916;
srom_1(57695) <= 4605452;
srom_1(57696) <= 5126728;
srom_1(57697) <= 5663300;
srom_1(57698) <= 6212652;
srom_1(57699) <= 6772208;
srom_1(57700) <= 7339344;
srom_1(57701) <= 7911400;
srom_1(57702) <= 8485694;
srom_1(57703) <= 9059533;
srom_1(57704) <= 9630225;
srom_1(57705) <= 10195095;
srom_1(57706) <= 10751494;
srom_1(57707) <= 11296813;
srom_1(57708) <= 11828494;
srom_1(57709) <= 12344044;
srom_1(57710) <= 12841045;
srom_1(57711) <= 13317168;
srom_1(57712) <= 13770179;
srom_1(57713) <= 14197954;
srom_1(57714) <= 14598487;
srom_1(57715) <= 14969899;
srom_1(57716) <= 15310450;
srom_1(57717) <= 15618542;
srom_1(57718) <= 15892730;
srom_1(57719) <= 16131728;
srom_1(57720) <= 16334417;
srom_1(57721) <= 16499845;
srom_1(57722) <= 16627236;
srom_1(57723) <= 16715994;
srom_1(57724) <= 16765702;
srom_1(57725) <= 16776127;
srom_1(57726) <= 16747219;
srom_1(57727) <= 16679116;
srom_1(57728) <= 16572135;
srom_1(57729) <= 16426779;
srom_1(57730) <= 16243729;
srom_1(57731) <= 16023844;
srom_1(57732) <= 15768154;
srom_1(57733) <= 15477860;
srom_1(57734) <= 15154321;
srom_1(57735) <= 14799056;
srom_1(57736) <= 14413729;
srom_1(57737) <= 14000149;
srom_1(57738) <= 13560255;
srom_1(57739) <= 13096109;
srom_1(57740) <= 12609887;
srom_1(57741) <= 12103871;
srom_1(57742) <= 11580433;
srom_1(57743) <= 11042027;
srom_1(57744) <= 10491178;
srom_1(57745) <= 9930469;
srom_1(57746) <= 9362530;
srom_1(57747) <= 8790025;
srom_1(57748) <= 8215636;
srom_1(57749) <= 7642059;
srom_1(57750) <= 7071983;
srom_1(57751) <= 6508081;
srom_1(57752) <= 5952997;
srom_1(57753) <= 5409334;
srom_1(57754) <= 4879643;
srom_1(57755) <= 4366406;
srom_1(57756) <= 3872031;
srom_1(57757) <= 3398835;
srom_1(57758) <= 2949038;
srom_1(57759) <= 2524749;
srom_1(57760) <= 2127958;
srom_1(57761) <= 1760525;
srom_1(57762) <= 1424174;
srom_1(57763) <= 1120481;
srom_1(57764) <= 850871;
srom_1(57765) <= 616608;
srom_1(57766) <= 418790;
srom_1(57767) <= 258346;
srom_1(57768) <= 136027;
srom_1(57769) <= 52408;
srom_1(57770) <= 7879;
srom_1(57771) <= 2651;
srom_1(57772) <= 36748;
srom_1(57773) <= 110009;
srom_1(57774) <= 222091;
srom_1(57775) <= 372469;
srom_1(57776) <= 560438;
srom_1(57777) <= 785115;
srom_1(57778) <= 1045448;
srom_1(57779) <= 1340215;
srom_1(57780) <= 1668035;
srom_1(57781) <= 2027370;
srom_1(57782) <= 2416534;
srom_1(57783) <= 2833704;
srom_1(57784) <= 3276923;
srom_1(57785) <= 3744112;
srom_1(57786) <= 4233081;
srom_1(57787) <= 4741537;
srom_1(57788) <= 5267094;
srom_1(57789) <= 5807290;
srom_1(57790) <= 6359590;
srom_1(57791) <= 6921406;
srom_1(57792) <= 7490101;
srom_1(57793) <= 8063010;
srom_1(57794) <= 8637445;
srom_1(57795) <= 9210714;
srom_1(57796) <= 9780127;
srom_1(57797) <= 10343016;
srom_1(57798) <= 10896739;
srom_1(57799) <= 11438701;
srom_1(57800) <= 11966360;
srom_1(57801) <= 12477241;
srom_1(57802) <= 12968950;
srom_1(57803) <= 13439180;
srom_1(57804) <= 13885725;
srom_1(57805) <= 14306493;
srom_1(57806) <= 14699510;
srom_1(57807) <= 15062933;
srom_1(57808) <= 15395058;
srom_1(57809) <= 15694327;
srom_1(57810) <= 15959337;
srom_1(57811) <= 16188846;
srom_1(57812) <= 16381776;
srom_1(57813) <= 16537224;
srom_1(57814) <= 16654460;
srom_1(57815) <= 16732934;
srom_1(57816) <= 16772279;
srom_1(57817) <= 16772311;
srom_1(57818) <= 16733028;
srom_1(57819) <= 16654615;
srom_1(57820) <= 16537440;
srom_1(57821) <= 16382052;
srom_1(57822) <= 16189181;
srom_1(57823) <= 15959730;
srom_1(57824) <= 15694775;
srom_1(57825) <= 15395559;
srom_1(57826) <= 15063485;
srom_1(57827) <= 14700110;
srom_1(57828) <= 14307139;
srom_1(57829) <= 13886413;
srom_1(57830) <= 13439907;
srom_1(57831) <= 12969713;
srom_1(57832) <= 12478036;
srom_1(57833) <= 11967183;
srom_1(57834) <= 11439549;
srom_1(57835) <= 10897608;
srom_1(57836) <= 10343901;
srom_1(57837) <= 9781026;
srom_1(57838) <= 9211620;
srom_1(57839) <= 8638356;
srom_1(57840) <= 8063920;
srom_1(57841) <= 7491006;
srom_1(57842) <= 6922302;
srom_1(57843) <= 6360474;
srom_1(57844) <= 5808157;
srom_1(57845) <= 5267940;
srom_1(57846) <= 4742357;
srom_1(57847) <= 4233872;
srom_1(57848) <= 3744871;
srom_1(57849) <= 3277645;
srom_1(57850) <= 2834387;
srom_1(57851) <= 2417174;
srom_1(57852) <= 2027963;
srom_1(57853) <= 1668580;
srom_1(57854) <= 1340709;
srom_1(57855) <= 1045888;
srom_1(57856) <= 785500;
srom_1(57857) <= 560765;
srom_1(57858) <= 372738;
srom_1(57859) <= 222300;
srom_1(57860) <= 110156;
srom_1(57861) <= 36833;
srom_1(57862) <= 2674;
srom_1(57863) <= 7840;
srom_1(57864) <= 52306;
srom_1(57865) <= 135864;
srom_1(57866) <= 258122;
srom_1(57867) <= 418506;
srom_1(57868) <= 616265;
srom_1(57869) <= 850471;
srom_1(57870) <= 1120026;
srom_1(57871) <= 1423666;
srom_1(57872) <= 1759967;
srom_1(57873) <= 2127352;
srom_1(57874) <= 2524098;
srom_1(57875) <= 2948345;
srom_1(57876) <= 3398103;
srom_1(57877) <= 3871263;
srom_1(57878) <= 4365607;
srom_1(57879) <= 4878816;
srom_1(57880) <= 5408483;
srom_1(57881) <= 5952125;
srom_1(57882) <= 6507193;
srom_1(57883) <= 7071083;
srom_1(57884) <= 7641152;
srom_1(57885) <= 8214726;
srom_1(57886) <= 8789115;
srom_1(57887) <= 9361626;
srom_1(57888) <= 9929574;
srom_1(57889) <= 10490296;
srom_1(57890) <= 11041163;
srom_1(57891) <= 11579590;
srom_1(57892) <= 12103054;
srom_1(57893) <= 12609100;
srom_1(57894) <= 13095355;
srom_1(57895) <= 13559538;
srom_1(57896) <= 13999472;
srom_1(57897) <= 14413096;
srom_1(57898) <= 14798468;
srom_1(57899) <= 15153782;
srom_1(57900) <= 15477373;
srom_1(57901) <= 15767721;
srom_1(57902) <= 16023467;
srom_1(57903) <= 16243409;
srom_1(57904) <= 16426518;
srom_1(57905) <= 16571935;
srom_1(57906) <= 16678977;
srom_1(57907) <= 16747142;
srom_1(57908) <= 16776112;
srom_1(57909) <= 16765750;
srom_1(57910) <= 16716104;
srom_1(57911) <= 16627408;
srom_1(57912) <= 16500077;
srom_1(57913) <= 16334709;
srom_1(57914) <= 16132079;
srom_1(57915) <= 15893137;
srom_1(57916) <= 15619003;
srom_1(57917) <= 15310964;
srom_1(57918) <= 14970464;
srom_1(57919) <= 14599099;
srom_1(57920) <= 14198611;
srom_1(57921) <= 13770878;
srom_1(57922) <= 13317905;
srom_1(57923) <= 12841817;
srom_1(57924) <= 12344847;
srom_1(57925) <= 11829324;
srom_1(57926) <= 11297667;
srom_1(57927) <= 10752368;
srom_1(57928) <= 10195985;
srom_1(57929) <= 9631126;
srom_1(57930) <= 9060441;
srom_1(57931) <= 8486605;
srom_1(57932) <= 7912309;
srom_1(57933) <= 7340248;
srom_1(57934) <= 6773102;
srom_1(57935) <= 6213532;
srom_1(57936) <= 5664161;
srom_1(57937) <= 5127567;
srom_1(57938) <= 4606264;
srom_1(57939) <= 4102699;
srom_1(57940) <= 3619231;
srom_1(57941) <= 3158129;
srom_1(57942) <= 2721554;
srom_1(57943) <= 2311554;
srom_1(57944) <= 1930051;
srom_1(57945) <= 1578835;
srom_1(57946) <= 1259552;
srom_1(57947) <= 973699;
srom_1(57948) <= 722618;
srom_1(57949) <= 507485;
srom_1(57950) <= 329310;
srom_1(57951) <= 188927;
srom_1(57952) <= 86995;
srom_1(57953) <= 23992;
srom_1(57954) <= 214;
srom_1(57955) <= 15772;
srom_1(57956) <= 70594;
srom_1(57957) <= 164421;
srom_1(57958) <= 296814;
srom_1(57959) <= 467152;
srom_1(57960) <= 674637;
srom_1(57961) <= 918295;
srom_1(57962) <= 1196984;
srom_1(57963) <= 1509398;
srom_1(57964) <= 1854070;
srom_1(57965) <= 2229384;
srom_1(57966) <= 2633582;
srom_1(57967) <= 3064767;
srom_1(57968) <= 3520917;
srom_1(57969) <= 3999893;
srom_1(57970) <= 4499450;
srom_1(57971) <= 5017244;
srom_1(57972) <= 5550847;
srom_1(57973) <= 6097758;
srom_1(57974) <= 6655411;
srom_1(57975) <= 7221192;
srom_1(57976) <= 7792448;
srom_1(57977) <= 8366499;
srom_1(57978) <= 8940653;
srom_1(57979) <= 9512219;
srom_1(57980) <= 10078516;
srom_1(57981) <= 10636888;
srom_1(57982) <= 11184718;
srom_1(57983) <= 11719435;
srom_1(57984) <= 12238533;
srom_1(57985) <= 12739577;
srom_1(57986) <= 13220219;
srom_1(57987) <= 13678203;
srom_1(57988) <= 14111382;
srom_1(57989) <= 14517725;
srom_1(57990) <= 14895327;
srom_1(57991) <= 15242417;
srom_1(57992) <= 15557366;
srom_1(57993) <= 15838699;
srom_1(57994) <= 16085096;
srom_1(57995) <= 16295401;
srom_1(57996) <= 16468629;
srom_1(57997) <= 16603967;
srom_1(57998) <= 16700780;
srom_1(57999) <= 16758614;
srom_1(58000) <= 16777199;
srom_1(58001) <= 16756446;
srom_1(58002) <= 16696454;
srom_1(58003) <= 16597503;
srom_1(58004) <= 16460059;
srom_1(58005) <= 16284764;
srom_1(58006) <= 16072442;
srom_1(58007) <= 15824087;
srom_1(58008) <= 15540865;
srom_1(58009) <= 15224103;
srom_1(58010) <= 14875288;
srom_1(58011) <= 14496054;
srom_1(58012) <= 14088180;
srom_1(58013) <= 13653580;
srom_1(58014) <= 13194289;
srom_1(58015) <= 12712464;
srom_1(58016) <= 12210362;
srom_1(58017) <= 11690339;
srom_1(58018) <= 11154832;
srom_1(58019) <= 10606354;
srom_1(58020) <= 10047476;
srom_1(58021) <= 9480820;
srom_1(58022) <= 8909041;
srom_1(58023) <= 8334822;
srom_1(58024) <= 7760855;
srom_1(58025) <= 7189832;
srom_1(58026) <= 6624430;
srom_1(58027) <= 6067302;
srom_1(58028) <= 5521058;
srom_1(58029) <= 4988262;
srom_1(58030) <= 4471410;
srom_1(58031) <= 3972928;
srom_1(58032) <= 3495153;
srom_1(58033) <= 3040325;
srom_1(58034) <= 2610576;
srom_1(58035) <= 2207923;
srom_1(58036) <= 1834253;
srom_1(58037) <= 1491319;
srom_1(58038) <= 1180728;
srom_1(58039) <= 903938;
srom_1(58040) <= 662246;
srom_1(58041) <= 456785;
srom_1(58042) <= 288520;
srom_1(58043) <= 158238;
srom_1(58044) <= 66552;
srom_1(58045) <= 13891;
srom_1(58046) <= 501;
srom_1(58047) <= 26446;
srom_1(58048) <= 91604;
srom_1(58049) <= 195670;
srom_1(58050) <= 338155;
srom_1(58051) <= 518392;
srom_1(58052) <= 735535;
srom_1(58053) <= 988565;
srom_1(58054) <= 1276297;
srom_1(58055) <= 1597381;
srom_1(58056) <= 1950311;
srom_1(58057) <= 2333433;
srom_1(58058) <= 2744950;
srom_1(58059) <= 3182931;
srom_1(58060) <= 3645324;
srom_1(58061) <= 4129960;
srom_1(58062) <= 4634566;
srom_1(58063) <= 5156775;
srom_1(58064) <= 5694141;
srom_1(58065) <= 6244141;
srom_1(58066) <= 6804197;
srom_1(58067) <= 7371684;
srom_1(58068) <= 7943939;
srom_1(58069) <= 8518279;
srom_1(58070) <= 9092011;
srom_1(58071) <= 9662445;
srom_1(58072) <= 10226905;
srom_1(58073) <= 10782745;
srom_1(58074) <= 11327357;
srom_1(58075) <= 11858189;
srom_1(58076) <= 12372751;
srom_1(58077) <= 12868630;
srom_1(58078) <= 13343501;
srom_1(58079) <= 13795136;
srom_1(58080) <= 14221418;
srom_1(58081) <= 14620349;
srom_1(58082) <= 14990056;
srom_1(58083) <= 15328807;
srom_1(58084) <= 15635013;
srom_1(58085) <= 15907238;
srom_1(58086) <= 16144206;
srom_1(58087) <= 16344805;
srom_1(58088) <= 16508094;
srom_1(58089) <= 16633309;
srom_1(58090) <= 16719861;
srom_1(58091) <= 16767345;
srom_1(58092) <= 16775539;
srom_1(58093) <= 16744403;
srom_1(58094) <= 16674084;
srom_1(58095) <= 16564912;
srom_1(58096) <= 16417398;
srom_1(58097) <= 16232234;
srom_1(58098) <= 16010289;
srom_1(58099) <= 15752603;
srom_1(58100) <= 15460385;
srom_1(58101) <= 15135005;
srom_1(58102) <= 14777988;
srom_1(58103) <= 14391010;
srom_1(58104) <= 13975884;
srom_1(58105) <= 13534558;
srom_1(58106) <= 13069100;
srom_1(58107) <= 12581694;
srom_1(58108) <= 12074626;
srom_1(58109) <= 11550272;
srom_1(58110) <= 11011092;
srom_1(58111) <= 10459614;
srom_1(58112) <= 9898425;
srom_1(58113) <= 9330156;
srom_1(58114) <= 8757471;
srom_1(58115) <= 8183057;
srom_1(58116) <= 7609606;
srom_1(58117) <= 7039809;
srom_1(58118) <= 6476336;
srom_1(58119) <= 5921831;
srom_1(58120) <= 5378894;
srom_1(58121) <= 4850070;
srom_1(58122) <= 4337839;
srom_1(58123) <= 3844604;
srom_1(58124) <= 3372677;
srom_1(58125) <= 2924272;
srom_1(58126) <= 2501490;
srom_1(58127) <= 2106316;
srom_1(58128) <= 1740601;
srom_1(58129) <= 1406061;
srom_1(58130) <= 1104265;
srom_1(58131) <= 836627;
srom_1(58132) <= 604403;
srom_1(58133) <= 408682;
srom_1(58134) <= 250382;
srom_1(58135) <= 130245;
srom_1(58136) <= 48834;
srom_1(58137) <= 6530;
srom_1(58138) <= 3534;
srom_1(58139) <= 39858;
srom_1(58140) <= 115332;
srom_1(58141) <= 229602;
srom_1(58142) <= 382133;
srom_1(58143) <= 572208;
srom_1(58144) <= 798938;
srom_1(58145) <= 1061258;
srom_1(58146) <= 1357938;
srom_1(58147) <= 1687588;
srom_1(58148) <= 2048661;
srom_1(58149) <= 2439464;
srom_1(58150) <= 2858165;
srom_1(58151) <= 3302800;
srom_1(58152) <= 3771284;
srom_1(58153) <= 4261421;
srom_1(58154) <= 4770911;
srom_1(58155) <= 5297365;
srom_1(58156) <= 5838316;
srom_1(58157) <= 6391226;
srom_1(58158) <= 6953502;
srom_1(58159) <= 7522508;
srom_1(58160) <= 8095575;
srom_1(58161) <= 8670017;
srom_1(58162) <= 9243139;
srom_1(58163) <= 9812253;
srom_1(58164) <= 10374692;
srom_1(58165) <= 10927817;
srom_1(58166) <= 11469035;
srom_1(58167) <= 11995808;
srom_1(58168) <= 12505665;
srom_1(58169) <= 12996216;
srom_1(58170) <= 13465161;
srom_1(58171) <= 13910299;
srom_1(58172) <= 14329545;
srom_1(58173) <= 14720932;
srom_1(58174) <= 15082624;
srom_1(58175) <= 15412925;
srom_1(58176) <= 15710287;
srom_1(58177) <= 15973315;
srom_1(58178) <= 16200776;
srom_1(58179) <= 16391603;
srom_1(58180) <= 16544901;
srom_1(58181) <= 16659952;
srom_1(58182) <= 16736215;
srom_1(58183) <= 16773334;
srom_1(58184) <= 16771133;
srom_1(58185) <= 16729624;
srom_1(58186) <= 16649001;
srom_1(58187) <= 16529643;
srom_1(58188) <= 16372108;
srom_1(58189) <= 16177136;
srom_1(58190) <= 15945641;
srom_1(58191) <= 15678708;
srom_1(58192) <= 15377589;
srom_1(58193) <= 15043697;
srom_1(58194) <= 14678597;
srom_1(58195) <= 14284000;
srom_1(58196) <= 13861759;
srom_1(58197) <= 13413851;
srom_1(58198) <= 12942379;
srom_1(58199) <= 12449552;
srom_1(58200) <= 11937683;
srom_1(58201) <= 11409170;
srom_1(58202) <= 10866493;
srom_1(58203) <= 10312196;
srom_1(58204) <= 9748879;
srom_1(58205) <= 9179184;
srom_1(58206) <= 8605780;
srom_1(58207) <= 8031359;
srom_1(58208) <= 7458613;
srom_1(58209) <= 6890227;
srom_1(58210) <= 6328869;
srom_1(58211) <= 5777169;
srom_1(58212) <= 5237714;
srom_1(58213) <= 4713036;
srom_1(58214) <= 4205594;
srom_1(58215) <= 3717767;
srom_1(58216) <= 3251843;
srom_1(58217) <= 2810007;
srom_1(58218) <= 2394332;
srom_1(58219) <= 2006765;
srom_1(58220) <= 1649126;
srom_1(58221) <= 1323089;
srom_1(58222) <= 1030186;
srom_1(58223) <= 771789;
srom_1(58224) <= 549109;
srom_1(58225) <= 363192;
srom_1(58226) <= 214909;
srom_1(58227) <= 104955;
srom_1(58228) <= 33845;
srom_1(58229) <= 1915;
srom_1(58230) <= 9312;
srom_1(58231) <= 56002;
srom_1(58232) <= 141767;
srom_1(58233) <= 266205;
srom_1(58234) <= 428731;
srom_1(58235) <= 628584;
srom_1(58236) <= 864826;
srom_1(58237) <= 1136349;
srom_1(58238) <= 1441881;
srom_1(58239) <= 1779989;
srom_1(58240) <= 2149086;
srom_1(58241) <= 2547443;
srom_1(58242) <= 2973191;
srom_1(58243) <= 3424334;
srom_1(58244) <= 3898756;
srom_1(58245) <= 4394233;
srom_1(58246) <= 4908440;
srom_1(58247) <= 5438967;
srom_1(58248) <= 5983326;
srom_1(58249) <= 6538965;
srom_1(58250) <= 7103277;
srom_1(58251) <= 7673616;
srom_1(58252) <= 8247308;
srom_1(58253) <= 8821662;
srom_1(58254) <= 9393986;
srom_1(58255) <= 9961596;
srom_1(58256) <= 10521829;
srom_1(58257) <= 11072058;
srom_1(58258) <= 11609704;
srom_1(58259) <= 12132245;
srom_1(58260) <= 12637231;
srom_1(58261) <= 13122294;
srom_1(58262) <= 13585159;
srom_1(58263) <= 14023655;
srom_1(58264) <= 14435727;
srom_1(58265) <= 14819441;
srom_1(58266) <= 15173000;
srom_1(58267) <= 15494744;
srom_1(58268) <= 15783164;
srom_1(58269) <= 16036910;
srom_1(58270) <= 16254789;
srom_1(58271) <= 16435782;
srom_1(58272) <= 16579038;
srom_1(58273) <= 16683887;
srom_1(58274) <= 16749836;
srom_1(58275) <= 16776577;
srom_1(58276) <= 16763983;
srom_1(58277) <= 16712115;
srom_1(58278) <= 16621215;
srom_1(58279) <= 16491709;
srom_1(58280) <= 16324205;
srom_1(58281) <= 16119488;
srom_1(58282) <= 15878518;
srom_1(58283) <= 15602426;
srom_1(58284) <= 15292506;
srom_1(58285) <= 14950211;
srom_1(58286) <= 14577146;
srom_1(58287) <= 14175061;
srom_1(58288) <= 13745841;
srom_1(58289) <= 13291500;
srom_1(58290) <= 12814167;
srom_1(58291) <= 12316081;
srom_1(58292) <= 11799578;
srom_1(58293) <= 11267080;
srom_1(58294) <= 10721083;
srom_1(58295) <= 10164149;
srom_1(58296) <= 9598888;
srom_1(58297) <= 9027953;
srom_1(58298) <= 8454019;
srom_1(58299) <= 7879778;
srom_1(58300) <= 7307923;
srom_1(58301) <= 6741136;
srom_1(58302) <= 6182075;
srom_1(58303) <= 5633361;
srom_1(58304) <= 5097567;
srom_1(58305) <= 4577206;
srom_1(58306) <= 4074718;
srom_1(58307) <= 3592459;
srom_1(58308) <= 3132691;
srom_1(58309) <= 2697570;
srom_1(58310) <= 2289136;
srom_1(58311) <= 1909304;
srom_1(58312) <= 1559856;
srom_1(58313) <= 1242431;
srom_1(58314) <= 958516;
srom_1(58315) <= 709444;
srom_1(58316) <= 496382;
srom_1(58317) <= 320329;
srom_1(58318) <= 182111;
srom_1(58319) <= 82377;
srom_1(58320) <= 21593;
srom_1(58321) <= 44;
srom_1(58322) <= 17833;
srom_1(58323) <= 74875;
srom_1(58324) <= 170903;
srom_1(58325) <= 305467;
srom_1(58326) <= 477935;
srom_1(58327) <= 687499;
srom_1(58328) <= 933177;
srom_1(58329) <= 1213815;
srom_1(58330) <= 1528098;
srom_1(58331) <= 1874553;
srom_1(58332) <= 2251554;
srom_1(58333) <= 2657335;
srom_1(58334) <= 3089991;
srom_1(58335) <= 3547494;
srom_1(58336) <= 4027698;
srom_1(58337) <= 4528353;
srom_1(58338) <= 5047109;
srom_1(58339) <= 5581535;
srom_1(58340) <= 6129124;
srom_1(58341) <= 6687309;
srom_1(58342) <= 7253472;
srom_1(58343) <= 7824958;
srom_1(58344) <= 8399086;
srom_1(58345) <= 8973166;
srom_1(58346) <= 9544505;
srom_1(58347) <= 10110423;
srom_1(58348) <= 10668267;
srom_1(58349) <= 11215421;
srom_1(58350) <= 11749319;
srom_1(58351) <= 12267457;
srom_1(58352) <= 12767406;
srom_1(58353) <= 13246822;
srom_1(58354) <= 13703455;
srom_1(58355) <= 14135166;
srom_1(58356) <= 14539929;
srom_1(58357) <= 14915846;
srom_1(58358) <= 15261155;
srom_1(58359) <= 15574236;
srom_1(58360) <= 15853621;
srom_1(58361) <= 16098000;
srom_1(58362) <= 16306227;
srom_1(58363) <= 16477326;
srom_1(58364) <= 16610493;
srom_1(58365) <= 16705106;
srom_1(58366) <= 16760720;
srom_1(58367) <= 16777074;
srom_1(58368) <= 16754091;
srom_1(58369) <= 16691880;
srom_1(58370) <= 16590732;
srom_1(58371) <= 16451122;
srom_1(58372) <= 16273703;
srom_1(58373) <= 16059309;
srom_1(58374) <= 15808944;
srom_1(58375) <= 15523783;
srom_1(58376) <= 15205162;
srom_1(58377) <= 14854576;
srom_1(58378) <= 14473669;
srom_1(58379) <= 14064227;
srom_1(58380) <= 13628170;
srom_1(58381) <= 13167543;
srom_1(58382) <= 12684506;
srom_1(58383) <= 12181324;
srom_1(58384) <= 11660356;
srom_1(58385) <= 11124046;
srom_1(58386) <= 10574909;
srom_1(58387) <= 10015520;
srom_1(58388) <= 9448501;
srom_1(58389) <= 8876512;
srom_1(58390) <= 8302235;
srom_1(58391) <= 7728364;
srom_1(58392) <= 7157588;
srom_1(58393) <= 6592585;
srom_1(58394) <= 6036004;
srom_1(58395) <= 5490455;
srom_1(58396) <= 4958497;
srom_1(58397) <= 4442623;
srom_1(58398) <= 3945254;
srom_1(58399) <= 3468721;
srom_1(58400) <= 3015260;
srom_1(58401) <= 2586995;
srom_1(58402) <= 2185937;
srom_1(58403) <= 1813964;
srom_1(58404) <= 1472823;
srom_1(58405) <= 1164112;
srom_1(58406) <= 889279;
srom_1(58407) <= 649613;
srom_1(58408) <= 446238;
srom_1(58409) <= 280108;
srom_1(58410) <= 152001;
srom_1(58411) <= 62518;
srom_1(58412) <= 12079;
srom_1(58413) <= 921;
srom_1(58414) <= 29095;
srom_1(58415) <= 96470;
srom_1(58416) <= 202729;
srom_1(58417) <= 347375;
srom_1(58418) <= 529730;
srom_1(58419) <= 748937;
srom_1(58420) <= 1003969;
srom_1(58421) <= 1293630;
srom_1(58422) <= 1616562;
srom_1(58423) <= 1971250;
srom_1(58424) <= 2356032;
srom_1(58425) <= 2769102;
srom_1(58426) <= 3208524;
srom_1(58427) <= 3672238;
srom_1(58428) <= 4158068;
srom_1(58429) <= 4663736;
srom_1(58430) <= 5186872;
srom_1(58431) <= 5725022;
srom_1(58432) <= 6275662;
srom_1(58433) <= 6836211;
srom_1(58434) <= 7404039;
srom_1(58435) <= 7976484;
srom_1(58436) <= 8550862;
srom_1(58437) <= 9124479;
srom_1(58438) <= 9694645;
srom_1(58439) <= 10258687;
srom_1(58440) <= 10813959;
srom_1(58441) <= 11357858;
srom_1(58442) <= 11887833;
srom_1(58443) <= 12401399;
srom_1(58444) <= 12896148;
srom_1(58445) <= 13369759;
srom_1(58446) <= 13820012;
srom_1(58447) <= 14244795;
srom_1(58448) <= 14642117;
srom_1(58449) <= 15010113;
srom_1(58450) <= 15347059;
srom_1(58451) <= 15651375;
srom_1(58452) <= 15921633;
srom_1(58453) <= 16156566;
srom_1(58454) <= 16355072;
srom_1(58455) <= 16516221;
srom_1(58456) <= 16639257;
srom_1(58457) <= 16723602;
srom_1(58458) <= 16768862;
srom_1(58459) <= 16774824;
srom_1(58460) <= 16741461;
srom_1(58461) <= 16668927;
srom_1(58462) <= 16557565;
srom_1(58463) <= 16407895;
srom_1(58464) <= 16220620;
srom_1(58465) <= 15996619;
srom_1(58466) <= 15736940;
srom_1(58467) <= 15442803;
srom_1(58468) <= 15115586;
srom_1(58469) <= 14756824;
srom_1(58470) <= 14368200;
srom_1(58471) <= 13951535;
srom_1(58472) <= 13508783;
srom_1(58473) <= 13042021;
srom_1(58474) <= 12553438;
srom_1(58475) <= 12045325;
srom_1(58476) <= 11520064;
srom_1(58477) <= 10980118;
srom_1(58478) <= 10428020;
srom_1(58479) <= 9866358;
srom_1(58480) <= 9297767;
srom_1(58481) <= 8724912;
srom_1(58482) <= 8150480;
srom_1(58483) <= 7577165;
srom_1(58484) <= 7007655;
srom_1(58485) <= 6444621;
srom_1(58486) <= 5890703;
srom_1(58487) <= 5348498;
srom_1(58488) <= 4820550;
srom_1(58489) <= 4309333;
srom_1(58490) <= 3817245;
srom_1(58491) <= 3346595;
srom_1(58492) <= 2899587;
srom_1(58493) <= 2478320;
srom_1(58494) <= 2084768;
srom_1(58495) <= 1720777;
srom_1(58496) <= 1388054;
srom_1(58497) <= 1088158;
srom_1(58498) <= 822497;
srom_1(58499) <= 592317;
srom_1(58500) <= 398695;
srom_1(58501) <= 242541;
srom_1(58502) <= 124587;
srom_1(58503) <= 45385;
srom_1(58504) <= 5308;
srom_1(58505) <= 4543;
srom_1(58506) <= 43094;
srom_1(58507) <= 120779;
srom_1(58508) <= 237236;
srom_1(58509) <= 391917;
srom_1(58510) <= 584097;
srom_1(58511) <= 812875;
srom_1(58512) <= 1077178;
srom_1(58513) <= 1375767;
srom_1(58514) <= 1707242;
srom_1(58515) <= 2070048;
srom_1(58516) <= 2462484;
srom_1(58517) <= 2882710;
srom_1(58518) <= 3328754;
srom_1(58519) <= 3798526;
srom_1(58520) <= 4289823;
srom_1(58521) <= 4800340;
srom_1(58522) <= 5327683;
srom_1(58523) <= 5869381;
srom_1(58524) <= 6422891;
srom_1(58525) <= 6985620;
srom_1(58526) <= 7554928;
srom_1(58527) <= 8128145;
srom_1(58528) <= 8702584;
srom_1(58529) <= 9275550;
srom_1(58530) <= 9844357;
srom_1(58531) <= 10406338;
srom_1(58532) <= 10958857;
srom_1(58533) <= 11499323;
srom_1(58534) <= 12025202;
srom_1(58535) <= 12534027;
srom_1(58536) <= 13023413;
srom_1(58537) <= 13491065;
srom_1(58538) <= 13934790;
srom_1(58539) <= 14352507;
srom_1(58540) <= 14742257;
srom_1(58541) <= 15102213;
srom_1(58542) <= 15430686;
srom_1(58543) <= 15726137;
srom_1(58544) <= 15987179;
srom_1(58545) <= 16212589;
srom_1(58546) <= 16401310;
srom_1(58547) <= 16552456;
srom_1(58548) <= 16665319;
srom_1(58549) <= 16739370;
srom_1(58550) <= 16774261;
srom_1(58551) <= 16769829;
srom_1(58552) <= 16726095;
srom_1(58553) <= 16643263;
srom_1(58554) <= 16521723;
srom_1(58555) <= 16362043;
srom_1(58556) <= 16164973;
srom_1(58557) <= 15931438;
srom_1(58558) <= 15662531;
srom_1(58559) <= 15359514;
srom_1(58560) <= 15023808;
srom_1(58561) <= 14656988;
srom_1(58562) <= 14260773;
srom_1(58563) <= 13837021;
srom_1(58564) <= 13387720;
srom_1(58565) <= 12914977;
srom_1(58566) <= 12421007;
srom_1(58567) <= 11908129;
srom_1(58568) <= 11378746;
srom_1(58569) <= 10835341;
srom_1(58570) <= 10280463;
srom_1(58571) <= 9716713;
srom_1(58572) <= 9146735;
srom_1(58573) <= 8573202;
srom_1(58574) <= 7998803;
srom_1(58575) <= 7426233;
srom_1(58576) <= 6858175;
srom_1(58577) <= 6297294;
srom_1(58578) <= 5746220;
srom_1(58579) <= 5207537;
srom_1(58580) <= 4683771;
srom_1(58581) <= 4177378;
srom_1(58582) <= 3690733;
srom_1(58583) <= 3226118;
srom_1(58584) <= 2785712;
srom_1(58585) <= 2371580;
srom_1(58586) <= 1985664;
srom_1(58587) <= 1629773;
srom_1(58588) <= 1305576;
srom_1(58589) <= 1014595;
srom_1(58590) <= 758193;
srom_1(58591) <= 537572;
srom_1(58592) <= 353768;
srom_1(58593) <= 207641;
srom_1(58594) <= 99878;
srom_1(58595) <= 30984;
srom_1(58596) <= 1282;
srom_1(58597) <= 10910;
srom_1(58598) <= 59825;
srom_1(58599) <= 147796;
srom_1(58600) <= 274411;
srom_1(58601) <= 439076;
srom_1(58602) <= 641019;
srom_1(58603) <= 879293;
srom_1(58604) <= 1152782;
srom_1(58605) <= 1460201;
srom_1(58606) <= 1800110;
srom_1(58607) <= 2170915;
srom_1(58608) <= 2570877;
srom_1(58609) <= 2998120;
srom_1(58610) <= 3450641;
srom_1(58611) <= 3926317;
srom_1(58612) <= 4422919;
srom_1(58613) <= 4938118;
srom_1(58614) <= 5469496;
srom_1(58615) <= 6014564;
srom_1(58616) <= 6570764;
srom_1(58617) <= 7135489;
srom_1(58618) <= 7706090;
srom_1(58619) <= 8279892;
srom_1(58620) <= 8854203;
srom_1(58621) <= 9426331;
srom_1(58622) <= 9993593;
srom_1(58623) <= 10553329;
srom_1(58624) <= 11102913;
srom_1(58625) <= 11639769;
srom_1(58626) <= 12161380;
srom_1(58627) <= 12665298;
srom_1(58628) <= 13149162;
srom_1(58629) <= 13610701;
srom_1(58630) <= 14047753;
srom_1(58631) <= 14458267;
srom_1(58632) <= 14840318;
srom_1(58633) <= 15192114;
srom_1(58634) <= 15512007;
srom_1(58635) <= 15798496;
srom_1(58636) <= 16050237;
srom_1(58637) <= 16266050;
srom_1(58638) <= 16444924;
srom_1(58639) <= 16586018;
srom_1(58640) <= 16688672;
srom_1(58641) <= 16752404;
srom_1(58642) <= 16776915;
srom_1(58643) <= 16762091;
srom_1(58644) <= 16708000;
srom_1(58645) <= 16614897;
srom_1(58646) <= 16483218;
srom_1(58647) <= 16313581;
srom_1(58648) <= 16106780;
srom_1(58649) <= 15863787;
srom_1(58650) <= 15585740;
srom_1(58651) <= 15273943;
srom_1(58652) <= 14929858;
srom_1(58653) <= 14555099;
srom_1(58654) <= 14151424;
srom_1(58655) <= 13720724;
srom_1(58656) <= 13265021;
srom_1(58657) <= 12786450;
srom_1(58658) <= 12287256;
srom_1(58659) <= 11769780;
srom_1(58660) <= 11236449;
srom_1(58661) <= 10689763;
srom_1(58662) <= 10132286;
srom_1(58663) <= 9566632;
srom_1(58664) <= 8995455;
srom_1(58665) <= 8421431;
srom_1(58666) <= 7847254;
srom_1(58667) <= 7275615;
srom_1(58668) <= 6709196;
srom_1(58669) <= 6150651;
srom_1(58670) <= 5602602;
srom_1(58671) <= 5067617;
srom_1(58672) <= 4548205;
srom_1(58673) <= 4046802;
srom_1(58674) <= 3565759;
srom_1(58675) <= 3107332;
srom_1(58676) <= 2673671;
srom_1(58677) <= 2266810;
srom_1(58678) <= 1888655;
srom_1(58679) <= 1540981;
srom_1(58680) <= 1225418;
srom_1(58681) <= 943446;
srom_1(58682) <= 696386;
srom_1(58683) <= 485398;
srom_1(58684) <= 311471;
srom_1(58685) <= 175420;
srom_1(58686) <= 77884;
srom_1(58687) <= 19319;
srom_1(58688) <= 1;
srom_1(58689) <= 20020;
srom_1(58690) <= 79282;
srom_1(58691) <= 177510;
srom_1(58692) <= 314242;
srom_1(58693) <= 488838;
srom_1(58694) <= 700478;
srom_1(58695) <= 948170;
srom_1(58696) <= 1230754;
srom_1(58697) <= 1546903;
srom_1(58698) <= 1895135;
srom_1(58699) <= 2273817;
srom_1(58700) <= 2681174;
srom_1(58701) <= 3115294;
srom_1(58702) <= 3574144;
srom_1(58703) <= 4055569;
srom_1(58704) <= 4557314;
srom_1(58705) <= 5077025;
srom_1(58706) <= 5612265;
srom_1(58707) <= 6160525;
srom_1(58708) <= 6719232;
srom_1(58709) <= 7285768;
srom_1(58710) <= 7857476;
srom_1(58711) <= 8431674;
srom_1(58712) <= 9005670;
srom_1(58713) <= 9576773;
srom_1(58714) <= 10142304;
srom_1(58715) <= 10699611;
srom_1(58716) <= 11246081;
srom_1(58717) <= 11779152;
srom_1(58718) <= 12296323;
srom_1(58719) <= 12795169;
srom_1(58720) <= 13273351;
srom_1(58721) <= 13728628;
srom_1(58722) <= 14158863;
srom_1(58723) <= 14562039;
srom_1(58724) <= 14936266;
srom_1(58725) <= 15279789;
srom_1(58726) <= 15590996;
srom_1(58727) <= 15868429;
srom_1(58728) <= 16110787;
srom_1(58729) <= 16316933;
srom_1(58730) <= 16485900;
srom_1(58731) <= 16616896;
srom_1(58732) <= 16709307;
srom_1(58733) <= 16762699;
srom_1(58734) <= 16776822;
srom_1(58735) <= 16751610;
srom_1(58736) <= 16687181;
srom_1(58737) <= 16583837;
srom_1(58738) <= 16442063;
srom_1(58739) <= 16262524;
srom_1(58740) <= 16046061;
srom_1(58741) <= 15793689;
srom_1(58742) <= 15506593;
srom_1(58743) <= 15186117;
srom_1(58744) <= 14833766;
srom_1(58745) <= 14451192;
srom_1(58746) <= 14040188;
srom_1(58747) <= 13602681;
srom_1(58748) <= 13140724;
srom_1(58749) <= 12656483;
srom_1(58750) <= 12152228;
srom_1(58751) <= 11630325;
srom_1(58752) <= 11093219;
srom_1(58753) <= 10543431;
srom_1(58754) <= 9983538;
srom_1(58755) <= 9416166;
srom_1(58756) <= 8843976;
srom_1(58757) <= 8269650;
srom_1(58758) <= 7695882;
srom_1(58759) <= 7125362;
srom_1(58760) <= 6560766;
srom_1(58761) <= 6004742;
srom_1(58762) <= 5459896;
srom_1(58763) <= 4928784;
srom_1(58764) <= 4413896;
srom_1(58765) <= 3917647;
srom_1(58766) <= 3442364;
srom_1(58767) <= 2990275;
srom_1(58768) <= 2563502;
srom_1(58769) <= 2164044;
srom_1(58770) <= 1793775;
srom_1(58771) <= 1454431;
srom_1(58772) <= 1147605;
srom_1(58773) <= 874734;
srom_1(58774) <= 637098;
srom_1(58775) <= 435811;
srom_1(58776) <= 271818;
srom_1(58777) <= 145887;
srom_1(58778) <= 58610;
srom_1(58779) <= 10394;
srom_1(58780) <= 1467;
srom_1(58781) <= 31870;
srom_1(58782) <= 101460;
srom_1(58783) <= 209912;
srom_1(58784) <= 356717;
srom_1(58785) <= 541186;
srom_1(58786) <= 762454;
srom_1(58787) <= 1019483;
srom_1(58788) <= 1311070;
srom_1(58789) <= 1635845;
srom_1(58790) <= 1992286;
srom_1(58791) <= 2378721;
srom_1(58792) <= 2793340;
srom_1(58793) <= 3234196;
srom_1(58794) <= 3699223;
srom_1(58795) <= 4186240;
srom_1(58796) <= 4692963;
srom_1(58797) <= 5217017;
srom_1(58798) <= 5755943;
srom_1(58799) <= 6307215;
srom_1(58800) <= 6868247;
srom_1(58801) <= 7436409;
srom_1(58802) <= 8009035;
srom_1(58803) <= 8583442;
srom_1(58804) <= 9156935;
srom_1(58805) <= 9726825;
srom_1(58806) <= 10290440;
srom_1(58807) <= 10845137;
srom_1(58808) <= 11388313;
srom_1(58809) <= 11917424;
srom_1(58810) <= 12429986;
srom_1(58811) <= 12923597;
srom_1(58812) <= 13395942;
srom_1(58813) <= 13844806;
srom_1(58814) <= 14268083;
srom_1(58815) <= 14663790;
srom_1(58816) <= 15030071;
srom_1(58817) <= 15365207;
srom_1(58818) <= 15667627;
srom_1(58819) <= 15935914;
srom_1(58820) <= 16168809;
srom_1(58821) <= 16365220;
srom_1(58822) <= 16524225;
srom_1(58823) <= 16645080;
srom_1(58824) <= 16727218;
srom_1(58825) <= 16770253;
srom_1(58826) <= 16773983;
srom_1(58827) <= 16738392;
srom_1(58828) <= 16663646;
srom_1(58829) <= 16550095;
srom_1(58830) <= 16398272;
srom_1(58831) <= 16208889;
srom_1(58832) <= 15982834;
srom_1(58833) <= 15721167;
srom_1(58834) <= 15425115;
srom_1(58835) <= 15096067;
srom_1(58836) <= 14735565;
srom_1(58837) <= 14345299;
srom_1(58838) <= 13927101;
srom_1(58839) <= 13482931;
srom_1(58840) <= 13014872;
srom_1(58841) <= 12525119;
srom_1(58842) <= 12015969;
srom_1(58843) <= 11489808;
srom_1(58844) <= 10949105;
srom_1(58845) <= 10396394;
srom_1(58846) <= 9834269;
srom_1(58847) <= 9265364;
srom_1(58848) <= 8692348;
srom_1(58849) <= 8117908;
srom_1(58850) <= 7544736;
srom_1(58851) <= 6975523;
srom_1(58852) <= 6412935;
srom_1(58853) <= 5859612;
srom_1(58854) <= 5318149;
srom_1(58855) <= 4791084;
srom_1(58856) <= 4280889;
srom_1(58857) <= 3789956;
srom_1(58858) <= 3320588;
srom_1(58859) <= 2874986;
srom_1(58860) <= 2455239;
srom_1(58861) <= 2063316;
srom_1(58862) <= 1701054;
srom_1(58863) <= 1370152;
srom_1(58864) <= 1072162;
srom_1(58865) <= 808482;
srom_1(58866) <= 580347;
srom_1(58867) <= 388828;
srom_1(58868) <= 234823;
srom_1(58869) <= 119054;
srom_1(58870) <= 42063;
srom_1(58871) <= 4212;
srom_1(58872) <= 5679;
srom_1(58873) <= 46456;
srom_1(58874) <= 126352;
srom_1(58875) <= 244992;
srom_1(58876) <= 401821;
srom_1(58877) <= 596103;
srom_1(58878) <= 826926;
srom_1(58879) <= 1093209;
srom_1(58880) <= 1393702;
srom_1(58881) <= 1726997;
srom_1(58882) <= 2091531;
srom_1(58883) <= 2485593;
srom_1(58884) <= 2907337;
srom_1(58885) <= 3354784;
srom_1(58886) <= 3825837;
srom_1(58887) <= 4318286;
srom_1(58888) <= 4829823;
srom_1(58889) <= 5358047;
srom_1(58890) <= 5900483;
srom_1(58891) <= 6454587;
srom_1(58892) <= 7017760;
srom_1(58893) <= 7587361;
srom_1(58894) <= 8160719;
srom_1(58895) <= 8735147;
srom_1(58896) <= 9307949;
srom_1(58897) <= 9876440;
srom_1(58898) <= 10437954;
srom_1(58899) <= 10989858;
srom_1(58900) <= 11529564;
srom_1(58901) <= 12054540;
srom_1(58902) <= 12562326;
srom_1(58903) <= 13050540;
srom_1(58904) <= 13516893;
srom_1(58905) <= 13959197;
srom_1(58906) <= 14375379;
srom_1(58907) <= 14763487;
srom_1(58908) <= 15121701;
srom_1(58909) <= 15448341;
srom_1(58910) <= 15741875;
srom_1(58911) <= 16000928;
srom_1(58912) <= 16224283;
srom_1(58913) <= 16410895;
srom_1(58914) <= 16559887;
srom_1(58915) <= 16670562;
srom_1(58916) <= 16742399;
srom_1(58917) <= 16775063;
srom_1(58918) <= 16768399;
srom_1(58919) <= 16722440;
srom_1(58920) <= 16637401;
srom_1(58921) <= 16513680;
srom_1(58922) <= 16351858;
srom_1(58923) <= 16152694;
srom_1(58924) <= 15917121;
srom_1(58925) <= 15646244;
srom_1(58926) <= 15341334;
srom_1(58927) <= 15003820;
srom_1(58928) <= 14635285;
srom_1(58929) <= 14237457;
srom_1(58930) <= 13812202;
srom_1(58931) <= 13361514;
srom_1(58932) <= 12887506;
srom_1(58933) <= 12392401;
srom_1(58934) <= 11878521;
srom_1(58935) <= 11348276;
srom_1(58936) <= 10804152;
srom_1(58937) <= 10248700;
srom_1(58938) <= 9684526;
srom_1(58939) <= 9114275;
srom_1(58940) <= 8540621;
srom_1(58941) <= 7966254;
srom_1(58942) <= 7393867;
srom_1(58943) <= 6826146;
srom_1(58944) <= 6265751;
srom_1(58945) <= 5715311;
srom_1(58946) <= 5177407;
srom_1(58947) <= 4654561;
srom_1(58948) <= 4149226;
srom_1(58949) <= 3663771;
srom_1(58950) <= 3200472;
srom_1(58951) <= 2761502;
srom_1(58952) <= 2348919;
srom_1(58953) <= 1964658;
srom_1(58954) <= 1610522;
srom_1(58955) <= 1288170;
srom_1(58956) <= 999115;
srom_1(58957) <= 744712;
srom_1(58958) <= 526153;
srom_1(58959) <= 344464;
srom_1(58960) <= 200497;
srom_1(58961) <= 94927;
srom_1(58962) <= 28249;
srom_1(58963) <= 775;
srom_1(58964) <= 12635;
srom_1(58965) <= 63772;
srom_1(58966) <= 153948;
srom_1(58967) <= 282739;
srom_1(58968) <= 449541;
srom_1(58969) <= 653571;
srom_1(58970) <= 893875;
srom_1(58971) <= 1169323;
srom_1(58972) <= 1478625;
srom_1(58973) <= 1820331;
srom_1(58974) <= 2192837;
srom_1(58975) <= 2594398;
srom_1(58976) <= 3023129;
srom_1(58977) <= 3477021;
srom_1(58978) <= 3953945;
srom_1(58979) <= 4451665;
srom_1(58980) <= 4967847;
srom_1(58981) <= 5500069;
srom_1(58982) <= 6045837;
srom_1(58983) <= 6602591;
srom_1(58984) <= 7167721;
srom_1(58985) <= 7738575;
srom_1(58986) <= 8312478;
srom_1(58987) <= 8886737;
srom_1(58988) <= 9458661;
srom_1(58989) <= 10025567;
srom_1(58990) <= 10584797;
srom_1(58991) <= 11133727;
srom_1(58992) <= 11669786;
srom_1(58993) <= 12190457;
srom_1(58994) <= 12693300;
srom_1(58995) <= 13175958;
srom_1(58996) <= 13636165;
srom_1(58997) <= 14071765;
srom_1(58998) <= 14480715;
srom_1(58999) <= 14861097;
srom_1(59000) <= 15211127;
srom_1(59001) <= 15529163;
srom_1(59002) <= 15813716;
srom_1(59003) <= 16063449;
srom_1(59004) <= 16277193;
srom_1(59005) <= 16453944;
srom_1(59006) <= 16592874;
srom_1(59007) <= 16693331;
srom_1(59008) <= 16754845;
srom_1(59009) <= 16777127;
srom_1(59010) <= 16760071;
srom_1(59011) <= 16703760;
srom_1(59012) <= 16608455;
srom_1(59013) <= 16474605;
srom_1(59014) <= 16302837;
srom_1(59015) <= 16093956;
srom_1(59016) <= 15848943;
srom_1(59017) <= 15568945;
srom_1(59018) <= 15255276;
srom_1(59019) <= 14909407;
srom_1(59020) <= 14532960;
srom_1(59021) <= 14127699;
srom_1(59022) <= 13695527;
srom_1(59023) <= 13238468;
srom_1(59024) <= 12758666;
srom_1(59025) <= 12258372;
srom_1(59026) <= 11739931;
srom_1(59027) <= 11205775;
srom_1(59028) <= 10658408;
srom_1(59029) <= 10100397;
srom_1(59030) <= 9534359;
srom_1(59031) <= 8962948;
srom_1(59032) <= 8388844;
srom_1(59033) <= 7814738;
srom_1(59034) <= 7243324;
srom_1(59035) <= 6677280;
srom_1(59036) <= 6119262;
srom_1(59037) <= 5571885;
srom_1(59038) <= 5037716;
srom_1(59039) <= 4519262;
srom_1(59040) <= 4018951;
srom_1(59041) <= 3539132;
srom_1(59042) <= 3082054;
srom_1(59043) <= 2649859;
srom_1(59044) <= 2244576;
srom_1(59045) <= 1868104;
srom_1(59046) <= 1522209;
srom_1(59047) <= 1208513;
srom_1(59048) <= 928487;
srom_1(59049) <= 683444;
srom_1(59050) <= 474533;
srom_1(59051) <= 302734;
srom_1(59052) <= 168852;
srom_1(59053) <= 73516;
srom_1(59054) <= 17172;
srom_1(59055) <= 84;
srom_1(59056) <= 22333;
srom_1(59057) <= 83815;
srom_1(59058) <= 184240;
srom_1(59059) <= 323139;
srom_1(59060) <= 499859;
srom_1(59061) <= 713572;
srom_1(59062) <= 963277;
srom_1(59063) <= 1247801;
srom_1(59064) <= 1565811;
srom_1(59065) <= 1915815;
srom_1(59066) <= 2296172;
srom_1(59067) <= 2705099;
srom_1(59068) <= 3140678;
srom_1(59069) <= 3600866;
srom_1(59070) <= 4083506;
srom_1(59071) <= 4586333;
srom_1(59072) <= 5106991;
srom_1(59073) <= 5643037;
srom_1(59074) <= 6191959;
srom_1(59075) <= 6751181;
srom_1(59076) <= 7318082;
srom_1(59077) <= 7890002;
srom_1(59078) <= 8464261;
srom_1(59079) <= 9038165;
srom_1(59080) <= 9609023;
srom_1(59081) <= 10174158;
srom_1(59082) <= 10730920;
srom_1(59083) <= 11276698;
srom_1(59084) <= 11808933;
srom_1(59085) <= 12325129;
srom_1(59086) <= 12822865;
srom_1(59087) <= 13299807;
srom_1(59088) <= 13753719;
srom_1(59089) <= 14182472;
srom_1(59090) <= 14584056;
srom_1(59091) <= 14956587;
srom_1(59092) <= 15298319;
srom_1(59093) <= 15607648;
srom_1(59094) <= 15883125;
srom_1(59095) <= 16123458;
srom_1(59096) <= 16327519;
srom_1(59097) <= 16494352;
srom_1(59098) <= 16623175;
srom_1(59099) <= 16713382;
srom_1(59100) <= 16764552;
srom_1(59101) <= 16776444;
srom_1(59102) <= 16749003;
srom_1(59103) <= 16682357;
srom_1(59104) <= 16576819;
srom_1(59105) <= 16432883;
srom_1(59106) <= 16251225;
srom_1(59107) <= 16032697;
srom_1(59108) <= 15778322;
srom_1(59109) <= 15489295;
srom_1(59110) <= 15166970;
srom_1(59111) <= 14812860;
srom_1(59112) <= 14428623;
srom_1(59113) <= 14016063;
srom_1(59114) <= 13577114;
srom_1(59115) <= 13113834;
srom_1(59116) <= 12628396;
srom_1(59117) <= 12123076;
srom_1(59118) <= 11600244;
srom_1(59119) <= 11062351;
srom_1(59120) <= 10511921;
srom_1(59121) <= 9951533;
srom_1(59122) <= 9383816;
srom_1(59123) <= 8811433;
srom_1(59124) <= 8237066;
srom_1(59125) <= 7663411;
srom_1(59126) <= 7093156;
srom_1(59127) <= 6528975;
srom_1(59128) <= 5973515;
srom_1(59129) <= 5429381;
srom_1(59130) <= 4899123;
srom_1(59131) <= 4385229;
srom_1(59132) <= 3890107;
srom_1(59133) <= 3416081;
srom_1(59134) <= 2965373;
srom_1(59135) <= 2540096;
srom_1(59136) <= 2142245;
srom_1(59137) <= 1773685;
srom_1(59138) <= 1436145;
srom_1(59139) <= 1131207;
srom_1(59140) <= 860302;
srom_1(59141) <= 624699;
srom_1(59142) <= 425504;
srom_1(59143) <= 263651;
srom_1(59144) <= 139898;
srom_1(59145) <= 54827;
srom_1(59146) <= 8836;
srom_1(59147) <= 2140;
srom_1(59148) <= 34771;
srom_1(59149) <= 106576;
srom_1(59150) <= 217219;
srom_1(59151) <= 366179;
srom_1(59152) <= 552760;
srom_1(59153) <= 776086;
srom_1(59154) <= 1035110;
srom_1(59155) <= 1328616;
srom_1(59156) <= 1655229;
srom_1(59157) <= 2013418;
srom_1(59158) <= 2401502;
srom_1(59159) <= 2817661;
srom_1(59160) <= 3259945;
srom_1(59161) <= 3726278;
srom_1(59162) <= 4214475;
srom_1(59163) <= 4722246;
srom_1(59164) <= 5247210;
srom_1(59165) <= 5786904;
srom_1(59166) <= 6338799;
srom_1(59167) <= 6900307;
srom_1(59168) <= 7468793;
srom_1(59169) <= 8041593;
srom_1(59170) <= 8616020;
srom_1(59171) <= 9189380;
srom_1(59172) <= 9758986;
srom_1(59173) <= 10322165;
srom_1(59174) <= 10876277;
srom_1(59175) <= 11418724;
srom_1(59176) <= 11946961;
srom_1(59177) <= 12458512;
srom_1(59178) <= 12950978;
srom_1(59179) <= 13422049;
srom_1(59180) <= 13869517;
srom_1(59181) <= 14291283;
srom_1(59182) <= 14685369;
srom_1(59183) <= 15049928;
srom_1(59184) <= 15383249;
srom_1(59185) <= 15683770;
srom_1(59186) <= 15950081;
srom_1(59187) <= 16180934;
srom_1(59188) <= 16375247;
srom_1(59189) <= 16532107;
srom_1(59190) <= 16650779;
srom_1(59191) <= 16730708;
srom_1(59192) <= 16771517;
srom_1(59193) <= 16773016;
srom_1(59194) <= 16735197;
srom_1(59195) <= 16658239;
srom_1(59196) <= 16542501;
srom_1(59197) <= 16388527;
srom_1(59198) <= 16197039;
srom_1(59199) <= 15968934;
srom_1(59200) <= 15705283;
srom_1(59201) <= 15407321;
srom_1(59202) <= 15076446;
srom_1(59203) <= 14714209;
srom_1(59204) <= 14322309;
srom_1(59205) <= 13902584;
srom_1(59206) <= 13457003;
srom_1(59207) <= 12987653;
srom_1(59208) <= 12496738;
srom_1(59209) <= 11986558;
srom_1(59210) <= 11459505;
srom_1(59211) <= 10918053;
srom_1(59212) <= 10364739;
srom_1(59213) <= 9802158;
srom_1(59214) <= 9232948;
srom_1(59215) <= 8659779;
srom_1(59216) <= 8085339;
srom_1(59217) <= 7512320;
srom_1(59218) <= 6943411;
srom_1(59219) <= 6381279;
srom_1(59220) <= 5828560;
srom_1(59221) <= 5287846;
srom_1(59222) <= 4761672;
srom_1(59223) <= 4252506;
srom_1(59224) <= 3762736;
srom_1(59225) <= 3294658;
srom_1(59226) <= 2850468;
srom_1(59227) <= 2432247;
srom_1(59228) <= 2041959;
srom_1(59229) <= 1681431;
srom_1(59230) <= 1352356;
srom_1(59231) <= 1056277;
srom_1(59232) <= 794581;
srom_1(59233) <= 568496;
srom_1(59234) <= 379082;
srom_1(59235) <= 227228;
srom_1(59236) <= 113645;
srom_1(59237) <= 38867;
srom_1(59238) <= 3243;
srom_1(59239) <= 6941;
srom_1(59240) <= 49943;
srom_1(59241) <= 132049;
srom_1(59242) <= 252872;
srom_1(59243) <= 411847;
srom_1(59244) <= 608227;
srom_1(59245) <= 841092;
srom_1(59246) <= 1109350;
srom_1(59247) <= 1411743;
srom_1(59248) <= 1746853;
srom_1(59249) <= 2113108;
srom_1(59250) <= 2508791;
srom_1(59251) <= 2932047;
srom_1(59252) <= 3380891;
srom_1(59253) <= 3853217;
srom_1(59254) <= 4346811;
srom_1(59255) <= 4859359;
srom_1(59256) <= 5388457;
srom_1(59257) <= 5931623;
srom_1(59258) <= 6486311;
srom_1(59259) <= 7049920;
srom_1(59260) <= 7619806;
srom_1(59261) <= 8193297;
srom_1(59262) <= 8767704;
srom_1(59263) <= 9340333;
srom_1(59264) <= 9908500;
srom_1(59265) <= 10469539;
srom_1(59266) <= 11020820;
srom_1(59267) <= 11559757;
srom_1(59268) <= 12083824;
srom_1(59269) <= 12590563;
srom_1(59270) <= 13077597;
srom_1(59271) <= 13542643;
srom_1(59272) <= 13983520;
srom_1(59273) <= 14398161;
srom_1(59274) <= 14784620;
srom_1(59275) <= 15141087;
srom_1(59276) <= 15465889;
srom_1(59277) <= 15757503;
srom_1(59278) <= 16014562;
srom_1(59279) <= 16235860;
srom_1(59280) <= 16420359;
srom_1(59281) <= 16567195;
srom_1(59282) <= 16675679;
srom_1(59283) <= 16745302;
srom_1(59284) <= 16775737;
srom_1(59285) <= 16766842;
srom_1(59286) <= 16718659;
srom_1(59287) <= 16631414;
srom_1(59288) <= 16505515;
srom_1(59289) <= 16341553;
srom_1(59290) <= 16140297;
srom_1(59291) <= 15902690;
srom_1(59292) <= 15629848;
srom_1(59293) <= 15323048;
srom_1(59294) <= 14983731;
srom_1(59295) <= 14613487;
srom_1(59296) <= 14214053;
srom_1(59297) <= 13787300;
srom_1(59298) <= 13335232;
srom_1(59299) <= 12859967;
srom_1(59300) <= 12363734;
srom_1(59301) <= 11848861;
srom_1(59302) <= 11317761;
srom_1(59303) <= 10772926;
srom_1(59304) <= 10216910;
srom_1(59305) <= 9652320;
srom_1(59306) <= 9081804;
srom_1(59307) <= 8508037;
srom_1(59308) <= 7933711;
srom_1(59309) <= 7361517;
srom_1(59310) <= 6794140;
srom_1(59311) <= 6234240;
srom_1(59312) <= 5684442;
srom_1(59313) <= 5147326;
srom_1(59314) <= 4625408;
srom_1(59315) <= 4121138;
srom_1(59316) <= 3636879;
srom_1(59317) <= 3174903;
srom_1(59318) <= 2737376;
srom_1(59319) <= 2326349;
srom_1(59320) <= 1943750;
srom_1(59321) <= 1591373;
srom_1(59322) <= 1270871;
srom_1(59323) <= 983747;
srom_1(59324) <= 731346;
srom_1(59325) <= 514853;
srom_1(59326) <= 335282;
srom_1(59327) <= 193477;
srom_1(59328) <= 90101;
srom_1(59329) <= 25640;
srom_1(59330) <= 395;
srom_1(59331) <= 14486;
srom_1(59332) <= 67846;
srom_1(59333) <= 160225;
srom_1(59334) <= 291189;
srom_1(59335) <= 460125;
srom_1(59336) <= 666241;
srom_1(59337) <= 908569;
srom_1(59338) <= 1185974;
srom_1(59339) <= 1497154;
srom_1(59340) <= 1840651;
srom_1(59341) <= 2214853;
srom_1(59342) <= 2618006;
srom_1(59343) <= 3048220;
srom_1(59344) <= 3503476;
srom_1(59345) <= 3981641;
srom_1(59346) <= 4480471;
srom_1(59347) <= 4997628;
srom_1(59348) <= 5530686;
srom_1(59349) <= 6077146;
srom_1(59350) <= 6634446;
srom_1(59351) <= 7199971;
srom_1(59352) <= 7771070;
srom_1(59353) <= 8345065;
srom_1(59354) <= 8919264;
srom_1(59355) <= 9490975;
srom_1(59356) <= 10057516;
srom_1(59357) <= 10616231;
srom_1(59358) <= 11164500;
srom_1(59359) <= 11699752;
srom_1(59360) <= 12219477;
srom_1(59361) <= 12721238;
srom_1(59362) <= 13202681;
srom_1(59363) <= 13661550;
srom_1(59364) <= 14095692;
srom_1(59365) <= 14503071;
srom_1(59366) <= 14881778;
srom_1(59367) <= 15230036;
srom_1(59368) <= 15546212;
srom_1(59369) <= 15828824;
srom_1(59370) <= 16076545;
srom_1(59371) <= 16288216;
srom_1(59372) <= 16462842;
srom_1(59373) <= 16599606;
srom_1(59374) <= 16697866;
srom_1(59375) <= 16757160;
srom_1(59376) <= 16777212;
srom_1(59377) <= 16757926;
srom_1(59378) <= 16699394;
srom_1(59379) <= 16601890;
srom_1(59380) <= 16465870;
srom_1(59381) <= 16291974;
srom_1(59382) <= 16081016;
srom_1(59383) <= 15833986;
srom_1(59384) <= 15552042;
srom_1(59385) <= 15236506;
srom_1(59386) <= 14888858;
srom_1(59387) <= 14510727;
srom_1(59388) <= 14103889;
srom_1(59389) <= 13670249;
srom_1(59390) <= 13211842;
srom_1(59391) <= 12730817;
srom_1(59392) <= 12229430;
srom_1(59393) <= 11710032;
srom_1(59394) <= 11175058;
srom_1(59395) <= 10627019;
srom_1(59396) <= 10068482;
srom_1(59397) <= 9502068;
srom_1(59398) <= 8930432;
srom_1(59399) <= 8356256;
srom_1(59400) <= 7782231;
srom_1(59401) <= 7211050;
srom_1(59402) <= 6645391;
srom_1(59403) <= 6087906;
srom_1(59404) <= 5541210;
srom_1(59405) <= 5007867;
srom_1(59406) <= 4490377;
srom_1(59407) <= 3991167;
srom_1(59408) <= 3512578;
srom_1(59409) <= 3056855;
srom_1(59410) <= 2626134;
srom_1(59411) <= 2222435;
srom_1(59412) <= 1847652;
srom_1(59413) <= 1503541;
srom_1(59414) <= 1191717;
srom_1(59415) <= 913641;
srom_1(59416) <= 670618;
srom_1(59417) <= 463788;
srom_1(59418) <= 294119;
srom_1(59419) <= 162409;
srom_1(59420) <= 69274;
srom_1(59421) <= 15151;
srom_1(59422) <= 294;
srom_1(59423) <= 24773;
srom_1(59424) <= 88473;
srom_1(59425) <= 191094;
srom_1(59426) <= 332157;
srom_1(59427) <= 511000;
srom_1(59428) <= 726783;
srom_1(59429) <= 978495;
srom_1(59430) <= 1264955;
srom_1(59431) <= 1584821;
srom_1(59432) <= 1936592;
srom_1(59433) <= 2318619;
srom_1(59434) <= 2729110;
srom_1(59435) <= 3166141;
srom_1(59436) <= 3627661;
srom_1(59437) <= 4111507;
srom_1(59438) <= 4615410;
srom_1(59439) <= 5137007;
srom_1(59440) <= 5673851;
srom_1(59441) <= 6223426;
srom_1(59442) <= 6783154;
srom_1(59443) <= 7350411;
srom_1(59444) <= 7922536;
srom_1(59445) <= 8496847;
srom_1(59446) <= 9070650;
srom_1(59447) <= 9641255;
srom_1(59448) <= 10205986;
srom_1(59449) <= 10762194;
srom_1(59450) <= 11307272;
srom_1(59451) <= 11838663;
srom_1(59452) <= 12353876;
srom_1(59453) <= 12850494;
srom_1(59454) <= 13326189;
srom_1(59455) <= 13778730;
srom_1(59456) <= 14205995;
srom_1(59457) <= 14605980;
srom_1(59458) <= 14976809;
srom_1(59459) <= 15316745;
srom_1(59460) <= 15624192;
srom_1(59461) <= 15897708;
srom_1(59462) <= 16136012;
srom_1(59463) <= 16337986;
srom_1(59464) <= 16502682;
srom_1(59465) <= 16629329;
srom_1(59466) <= 16717332;
srom_1(59467) <= 16766279;
srom_1(59468) <= 16775940;
srom_1(59469) <= 16746270;
srom_1(59470) <= 16677408;
srom_1(59471) <= 16569677;
srom_1(59472) <= 16423582;
srom_1(59473) <= 16239808;
srom_1(59474) <= 16019217;
srom_1(59475) <= 15762844;
srom_1(59476) <= 15471891;
srom_1(59477) <= 15147721;
srom_1(59478) <= 14791856;
srom_1(59479) <= 14405963;
srom_1(59480) <= 13991854;
srom_1(59481) <= 13551468;
srom_1(59482) <= 13086873;
srom_1(59483) <= 12600245;
srom_1(59484) <= 12093868;
srom_1(59485) <= 11570115;
srom_1(59486) <= 11031443;
srom_1(59487) <= 10480378;
srom_1(59488) <= 9919504;
srom_1(59489) <= 9351451;
srom_1(59490) <= 8778883;
srom_1(59491) <= 8204485;
srom_1(59492) <= 7630950;
srom_1(59493) <= 7060968;
srom_1(59494) <= 6497212;
srom_1(59495) <= 5942326;
srom_1(59496) <= 5398910;
srom_1(59497) <= 4869515;
srom_1(59498) <= 4356622;
srom_1(59499) <= 3862636;
srom_1(59500) <= 3389874;
srom_1(59501) <= 2940552;
srom_1(59502) <= 2516779;
srom_1(59503) <= 2120540;
srom_1(59504) <= 1753695;
srom_1(59505) <= 1417963;
srom_1(59506) <= 1114918;
srom_1(59507) <= 845983;
srom_1(59508) <= 612417;
srom_1(59509) <= 415317;
srom_1(59510) <= 255606;
srom_1(59511) <= 134034;
srom_1(59512) <= 51170;
srom_1(59513) <= 7403;
srom_1(59514) <= 2939;
srom_1(59515) <= 37798;
srom_1(59516) <= 111817;
srom_1(59517) <= 224648;
srom_1(59518) <= 375763;
srom_1(59519) <= 564453;
srom_1(59520) <= 789833;
srom_1(59521) <= 1050847;
srom_1(59522) <= 1346269;
srom_1(59523) <= 1674716;
srom_1(59524) <= 2034646;
srom_1(59525) <= 2424372;
srom_1(59526) <= 2842067;
srom_1(59527) <= 3285771;
srom_1(59528) <= 3753404;
srom_1(59529) <= 4242774;
srom_1(59530) <= 4751584;
srom_1(59531) <= 5277450;
srom_1(59532) <= 5817905;
srom_1(59533) <= 6370415;
srom_1(59534) <= 6932389;
srom_1(59535) <= 7501191;
srom_1(59536) <= 8074155;
srom_1(59537) <= 8648594;
srom_1(59538) <= 9221813;
srom_1(59539) <= 9791125;
srom_1(59540) <= 10353861;
srom_1(59541) <= 10907380;
srom_1(59542) <= 11449088;
srom_1(59543) <= 11976445;
srom_1(59544) <= 12486977;
srom_1(59545) <= 12978290;
srom_1(59546) <= 13448081;
srom_1(59547) <= 13894146;
srom_1(59548) <= 14314393;
srom_1(59549) <= 14706853;
srom_1(59550) <= 15069684;
srom_1(59551) <= 15401185;
srom_1(59552) <= 15699802;
srom_1(59553) <= 15964135;
srom_1(59554) <= 16192942;
srom_1(59555) <= 16385153;
srom_1(59556) <= 16539865;
srom_1(59557) <= 16656354;
srom_1(59558) <= 16734071;
srom_1(59559) <= 16772654;
srom_1(59560) <= 16771922;
srom_1(59561) <= 16731877;
srom_1(59562) <= 16652708;
srom_1(59563) <= 16534785;
srom_1(59564) <= 16378662;
srom_1(59565) <= 16185071;
srom_1(59566) <= 15954920;
srom_1(59567) <= 15689288;
srom_1(59568) <= 15389420;
srom_1(59569) <= 15056724;
srom_1(59570) <= 14692758;
srom_1(59571) <= 14299229;
srom_1(59572) <= 13877984;
srom_1(59573) <= 13430997;
srom_1(59574) <= 12960365;
srom_1(59575) <= 12468294;
srom_1(59576) <= 11957092;
srom_1(59577) <= 11429157;
srom_1(59578) <= 10886963;
srom_1(59579) <= 10333053;
srom_1(59580) <= 9770025;
srom_1(59581) <= 9200520;
srom_1(59582) <= 8627207;
srom_1(59583) <= 8052775;
srom_1(59584) <= 7479918;
srom_1(59585) <= 6911322;
srom_1(59586) <= 6349653;
srom_1(59587) <= 5797546;
srom_1(59588) <= 5257589;
srom_1(59589) <= 4732315;
srom_1(59590) <= 4224186;
srom_1(59591) <= 3735586;
srom_1(59592) <= 3268805;
srom_1(59593) <= 2826033;
srom_1(59594) <= 2409346;
srom_1(59595) <= 2020697;
srom_1(59596) <= 1661910;
srom_1(59597) <= 1334667;
srom_1(59598) <= 1040501;
srom_1(59599) <= 780794;
srom_1(59600) <= 556762;
srom_1(59601) <= 369457;
srom_1(59602) <= 219756;
srom_1(59603) <= 108362;
srom_1(59604) <= 35796;
srom_1(59605) <= 2400;
srom_1(59606) <= 8329;
srom_1(59607) <= 53557;
srom_1(59608) <= 137870;
srom_1(59609) <= 260874;
srom_1(59610) <= 421992;
srom_1(59611) <= 620468;
srom_1(59612) <= 855371;
srom_1(59613) <= 1125601;
srom_1(59614) <= 1429889;
srom_1(59615) <= 1766809;
srom_1(59616) <= 2134780;
srom_1(59617) <= 2532078;
srom_1(59618) <= 2956840;
srom_1(59619) <= 3407073;
srom_1(59620) <= 3880665;
srom_1(59621) <= 4375398;
srom_1(59622) <= 4888949;
srom_1(59623) <= 5418912;
srom_1(59624) <= 5962800;
srom_1(59625) <= 6518064;
srom_1(59626) <= 7082100;
srom_1(59627) <= 7652262;
srom_1(59628) <= 8225877;
srom_1(59629) <= 8800255;
srom_1(59630) <= 9372703;
srom_1(59631) <= 9940537;
srom_1(59632) <= 10501092;
srom_1(59633) <= 11051742;
srom_1(59634) <= 11589903;
srom_1(59635) <= 12113052;
srom_1(59636) <= 12618736;
srom_1(59637) <= 13104583;
srom_1(59638) <= 13568316;
srom_1(59639) <= 14007759;
srom_1(59640) <= 14420852;
srom_1(59641) <= 14805657;
srom_1(59642) <= 15160371;
srom_1(59643) <= 15483330;
srom_1(59644) <= 15773019;
srom_1(59645) <= 16028081;
srom_1(59646) <= 16247318;
srom_1(59647) <= 16429703;
srom_1(59648) <= 16574380;
srom_1(59649) <= 16680671;
srom_1(59650) <= 16748079;
srom_1(59651) <= 16776285;
srom_1(59652) <= 16765159;
srom_1(59653) <= 16714753;
srom_1(59654) <= 16625302;
srom_1(59655) <= 16497227;
srom_1(59656) <= 16331127;
srom_1(59657) <= 16127782;
srom_1(59658) <= 15888146;
srom_1(59659) <= 15613342;
srom_1(59660) <= 15304658;
srom_1(59661) <= 14963543;
srom_1(59662) <= 14591596;
srom_1(59663) <= 14190560;
srom_1(59664) <= 13762318;
srom_1(59665) <= 13308876;
srom_1(59666) <= 12832361;
srom_1(59667) <= 12335008;
srom_1(59668) <= 11819149;
srom_1(59669) <= 11287203;
srom_1(59670) <= 10741664;
srom_1(59671) <= 10185091;
srom_1(59672) <= 9620094;
srom_1(59673) <= 9049322;
srom_1(59674) <= 8475452;
srom_1(59675) <= 7901174;
srom_1(59676) <= 7329182;
srom_1(59677) <= 6762158;
srom_1(59678) <= 6202761;
srom_1(59679) <= 5653615;
srom_1(59680) <= 5117293;
srom_1(59681) <= 4596312;
srom_1(59682) <= 4093114;
srom_1(59683) <= 3610060;
srom_1(59684) <= 3149413;
srom_1(59685) <= 2713335;
srom_1(59686) <= 2303870;
srom_1(59687) <= 1922939;
srom_1(59688) <= 1572328;
srom_1(59689) <= 1253680;
srom_1(59690) <= 968490;
srom_1(59691) <= 718096;
srom_1(59692) <= 503671;
srom_1(59693) <= 326222;
srom_1(59694) <= 186580;
srom_1(59695) <= 85400;
srom_1(59696) <= 23157;
srom_1(59697) <= 142;
srom_1(59698) <= 16464;
srom_1(59699) <= 72045;
srom_1(59700) <= 166626;
srom_1(59701) <= 299762;
srom_1(59702) <= 470830;
srom_1(59703) <= 679026;
srom_1(59704) <= 923376;
srom_1(59705) <= 1202733;
srom_1(59706) <= 1515787;
srom_1(59707) <= 1861069;
srom_1(59708) <= 2236962;
srom_1(59709) <= 2641702;
srom_1(59710) <= 3073391;
srom_1(59711) <= 3530005;
srom_1(59712) <= 4009402;
srom_1(59713) <= 4509336;
srom_1(59714) <= 5027460;
srom_1(59715) <= 5561346;
srom_1(59716) <= 6108490;
srom_1(59717) <= 6666326;
srom_1(59718) <= 7232239;
srom_1(59719) <= 7803574;
srom_1(59720) <= 8377652;
srom_1(59721) <= 8951782;
srom_1(59722) <= 9523271;
srom_1(59723) <= 10089440;
srom_1(59724) <= 10647632;
srom_1(59725) <= 11195231;
srom_1(59726) <= 11729669;
srom_1(59727) <= 12248439;
srom_1(59728) <= 12749110;
srom_1(59729) <= 13229332;
srom_1(59730) <= 13686855;
srom_1(59731) <= 14119532;
srom_1(59732) <= 14525335;
srom_1(59733) <= 14902361;
srom_1(59734) <= 15248842;
srom_1(59735) <= 15563152;
srom_1(59736) <= 15843819;
srom_1(59737) <= 16089526;
srom_1(59738) <= 16299120;
srom_1(59739) <= 16471619;
srom_1(59740) <= 16606214;
srom_1(59741) <= 16702275;
srom_1(59742) <= 16759349;
srom_1(59743) <= 16777170;
srom_1(59744) <= 16755654;
srom_1(59745) <= 16694903;
srom_1(59746) <= 16595200;
srom_1(59747) <= 16457014;
srom_1(59748) <= 16280992;
srom_1(59749) <= 16067960;
srom_1(59750) <= 15818917;
srom_1(59751) <= 15535030;
srom_1(59752) <= 15217632;
srom_1(59753) <= 14868210;
srom_1(59754) <= 14488403;
srom_1(59755) <= 14079992;
srom_1(59756) <= 13644892;
srom_1(59757) <= 13185143;
srom_1(59758) <= 12702902;
srom_1(59759) <= 12200430;
srom_1(59760) <= 11680082;
srom_1(59761) <= 11144300;
srom_1(59762) <= 10595595;
srom_1(59763) <= 10036542;
srom_1(59764) <= 9469760;
srom_1(59765) <= 8897908;
srom_1(59766) <= 8323669;
srom_1(59767) <= 7749733;
srom_1(59768) <= 7178794;
srom_1(59769) <= 6613528;
srom_1(59770) <= 6056585;
srom_1(59771) <= 5510579;
srom_1(59772) <= 4978068;
srom_1(59773) <= 4461551;
srom_1(59774) <= 3963449;
srom_1(59775) <= 3486098;
srom_1(59776) <= 3031737;
srom_1(59777) <= 2602495;
srom_1(59778) <= 2200387;
srom_1(59779) <= 1827298;
srom_1(59780) <= 1484977;
srom_1(59781) <= 1175029;
srom_1(59782) <= 898908;
srom_1(59783) <= 657909;
srom_1(59784) <= 453162;
srom_1(59785) <= 285627;
srom_1(59786) <= 156089;
srom_1(59787) <= 65157;
srom_1(59788) <= 13256;
srom_1(59789) <= 630;
srom_1(59790) <= 27339;
srom_1(59791) <= 93256;
srom_1(59792) <= 198072;
srom_1(59793) <= 341297;
srom_1(59794) <= 522259;
srom_1(59795) <= 740109;
srom_1(59796) <= 993825;
srom_1(59797) <= 1282217;
srom_1(59798) <= 1603934;
srom_1(59799) <= 1957467;
srom_1(59800) <= 2341158;
srom_1(59801) <= 2753207;
srom_1(59802) <= 3191682;
srom_1(59803) <= 3654528;
srom_1(59804) <= 4139573;
srom_1(59805) <= 4644543;
srom_1(59806) <= 5167071;
srom_1(59807) <= 5704706;
srom_1(59808) <= 6254926;
srom_1(59809) <= 6815152;
srom_1(59810) <= 7382756;
srom_1(59811) <= 7955077;
srom_1(59812) <= 8529431;
srom_1(59813) <= 9103125;
srom_1(59814) <= 9673468;
srom_1(59815) <= 10237786;
srom_1(59816) <= 10793432;
srom_1(59817) <= 11337802;
srom_1(59818) <= 11868341;
srom_1(59819) <= 12382563;
srom_1(59820) <= 12878056;
srom_1(59821) <= 13352497;
srom_1(59822) <= 13803659;
srom_1(59823) <= 14229429;
srom_1(59824) <= 14627810;
srom_1(59825) <= 14996932;
srom_1(59826) <= 15335066;
srom_1(59827) <= 15640625;
srom_1(59828) <= 15912178;
srom_1(59829) <= 16148449;
srom_1(59830) <= 16348332;
srom_1(59831) <= 16510890;
srom_1(59832) <= 16635359;
srom_1(59833) <= 16721156;
srom_1(59834) <= 16767879;
srom_1(59835) <= 16775309;
srom_1(59836) <= 16743410;
srom_1(59837) <= 16672333;
srom_1(59838) <= 16562411;
srom_1(59839) <= 16414159;
srom_1(59840) <= 16228272;
srom_1(59841) <= 16005623;
srom_1(59842) <= 15747255;
srom_1(59843) <= 15454379;
srom_1(59844) <= 15128370;
srom_1(59845) <= 14770755;
srom_1(59846) <= 14383213;
srom_1(59847) <= 13967560;
srom_1(59848) <= 13525745;
srom_1(59849) <= 13059840;
srom_1(59850) <= 12572030;
srom_1(59851) <= 12064603;
srom_1(59852) <= 11539938;
srom_1(59853) <= 11000495;
srom_1(59854) <= 10448804;
srom_1(59855) <= 9887452;
srom_1(59856) <= 9319072;
srom_1(59857) <= 8746328;
srom_1(59858) <= 8171907;
srom_1(59859) <= 7598502;
srom_1(59860) <= 7028801;
srom_1(59861) <= 6465478;
srom_1(59862) <= 5911173;
srom_1(59863) <= 5368485;
srom_1(59864) <= 4839960;
srom_1(59865) <= 4328075;
srom_1(59866) <= 3835232;
srom_1(59867) <= 3363741;
srom_1(59868) <= 2915814;
srom_1(59869) <= 2493550;
srom_1(59870) <= 2098930;
srom_1(59871) <= 1733805;
srom_1(59872) <= 1399886;
srom_1(59873) <= 1098740;
srom_1(59874) <= 831778;
srom_1(59875) <= 600253;
srom_1(59876) <= 405251;
srom_1(59877) <= 247685;
srom_1(59878) <= 128294;
srom_1(59879) <= 47639;
srom_1(59880) <= 6098;
srom_1(59881) <= 3865;
srom_1(59882) <= 40951;
srom_1(59883) <= 117182;
srom_1(59884) <= 232201;
srom_1(59885) <= 385468;
srom_1(59886) <= 576264;
srom_1(59887) <= 803695;
srom_1(59888) <= 1066694;
srom_1(59889) <= 1364029;
srom_1(59890) <= 1694304;
srom_1(59891) <= 2055970;
srom_1(59892) <= 2447333;
srom_1(59893) <= 2866557;
srom_1(59894) <= 3311675;
srom_1(59895) <= 3780600;
srom_1(59896) <= 4271135;
srom_1(59897) <= 4780977;
srom_1(59898) <= 5307737;
srom_1(59899) <= 5848944;
srom_1(59900) <= 6402061;
srom_1(59901) <= 6964493;
srom_1(59902) <= 7533603;
srom_1(59903) <= 8106722;
srom_1(59904) <= 8681164;
srom_1(59905) <= 9254233;
srom_1(59906) <= 9823244;
srom_1(59907) <= 10385527;
srom_1(59908) <= 10938445;
srom_1(59909) <= 11479407;
srom_1(59910) <= 12005874;
srom_1(59911) <= 12515380;
srom_1(59912) <= 13005533;
srom_1(59913) <= 13474036;
srom_1(59914) <= 13918691;
srom_1(59915) <= 14337414;
srom_1(59916) <= 14728241;
srom_1(59917) <= 15089340;
srom_1(59918) <= 15419016;
srom_1(59919) <= 15715724;
srom_1(59920) <= 15978073;
srom_1(59921) <= 16204833;
srom_1(59922) <= 16394939;
srom_1(59923) <= 16547501;
srom_1(59924) <= 16661803;
srom_1(59925) <= 16737309;
srom_1(59926) <= 16773665;
srom_1(59927) <= 16770701;
srom_1(59928) <= 16728431;
srom_1(59929) <= 16647052;
srom_1(59930) <= 16526946;
srom_1(59931) <= 16368677;
srom_1(59932) <= 16172986;
srom_1(59933) <= 15940792;
srom_1(59934) <= 15673183;
srom_1(59935) <= 15371415;
srom_1(59936) <= 15036901;
srom_1(59937) <= 14671211;
srom_1(59938) <= 14276060;
srom_1(59939) <= 13853301;
srom_1(59940) <= 13404916;
srom_1(59941) <= 12933008;
srom_1(59942) <= 12439789;
srom_1(59943) <= 11927573;
srom_1(59944) <= 11398762;
srom_1(59945) <= 10855835;
srom_1(59946) <= 10301338;
srom_1(59947) <= 9737872;
srom_1(59948) <= 9168079;
srom_1(59949) <= 8594630;
srom_1(59950) <= 8020216;
srom_1(59951) <= 7447528;
srom_1(59952) <= 6879254;
srom_1(59953) <= 6318058;
srom_1(59954) <= 5766571;
srom_1(59955) <= 5227380;
srom_1(59956) <= 4703013;
srom_1(59957) <= 4195929;
srom_1(59958) <= 3708506;
srom_1(59959) <= 3243030;
srom_1(59960) <= 2801682;
srom_1(59961) <= 2386534;
srom_1(59962) <= 1999532;
srom_1(59963) <= 1642490;
srom_1(59964) <= 1317083;
srom_1(59965) <= 1024837;
srom_1(59966) <= 767122;
srom_1(59967) <= 545147;
srom_1(59968) <= 359953;
srom_1(59969) <= 212407;
srom_1(59970) <= 103203;
srom_1(59971) <= 32852;
srom_1(59972) <= 1684;
srom_1(59973) <= 9845;
srom_1(59974) <= 57296;
srom_1(59975) <= 143817;
srom_1(59976) <= 269000;
srom_1(59977) <= 432258;
srom_1(59978) <= 632827;
srom_1(59979) <= 869765;
srom_1(59980) <= 1141961;
srom_1(59981) <= 1448140;
srom_1(59982) <= 1786864;
srom_1(59983) <= 2156547;
srom_1(59984) <= 2555454;
srom_1(59985) <= 2981714;
srom_1(59986) <= 3433330;
srom_1(59987) <= 3908182;
srom_1(59988) <= 4404044;
srom_1(59989) <= 4918592;
srom_1(59990) <= 5449411;
srom_1(59991) <= 5994014;
srom_1(59992) <= 6549846;
srom_1(59993) <= 7114300;
srom_1(59994) <= 7684729;
srom_1(59995) <= 8258460;
srom_1(59996) <= 8832801;
srom_1(59997) <= 9405059;
srom_1(59998) <= 9972550;
srom_1(59999) <= 10532614;
srom_1(60000) <= 11082623;
srom_1(60001) <= 11620000;
srom_1(60002) <= 12142223;
srom_1(60003) <= 12646845;
srom_1(60004) <= 13131498;
srom_1(60005) <= 13593910;
srom_1(60006) <= 14031912;
srom_1(60007) <= 14443452;
srom_1(60008) <= 14826598;
srom_1(60009) <= 15179554;
srom_1(60010) <= 15500664;
srom_1(60011) <= 15788424;
srom_1(60012) <= 16041484;
srom_1(60013) <= 16258657;
srom_1(60014) <= 16438924;
srom_1(60015) <= 16581441;
srom_1(60016) <= 16685539;
srom_1(60017) <= 16750729;
srom_1(60018) <= 16776707;
srom_1(60019) <= 16763350;
srom_1(60020) <= 16710721;
srom_1(60021) <= 16619066;
srom_1(60022) <= 16488816;
srom_1(60023) <= 16320582;
srom_1(60024) <= 16115152;
srom_1(60025) <= 15873489;
srom_1(60026) <= 15596727;
srom_1(60027) <= 15286164;
srom_1(60028) <= 14943256;
srom_1(60029) <= 14569611;
srom_1(60030) <= 14166980;
srom_1(60031) <= 13737254;
srom_1(60032) <= 13282445;
srom_1(60033) <= 12804688;
srom_1(60034) <= 12306222;
srom_1(60035) <= 11789385;
srom_1(60036) <= 11256600;
srom_1(60037) <= 10710367;
srom_1(60038) <= 10153246;
srom_1(60039) <= 9587850;
srom_1(60040) <= 9016831;
srom_1(60041) <= 8442865;
srom_1(60042) <= 7868645;
srom_1(60043) <= 7296863;
srom_1(60044) <= 6730201;
srom_1(60045) <= 6171316;
srom_1(60046) <= 5622828;
srom_1(60047) <= 5087310;
srom_1(60048) <= 4567273;
srom_1(60049) <= 4065156;
srom_1(60050) <= 3583312;
srom_1(60051) <= 3124003;
srom_1(60052) <= 2689380;
srom_1(60053) <= 2281484;
srom_1(60054) <= 1902226;
srom_1(60055) <= 1553384;
srom_1(60056) <= 1236596;
srom_1(60057) <= 953346;
srom_1(60058) <= 704962;
srom_1(60059) <= 492609;
srom_1(60060) <= 317284;
srom_1(60061) <= 179807;
srom_1(60062) <= 80825;
srom_1(60063) <= 20800;
srom_1(60064) <= 15;
srom_1(60065) <= 18567;
srom_1(60066) <= 76370;
srom_1(60067) <= 173151;
srom_1(60068) <= 308457;
srom_1(60069) <= 481653;
srom_1(60070) <= 691928;
srom_1(60071) <= 938296;
srom_1(60072) <= 1219600;
srom_1(60073) <= 1534523;
srom_1(60074) <= 1881587;
srom_1(60075) <= 2259164;
srom_1(60076) <= 2665484;
srom_1(60077) <= 3098642;
srom_1(60078) <= 3556607;
srom_1(60079) <= 4037230;
srom_1(60080) <= 4538259;
srom_1(60081) <= 5057343;
srom_1(60082) <= 5592048;
srom_1(60083) <= 6139868;
srom_1(60084) <= 6698233;
srom_1(60085) <= 7264524;
srom_1(60086) <= 7836087;
srom_1(60087) <= 8410240;
srom_1(60088) <= 8984292;
srom_1(60089) <= 9555551;
srom_1(60090) <= 10121338;
srom_1(60091) <= 10678999;
srom_1(60092) <= 11225920;
srom_1(60093) <= 11759535;
srom_1(60094) <= 12277343;
srom_1(60095) <= 12776916;
srom_1(60096) <= 13255910;
srom_1(60097) <= 13712080;
srom_1(60098) <= 14143286;
srom_1(60099) <= 14547507;
srom_1(60100) <= 14922846;
srom_1(60101) <= 15267544;
srom_1(60102) <= 15579984;
srom_1(60103) <= 15858702;
srom_1(60104) <= 16102390;
srom_1(60105) <= 16309905;
srom_1(60106) <= 16480274;
srom_1(60107) <= 16612699;
srom_1(60108) <= 16706558;
srom_1(60109) <= 16761411;
srom_1(60110) <= 16777002;
srom_1(60111) <= 16753256;
srom_1(60112) <= 16690286;
srom_1(60113) <= 16588386;
srom_1(60114) <= 16448035;
srom_1(60115) <= 16269890;
srom_1(60116) <= 16054787;
srom_1(60117) <= 15803735;
srom_1(60118) <= 15517911;
srom_1(60119) <= 15198655;
srom_1(60120) <= 14847465;
srom_1(60121) <= 14465986;
srom_1(60122) <= 14056009;
srom_1(60123) <= 13619455;
srom_1(60124) <= 13158372;
srom_1(60125) <= 12674922;
srom_1(60126) <= 12171372;
srom_1(60127) <= 11650083;
srom_1(60128) <= 11113500;
srom_1(60129) <= 10564139;
srom_1(60130) <= 10004576;
srom_1(60131) <= 9437436;
srom_1(60132) <= 8865377;
srom_1(60133) <= 8291082;
srom_1(60134) <= 7717245;
srom_1(60135) <= 7146556;
srom_1(60136) <= 6581691;
srom_1(60137) <= 6025300;
srom_1(60138) <= 5479991;
srom_1(60139) <= 4948321;
srom_1(60140) <= 4432784;
srom_1(60141) <= 3935798;
srom_1(60142) <= 3459692;
srom_1(60143) <= 3006699;
srom_1(60144) <= 2578944;
srom_1(60145) <= 2178433;
srom_1(60146) <= 1807043;
srom_1(60147) <= 1466516;
srom_1(60148) <= 1158450;
srom_1(60149) <= 884288;
srom_1(60150) <= 645317;
srom_1(60151) <= 442656;
srom_1(60152) <= 277257;
srom_1(60153) <= 149894;
srom_1(60154) <= 61166;
srom_1(60155) <= 11488;
srom_1(60156) <= 1093;
srom_1(60157) <= 30031;
srom_1(60158) <= 98164;
srom_1(60159) <= 205174;
srom_1(60160) <= 350559;
srom_1(60161) <= 533637;
srom_1(60162) <= 753550;
srom_1(60163) <= 1009266;
srom_1(60164) <= 1299587;
srom_1(60165) <= 1623150;
srom_1(60166) <= 1978439;
srom_1(60167) <= 2363787;
srom_1(60168) <= 2777388;
srom_1(60169) <= 3217302;
srom_1(60170) <= 3681466;
srom_1(60171) <= 4167703;
srom_1(60172) <= 4673733;
srom_1(60173) <= 5197184;
srom_1(60174) <= 5735601;
srom_1(60175) <= 6286458;
srom_1(60176) <= 6847173;
srom_1(60177) <= 7415116;
srom_1(60178) <= 7987625;
srom_1(60179) <= 8562013;
srom_1(60180) <= 9135589;
srom_1(60181) <= 9705661;
srom_1(60182) <= 10269558;
srom_1(60183) <= 10824634;
srom_1(60184) <= 11368287;
srom_1(60185) <= 11897967;
srom_1(60186) <= 12411190;
srom_1(60187) <= 12905550;
srom_1(60188) <= 13378729;
srom_1(60189) <= 13828507;
srom_1(60190) <= 14252776;
srom_1(60191) <= 14649545;
srom_1(60192) <= 15016955;
srom_1(60193) <= 15353282;
srom_1(60194) <= 15656950;
srom_1(60195) <= 15926534;
srom_1(60196) <= 16160769;
srom_1(60197) <= 16358559;
srom_1(60198) <= 16518975;
srom_1(60199) <= 16641264;
srom_1(60200) <= 16724854;
srom_1(60201) <= 16769353;
srom_1(60202) <= 16774551;
srom_1(60203) <= 16740424;
srom_1(60204) <= 16667134;
srom_1(60205) <= 16555022;
srom_1(60206) <= 16404615;
srom_1(60207) <= 16216618;
srom_1(60208) <= 15991913;
srom_1(60209) <= 15731554;
srom_1(60210) <= 15436761;
srom_1(60211) <= 15108917;
srom_1(60212) <= 14749559;
srom_1(60213) <= 14360372;
srom_1(60214) <= 13943181;
srom_1(60215) <= 13499944;
srom_1(60216) <= 13032737;
srom_1(60217) <= 12543753;
srom_1(60218) <= 12035283;
srom_1(60219) <= 11509713;
srom_1(60220) <= 10969507;
srom_1(60221) <= 10417199;
srom_1(60222) <= 9855378;
srom_1(60223) <= 9286678;
srom_1(60224) <= 8713767;
srom_1(60225) <= 8139331;
srom_1(60226) <= 7566065;
srom_1(60227) <= 6996655;
srom_1(60228) <= 6433773;
srom_1(60229) <= 5880057;
srom_1(60230) <= 5338105;
srom_1(60231) <= 4810458;
srom_1(60232) <= 4299591;
srom_1(60233) <= 3807897;
srom_1(60234) <= 3337685;
srom_1(60235) <= 2891158;
srom_1(60236) <= 2470410;
srom_1(60237) <= 2077415;
srom_1(60238) <= 1714015;
srom_1(60239) <= 1381915;
srom_1(60240) <= 1082671;
srom_1(60241) <= 817688;
srom_1(60242) <= 588207;
srom_1(60243) <= 395304;
srom_1(60244) <= 239886;
srom_1(60245) <= 122679;
srom_1(60246) <= 44234;
srom_1(60247) <= 4919;
srom_1(60248) <= 4917;
srom_1(60249) <= 44230;
srom_1(60250) <= 122673;
srom_1(60251) <= 239877;
srom_1(60252) <= 395293;
srom_1(60253) <= 588193;
srom_1(60254) <= 817671;
srom_1(60255) <= 1082653;
srom_1(60256) <= 1381894;
srom_1(60257) <= 1713992;
srom_1(60258) <= 2077390;
srom_1(60259) <= 2470384;
srom_1(60260) <= 2891129;
srom_1(60261) <= 3337655;
srom_1(60262) <= 3807866;
srom_1(60263) <= 4299558;
srom_1(60264) <= 4810425;
srom_1(60265) <= 5338071;
srom_1(60266) <= 5880022;
srom_1(60267) <= 6433736;
srom_1(60268) <= 6996618;
srom_1(60269) <= 7566027;
srom_1(60270) <= 8139294;
srom_1(60271) <= 8713730;
srom_1(60272) <= 9286641;
srom_1(60273) <= 9855341;
srom_1(60274) <= 10417163;
srom_1(60275) <= 10969472;
srom_1(60276) <= 11509679;
srom_1(60277) <= 12035249;
srom_1(60278) <= 12543720;
srom_1(60279) <= 13032706;
srom_1(60280) <= 13499914;
srom_1(60281) <= 13943153;
srom_1(60282) <= 14360346;
srom_1(60283) <= 14749534;
srom_1(60284) <= 15108894;
srom_1(60285) <= 15436741;
srom_1(60286) <= 15731536;
srom_1(60287) <= 15991898;
srom_1(60288) <= 16216605;
srom_1(60289) <= 16404604;
srom_1(60290) <= 16555013;
srom_1(60291) <= 16667128;
srom_1(60292) <= 16740421;
srom_1(60293) <= 16774550;
srom_1(60294) <= 16769354;
srom_1(60295) <= 16724858;
srom_1(60296) <= 16641271;
srom_1(60297) <= 16518984;
srom_1(60298) <= 16358571;
srom_1(60299) <= 16160784;
srom_1(60300) <= 15926550;
srom_1(60301) <= 15656969;
srom_1(60302) <= 15353303;
srom_1(60303) <= 15016978;
srom_1(60304) <= 14649570;
srom_1(60305) <= 14252803;
srom_1(60306) <= 13828536;
srom_1(60307) <= 13378759;
srom_1(60308) <= 12905582;
srom_1(60309) <= 12411223;
srom_1(60310) <= 11898001;
srom_1(60311) <= 11368322;
srom_1(60312) <= 10824670;
srom_1(60313) <= 10269595;
srom_1(60314) <= 9705698;
srom_1(60315) <= 9135626;
srom_1(60316) <= 8562051;
srom_1(60317) <= 7987662;
srom_1(60318) <= 7415153;
srom_1(60319) <= 6847210;
srom_1(60320) <= 6286494;
srom_1(60321) <= 5735636;
srom_1(60322) <= 5197219;
srom_1(60323) <= 4673767;
srom_1(60324) <= 4167735;
srom_1(60325) <= 3681497;
srom_1(60326) <= 3217332;
srom_1(60327) <= 2777416;
srom_1(60328) <= 2363814;
srom_1(60329) <= 1978463;
srom_1(60330) <= 1623172;
srom_1(60331) <= 1299607;
srom_1(60332) <= 1009284;
srom_1(60333) <= 753566;
srom_1(60334) <= 533650;
srom_1(60335) <= 350570;
srom_1(60336) <= 205182;
srom_1(60337) <= 98170;
srom_1(60338) <= 30034;
srom_1(60339) <= 1094;
srom_1(60340) <= 11486;
srom_1(60341) <= 61162;
srom_1(60342) <= 149887;
srom_1(60343) <= 277247;
srom_1(60344) <= 442644;
srom_1(60345) <= 645302;
srom_1(60346) <= 884271;
srom_1(60347) <= 1158431;
srom_1(60348) <= 1466495;
srom_1(60349) <= 1807020;
srom_1(60350) <= 2178408;
srom_1(60351) <= 2578917;
srom_1(60352) <= 3006670;
srom_1(60353) <= 3459661;
srom_1(60354) <= 3935766;
srom_1(60355) <= 4432751;
srom_1(60356) <= 4948287;
srom_1(60357) <= 5479956;
srom_1(60358) <= 6025264;
srom_1(60359) <= 6581655;
srom_1(60360) <= 7146519;
srom_1(60361) <= 7717208;
srom_1(60362) <= 8291045;
srom_1(60363) <= 8865339;
srom_1(60364) <= 9437399;
srom_1(60365) <= 10004540;
srom_1(60366) <= 10564103;
srom_1(60367) <= 11113465;
srom_1(60368) <= 11650048;
srom_1(60369) <= 12171338;
srom_1(60370) <= 12674890;
srom_1(60371) <= 13158341;
srom_1(60372) <= 13619426;
srom_1(60373) <= 14055981;
srom_1(60374) <= 14465960;
srom_1(60375) <= 14847441;
srom_1(60376) <= 15198633;
srom_1(60377) <= 15517891;
srom_1(60378) <= 15803718;
srom_1(60379) <= 16054772;
srom_1(60380) <= 16269877;
srom_1(60381) <= 16448025;
srom_1(60382) <= 16588378;
srom_1(60383) <= 16690281;
srom_1(60384) <= 16753254;
srom_1(60385) <= 16777002;
srom_1(60386) <= 16761414;
srom_1(60387) <= 16706563;
srom_1(60388) <= 16612706;
srom_1(60389) <= 16480284;
srom_1(60390) <= 16309917;
srom_1(60391) <= 16102404;
srom_1(60392) <= 15858719;
srom_1(60393) <= 15580004;
srom_1(60394) <= 15267566;
srom_1(60395) <= 14922870;
srom_1(60396) <= 14547532;
srom_1(60397) <= 14143313;
srom_1(60398) <= 13712109;
srom_1(60399) <= 13255941;
srom_1(60400) <= 12776948;
srom_1(60401) <= 12277377;
srom_1(60402) <= 11759570;
srom_1(60403) <= 11225955;
srom_1(60404) <= 10679035;
srom_1(60405) <= 10121374;
srom_1(60406) <= 9555588;
srom_1(60407) <= 8984330;
srom_1(60408) <= 8410278;
srom_1(60409) <= 7836124;
srom_1(60410) <= 7264561;
srom_1(60411) <= 6698269;
srom_1(60412) <= 6139904;
srom_1(60413) <= 5592084;
srom_1(60414) <= 5057377;
srom_1(60415) <= 4538292;
srom_1(60416) <= 4037262;
srom_1(60417) <= 3556637;
srom_1(60418) <= 3098671;
srom_1(60419) <= 2665512;
srom_1(60420) <= 2259189;
srom_1(60421) <= 1881610;
srom_1(60422) <= 1534545;
srom_1(60423) <= 1219620;
srom_1(60424) <= 938313;
srom_1(60425) <= 691943;
srom_1(60426) <= 481666;
srom_1(60427) <= 308467;
srom_1(60428) <= 173158;
srom_1(60429) <= 76375;
srom_1(60430) <= 18570;
srom_1(60431) <= 15;
srom_1(60432) <= 20798;
srom_1(60433) <= 80820;
srom_1(60434) <= 179799;
srom_1(60435) <= 317273;
srom_1(60436) <= 492596;
srom_1(60437) <= 704947;
srom_1(60438) <= 953328;
srom_1(60439) <= 1236576;
srom_1(60440) <= 1553363;
srom_1(60441) <= 1902202;
srom_1(60442) <= 2281458;
srom_1(60443) <= 2689353;
srom_1(60444) <= 3123973;
srom_1(60445) <= 3583282;
srom_1(60446) <= 4065124;
srom_1(60447) <= 4567240;
srom_1(60448) <= 5087276;
srom_1(60449) <= 5622793;
srom_1(60450) <= 6171280;
srom_1(60451) <= 6730165;
srom_1(60452) <= 7296826;
srom_1(60453) <= 7868608;
srom_1(60454) <= 8442828;
srom_1(60455) <= 9016793;
srom_1(60456) <= 9587813;
srom_1(60457) <= 10153210;
srom_1(60458) <= 10710331;
srom_1(60459) <= 11256565;
srom_1(60460) <= 11789351;
srom_1(60461) <= 12306189;
srom_1(60462) <= 12804656;
srom_1(60463) <= 13282415;
srom_1(60464) <= 13737225;
srom_1(60465) <= 14166953;
srom_1(60466) <= 14569585;
srom_1(60467) <= 14943232;
srom_1(60468) <= 15286143;
srom_1(60469) <= 15596708;
srom_1(60470) <= 15873472;
srom_1(60471) <= 16115137;
srom_1(60472) <= 16320570;
srom_1(60473) <= 16488807;
srom_1(60474) <= 16619059;
srom_1(60475) <= 16710716;
srom_1(60476) <= 16763348;
srom_1(60477) <= 16776707;
srom_1(60478) <= 16750732;
srom_1(60479) <= 16685544;
srom_1(60480) <= 16581449;
srom_1(60481) <= 16438935;
srom_1(60482) <= 16258670;
srom_1(60483) <= 16041500;
srom_1(60484) <= 15788442;
srom_1(60485) <= 15500684;
srom_1(60486) <= 15179576;
srom_1(60487) <= 14826622;
srom_1(60488) <= 14443478;
srom_1(60489) <= 14031940;
srom_1(60490) <= 13593939;
srom_1(60491) <= 13131529;
srom_1(60492) <= 12646877;
srom_1(60493) <= 12142257;
srom_1(60494) <= 11620035;
srom_1(60495) <= 11082659;
srom_1(60496) <= 10532650;
srom_1(60497) <= 9972587;
srom_1(60498) <= 9405096;
srom_1(60499) <= 8832838;
srom_1(60500) <= 8258497;
srom_1(60501) <= 7684767;
srom_1(60502) <= 7114337;
srom_1(60503) <= 6549882;
srom_1(60504) <= 5994050;
srom_1(60505) <= 5449447;
srom_1(60506) <= 4918626;
srom_1(60507) <= 4404077;
srom_1(60508) <= 3908214;
srom_1(60509) <= 3433360;
srom_1(60510) <= 2981743;
srom_1(60511) <= 2555481;
srom_1(60512) <= 2156572;
srom_1(60513) <= 1786888;
srom_1(60514) <= 1448161;
srom_1(60515) <= 1141980;
srom_1(60516) <= 869781;
srom_1(60517) <= 632841;
srom_1(60518) <= 432270;
srom_1(60519) <= 269009;
srom_1(60520) <= 143824;
srom_1(60521) <= 57301;
srom_1(60522) <= 9846;
srom_1(60523) <= 1683;
srom_1(60524) <= 32849;
srom_1(60525) <= 103197;
srom_1(60526) <= 212399;
srom_1(60527) <= 359942;
srom_1(60528) <= 545134;
srom_1(60529) <= 767107;
srom_1(60530) <= 1024819;
srom_1(60531) <= 1317063;
srom_1(60532) <= 1642468;
srom_1(60533) <= 1999508;
srom_1(60534) <= 2386508;
srom_1(60535) <= 2801655;
srom_1(60536) <= 3243000;
srom_1(60537) <= 3708475;
srom_1(60538) <= 4195897;
srom_1(60539) <= 4702980;
srom_1(60540) <= 5227346;
srom_1(60541) <= 5766536;
srom_1(60542) <= 6318022;
srom_1(60543) <= 6879217;
srom_1(60544) <= 7447491;
srom_1(60545) <= 8020178;
srom_1(60546) <= 8594593;
srom_1(60547) <= 9168041;
srom_1(60548) <= 9737835;
srom_1(60549) <= 10301302;
srom_1(60550) <= 10855799;
srom_1(60551) <= 11398727;
srom_1(60552) <= 11927539;
srom_1(60553) <= 12439756;
srom_1(60554) <= 12932976;
srom_1(60555) <= 13404886;
srom_1(60556) <= 13853273;
srom_1(60557) <= 14276034;
srom_1(60558) <= 14671187;
srom_1(60559) <= 15036878;
srom_1(60560) <= 15371394;
srom_1(60561) <= 15673165;
srom_1(60562) <= 15940776;
srom_1(60563) <= 16172972;
srom_1(60564) <= 16368665;
srom_1(60565) <= 16526937;
srom_1(60566) <= 16647045;
srom_1(60567) <= 16728426;
srom_1(60568) <= 16770700;
srom_1(60569) <= 16773666;
srom_1(60570) <= 16737313;
srom_1(60571) <= 16661809;
srom_1(60572) <= 16547510;
srom_1(60573) <= 16394950;
srom_1(60574) <= 16204846;
srom_1(60575) <= 15978089;
srom_1(60576) <= 15715743;
srom_1(60577) <= 15419037;
srom_1(60578) <= 15089362;
srom_1(60579) <= 14728266;
srom_1(60580) <= 14337441;
srom_1(60581) <= 13918719;
srom_1(60582) <= 13474065;
srom_1(60583) <= 13005564;
srom_1(60584) <= 12515412;
srom_1(60585) <= 12005908;
srom_1(60586) <= 11479442;
srom_1(60587) <= 10938481;
srom_1(60588) <= 10385563;
srom_1(60589) <= 9823281;
srom_1(60590) <= 9254271;
srom_1(60591) <= 8681201;
srom_1(60592) <= 8106760;
srom_1(60593) <= 7533640;
srom_1(60594) <= 6964530;
srom_1(60595) <= 6402097;
srom_1(60596) <= 5848980;
srom_1(60597) <= 5307772;
srom_1(60598) <= 4781011;
srom_1(60599) <= 4271167;
srom_1(60600) <= 3780632;
srom_1(60601) <= 3311705;
srom_1(60602) <= 2866585;
srom_1(60603) <= 2447360;
srom_1(60604) <= 2055995;
srom_1(60605) <= 1694326;
srom_1(60606) <= 1364049;
srom_1(60607) <= 1066713;
srom_1(60608) <= 803711;
srom_1(60609) <= 576278;
srom_1(60610) <= 385479;
srom_1(60611) <= 232210;
srom_1(60612) <= 117188;
srom_1(60613) <= 40955;
srom_1(60614) <= 3866;
srom_1(60615) <= 6096;
srom_1(60616) <= 47635;
srom_1(60617) <= 128288;
srom_1(60618) <= 247676;
srom_1(60619) <= 405239;
srom_1(60620) <= 600239;
srom_1(60621) <= 831762;
srom_1(60622) <= 1098721;
srom_1(60623) <= 1399865;
srom_1(60624) <= 1733782;
srom_1(60625) <= 2098905;
srom_1(60626) <= 2493523;
srom_1(60627) <= 2915785;
srom_1(60628) <= 3363711;
srom_1(60629) <= 3835201;
srom_1(60630) <= 4328043;
srom_1(60631) <= 4839926;
srom_1(60632) <= 5368450;
srom_1(60633) <= 5911137;
srom_1(60634) <= 6465442;
srom_1(60635) <= 7028764;
srom_1(60636) <= 7598464;
srom_1(60637) <= 8171869;
srom_1(60638) <= 8746290;
srom_1(60639) <= 9319034;
srom_1(60640) <= 9887415;
srom_1(60641) <= 10448768;
srom_1(60642) <= 11000459;
srom_1(60643) <= 11539903;
srom_1(60644) <= 12064569;
srom_1(60645) <= 12571998;
srom_1(60646) <= 13059809;
srom_1(60647) <= 13525715;
srom_1(60648) <= 13967532;
srom_1(60649) <= 14383187;
srom_1(60650) <= 14770731;
srom_1(60651) <= 15128347;
srom_1(60652) <= 15454359;
srom_1(60653) <= 15747237;
srom_1(60654) <= 16005607;
srom_1(60655) <= 16228259;
srom_1(60656) <= 16414148;
srom_1(60657) <= 16562402;
srom_1(60658) <= 16672327;
srom_1(60659) <= 16743407;
srom_1(60660) <= 16775308;
srom_1(60661) <= 16767881;
srom_1(60662) <= 16721160;
srom_1(60663) <= 16635366;
srom_1(60664) <= 16510899;
srom_1(60665) <= 16348344;
srom_1(60666) <= 16148464;
srom_1(60667) <= 15912194;
srom_1(60668) <= 15640644;
srom_1(60669) <= 15335087;
srom_1(60670) <= 14996955;
srom_1(60671) <= 14627835;
srom_1(60672) <= 14229456;
srom_1(60673) <= 13803688;
srom_1(60674) <= 13352527;
srom_1(60675) <= 12878088;
srom_1(60676) <= 12382596;
srom_1(60677) <= 11868375;
srom_1(60678) <= 11337837;
srom_1(60679) <= 10793468;
srom_1(60680) <= 10237822;
srom_1(60681) <= 9673505;
srom_1(60682) <= 9103162;
srom_1(60683) <= 8529469;
srom_1(60684) <= 7955115;
srom_1(60685) <= 7382793;
srom_1(60686) <= 6815189;
srom_1(60687) <= 6254962;
srom_1(60688) <= 5704741;
srom_1(60689) <= 5167106;
srom_1(60690) <= 4644577;
srom_1(60691) <= 4139605;
srom_1(60692) <= 3654559;
srom_1(60693) <= 3191712;
srom_1(60694) <= 2753234;
srom_1(60695) <= 2341184;
srom_1(60696) <= 1957491;
srom_1(60697) <= 1603957;
srom_1(60698) <= 1282237;
srom_1(60699) <= 993842;
srom_1(60700) <= 740124;
srom_1(60701) <= 522272;
srom_1(60702) <= 341308;
srom_1(60703) <= 198081;
srom_1(60704) <= 93261;
srom_1(60705) <= 27342;
srom_1(60706) <= 631;
srom_1(60707) <= 13254;
srom_1(60708) <= 65153;
srom_1(60709) <= 156082;
srom_1(60710) <= 285617;
srom_1(60711) <= 453150;
srom_1(60712) <= 657895;
srom_1(60713) <= 898891;
srom_1(60714) <= 1175010;
srom_1(60715) <= 1484955;
srom_1(60716) <= 1827274;
srom_1(60717) <= 2200362;
srom_1(60718) <= 2602468;
srom_1(60719) <= 3031708;
srom_1(60720) <= 3486068;
srom_1(60721) <= 3963417;
srom_1(60722) <= 4461518;
srom_1(60723) <= 4978034;
srom_1(60724) <= 5510544;
srom_1(60725) <= 6056549;
srom_1(60726) <= 6613491;
srom_1(60727) <= 7178757;
srom_1(60728) <= 7749696;
srom_1(60729) <= 8323631;
srom_1(60730) <= 8897871;
srom_1(60731) <= 9469723;
srom_1(60732) <= 10036505;
srom_1(60733) <= 10595559;
srom_1(60734) <= 11144265;
srom_1(60735) <= 11680048;
srom_1(60736) <= 12200396;
srom_1(60737) <= 12702870;
srom_1(60738) <= 13185112;
srom_1(60739) <= 13644862;
srom_1(60740) <= 14079964;
srom_1(60741) <= 14488377;
srom_1(60742) <= 14868186;
srom_1(60743) <= 15217610;
srom_1(60744) <= 15535011;
srom_1(60745) <= 15818899;
srom_1(60746) <= 16067945;
srom_1(60747) <= 16280979;
srom_1(60748) <= 16457003;
srom_1(60749) <= 16595192;
srom_1(60750) <= 16694897;
srom_1(60751) <= 16755652;
srom_1(60752) <= 16777170;
srom_1(60753) <= 16759351;
srom_1(60754) <= 16702280;
srom_1(60755) <= 16606222;
srom_1(60756) <= 16471629;
srom_1(60757) <= 16299132;
srom_1(60758) <= 16089540;
srom_1(60759) <= 15843836;
srom_1(60760) <= 15563172;
srom_1(60761) <= 15248863;
srom_1(60762) <= 14902385;
srom_1(60763) <= 14525361;
srom_1(60764) <= 14119560;
srom_1(60765) <= 13686884;
srom_1(60766) <= 13229363;
srom_1(60767) <= 12749142;
srom_1(60768) <= 12248473;
srom_1(60769) <= 11729703;
srom_1(60770) <= 11195266;
srom_1(60771) <= 10647668;
srom_1(60772) <= 10089476;
srom_1(60773) <= 9523309;
srom_1(60774) <= 8951820;
srom_1(60775) <= 8377690;
srom_1(60776) <= 7803611;
srom_1(60777) <= 7232276;
srom_1(60778) <= 6666363;
srom_1(60779) <= 6108526;
srom_1(60780) <= 5561381;
srom_1(60781) <= 5027494;
srom_1(60782) <= 4509369;
srom_1(60783) <= 4009434;
srom_1(60784) <= 3530035;
srom_1(60785) <= 3073420;
srom_1(60786) <= 2641729;
srom_1(60787) <= 2236988;
srom_1(60788) <= 1861093;
srom_1(60789) <= 1515808;
srom_1(60790) <= 1202752;
srom_1(60791) <= 923393;
srom_1(60792) <= 679041;
srom_1(60793) <= 470842;
srom_1(60794) <= 299772;
srom_1(60795) <= 166633;
srom_1(60796) <= 72050;
srom_1(60797) <= 16466;
srom_1(60798) <= 142;
srom_1(60799) <= 23154;
srom_1(60800) <= 85395;
srom_1(60801) <= 186572;
srom_1(60802) <= 326212;
srom_1(60803) <= 503659;
srom_1(60804) <= 718081;
srom_1(60805) <= 968473;
srom_1(60806) <= 1253660;
srom_1(60807) <= 1572306;
srom_1(60808) <= 1922915;
srom_1(60809) <= 2303845;
srom_1(60810) <= 2713308;
srom_1(60811) <= 3149384;
srom_1(60812) <= 3610029;
srom_1(60813) <= 4093082;
srom_1(60814) <= 4596279;
srom_1(60815) <= 5117259;
srom_1(60816) <= 5653579;
srom_1(60817) <= 6202725;
srom_1(60818) <= 6762122;
srom_1(60819) <= 7329145;
srom_1(60820) <= 7901137;
srom_1(60821) <= 8475414;
srom_1(60822) <= 9049285;
srom_1(60823) <= 9620057;
srom_1(60824) <= 10185055;
srom_1(60825) <= 10741628;
srom_1(60826) <= 11287168;
srom_1(60827) <= 11819115;
srom_1(60828) <= 12334975;
srom_1(60829) <= 12832329;
srom_1(60830) <= 13308845;
srom_1(60831) <= 13762289;
srom_1(60832) <= 14190533;
srom_1(60833) <= 14591570;
srom_1(60834) <= 14963520;
srom_1(60835) <= 15304637;
srom_1(60836) <= 15613323;
srom_1(60837) <= 15888129;
srom_1(60838) <= 16127768;
srom_1(60839) <= 16331115;
srom_1(60840) <= 16497217;
srom_1(60841) <= 16625295;
srom_1(60842) <= 16714748;
srom_1(60843) <= 16765157;
srom_1(60844) <= 16776286;
srom_1(60845) <= 16748082;
srom_1(60846) <= 16680677;
srom_1(60847) <= 16574388;
srom_1(60848) <= 16429713;
srom_1(60849) <= 16247331;
srom_1(60850) <= 16028096;
srom_1(60851) <= 15773037;
srom_1(60852) <= 15483350;
srom_1(60853) <= 15160394;
srom_1(60854) <= 14805682;
srom_1(60855) <= 14420878;
srom_1(60856) <= 14007787;
srom_1(60857) <= 13568345;
srom_1(60858) <= 13104614;
srom_1(60859) <= 12618768;
srom_1(60860) <= 12113085;
srom_1(60861) <= 11589937;
srom_1(60862) <= 11051777;
srom_1(60863) <= 10501128;
srom_1(60864) <= 9940573;
srom_1(60865) <= 9372741;
srom_1(60866) <= 8800293;
srom_1(60867) <= 8225915;
srom_1(60868) <= 7652299;
srom_1(60869) <= 7082137;
srom_1(60870) <= 6518101;
srom_1(60871) <= 5962836;
srom_1(60872) <= 5418947;
srom_1(60873) <= 4888983;
srom_1(60874) <= 4375431;
srom_1(60875) <= 3880697;
srom_1(60876) <= 3407103;
srom_1(60877) <= 2956868;
srom_1(60878) <= 2532105;
srom_1(60879) <= 2134805;
srom_1(60880) <= 1766832;
srom_1(60881) <= 1429910;
srom_1(60882) <= 1125620;
srom_1(60883) <= 855388;
srom_1(60884) <= 620482;
srom_1(60885) <= 422004;
srom_1(60886) <= 260884;
srom_1(60887) <= 137877;
srom_1(60888) <= 53561;
srom_1(60889) <= 8331;
srom_1(60890) <= 2399;
srom_1(60891) <= 35793;
srom_1(60892) <= 108356;
srom_1(60893) <= 219748;
srom_1(60894) <= 369446;
srom_1(60895) <= 556749;
srom_1(60896) <= 780778;
srom_1(60897) <= 1040483;
srom_1(60898) <= 1334646;
srom_1(60899) <= 1661888;
srom_1(60900) <= 2020673;
srom_1(60901) <= 2409319;
srom_1(60902) <= 2826005;
srom_1(60903) <= 3268776;
srom_1(60904) <= 3735555;
srom_1(60905) <= 4224154;
srom_1(60906) <= 4732281;
srom_1(60907) <= 5257555;
srom_1(60908) <= 5797510;
srom_1(60909) <= 6349617;
srom_1(60910) <= 6911285;
srom_1(60911) <= 7479880;
srom_1(60912) <= 8052737;
srom_1(60913) <= 8627169;
srom_1(60914) <= 9200482;
srom_1(60915) <= 9769988;
srom_1(60916) <= 10333017;
srom_1(60917) <= 10886927;
srom_1(60918) <= 11429122;
srom_1(60919) <= 11957058;
srom_1(60920) <= 12468262;
srom_1(60921) <= 12960334;
srom_1(60922) <= 13430967;
srom_1(60923) <= 13877956;
srom_1(60924) <= 14299203;
srom_1(60925) <= 14692733;
srom_1(60926) <= 15056701;
srom_1(60927) <= 15389400;
srom_1(60928) <= 15689270;
srom_1(60929) <= 15954904;
srom_1(60930) <= 16185058;
srom_1(60931) <= 16378651;
srom_1(60932) <= 16534776;
srom_1(60933) <= 16652701;
srom_1(60934) <= 16731873;
srom_1(60935) <= 16771920;
srom_1(60936) <= 16772656;
srom_1(60937) <= 16734075;
srom_1(60938) <= 16656360;
srom_1(60939) <= 16539874;
srom_1(60940) <= 16385165;
srom_1(60941) <= 16192956;
srom_1(60942) <= 15964151;
srom_1(60943) <= 15699821;
srom_1(60944) <= 15401206;
srom_1(60945) <= 15069707;
srom_1(60946) <= 14706878;
srom_1(60947) <= 14314420;
srom_1(60948) <= 13894174;
srom_1(60949) <= 13448111;
srom_1(60950) <= 12978321;
srom_1(60951) <= 12487009;
srom_1(60952) <= 11976479;
srom_1(60953) <= 11449123;
srom_1(60954) <= 10907416;
srom_1(60955) <= 10353897;
srom_1(60956) <= 9791162;
srom_1(60957) <= 9221850;
srom_1(60958) <= 8648631;
srom_1(60959) <= 8074193;
srom_1(60960) <= 7501228;
srom_1(60961) <= 6932426;
srom_1(60962) <= 6370451;
srom_1(60963) <= 5817941;
srom_1(60964) <= 5277485;
srom_1(60965) <= 4751618;
srom_1(60966) <= 4242806;
srom_1(60967) <= 3753436;
srom_1(60968) <= 3285801;
srom_1(60969) <= 2842095;
srom_1(60970) <= 2424399;
srom_1(60971) <= 2034671;
srom_1(60972) <= 1674738;
srom_1(60973) <= 1346290;
srom_1(60974) <= 1050865;
srom_1(60975) <= 789849;
srom_1(60976) <= 564467;
srom_1(60977) <= 375774;
srom_1(60978) <= 224657;
srom_1(60979) <= 111823;
srom_1(60980) <= 37802;
srom_1(60981) <= 2940;
srom_1(60982) <= 7402;
srom_1(60983) <= 51166;
srom_1(60984) <= 134027;
srom_1(60985) <= 255597;
srom_1(60986) <= 415306;
srom_1(60987) <= 612403;
srom_1(60988) <= 845967;
srom_1(60989) <= 1114900;
srom_1(60990) <= 1417942;
srom_1(60991) <= 1753672;
srom_1(60992) <= 2120515;
srom_1(60993) <= 2516752;
srom_1(60994) <= 2940524;
srom_1(60995) <= 3389843;
srom_1(60996) <= 3862604;
srom_1(60997) <= 4356589;
srom_1(60998) <= 4869481;
srom_1(60999) <= 5398875;
srom_1(61000) <= 5942290;
srom_1(61001) <= 6497176;
srom_1(61002) <= 7060931;
srom_1(61003) <= 7630913;
srom_1(61004) <= 8204448;
srom_1(61005) <= 8778846;
srom_1(61006) <= 9351414;
srom_1(61007) <= 9919467;
srom_1(61008) <= 10480342;
srom_1(61009) <= 11031408;
srom_1(61010) <= 11570080;
srom_1(61011) <= 12093834;
srom_1(61012) <= 12600213;
srom_1(61013) <= 13086842;
srom_1(61014) <= 13551439;
srom_1(61015) <= 13991826;
srom_1(61016) <= 14405937;
srom_1(61017) <= 14791832;
srom_1(61018) <= 15147699;
srom_1(61019) <= 15471871;
srom_1(61020) <= 15762826;
srom_1(61021) <= 16019202;
srom_1(61022) <= 16239795;
srom_1(61023) <= 16423571;
srom_1(61024) <= 16569668;
srom_1(61025) <= 16677402;
srom_1(61026) <= 16746266;
srom_1(61027) <= 16775939;
srom_1(61028) <= 16766281;
srom_1(61029) <= 16717336;
srom_1(61030) <= 16629336;
srom_1(61031) <= 16502692;
srom_1(61032) <= 16337998;
srom_1(61033) <= 16136027;
srom_1(61034) <= 15897725;
srom_1(61035) <= 15624210;
srom_1(61036) <= 15316766;
srom_1(61037) <= 14976833;
srom_1(61038) <= 14606005;
srom_1(61039) <= 14206022;
srom_1(61040) <= 13778759;
srom_1(61041) <= 13326219;
srom_1(61042) <= 12850526;
srom_1(61043) <= 12353909;
srom_1(61044) <= 11838697;
srom_1(61045) <= 11307307;
srom_1(61046) <= 10762230;
srom_1(61047) <= 10206022;
srom_1(61048) <= 9641292;
srom_1(61049) <= 9070688;
srom_1(61050) <= 8496884;
srom_1(61051) <= 7922574;
srom_1(61052) <= 7350448;
srom_1(61053) <= 6783191;
srom_1(61054) <= 6223462;
srom_1(61055) <= 5673887;
srom_1(61056) <= 5137041;
srom_1(61057) <= 4615443;
srom_1(61058) <= 4111539;
srom_1(61059) <= 3627692;
srom_1(61060) <= 3166170;
srom_1(61061) <= 2729138;
srom_1(61062) <= 2318645;
srom_1(61063) <= 1936616;
srom_1(61064) <= 1584843;
srom_1(61065) <= 1264975;
srom_1(61066) <= 978512;
srom_1(61067) <= 726798;
srom_1(61068) <= 511012;
srom_1(61069) <= 332168;
srom_1(61070) <= 191102;
srom_1(61071) <= 88478;
srom_1(61072) <= 24776;
srom_1(61073) <= 294;
srom_1(61074) <= 15149;
srom_1(61075) <= 69269;
srom_1(61076) <= 162402;
srom_1(61077) <= 294110;
srom_1(61078) <= 463775;
srom_1(61079) <= 670604;
srom_1(61080) <= 913624;
srom_1(61081) <= 1191698;
srom_1(61082) <= 1503520;
srom_1(61083) <= 1847628;
srom_1(61084) <= 2222410;
srom_1(61085) <= 2626107;
srom_1(61086) <= 3056826;
srom_1(61087) <= 3512548;
srom_1(61088) <= 3991135;
srom_1(61089) <= 4490344;
srom_1(61090) <= 5007833;
srom_1(61091) <= 5541175;
srom_1(61092) <= 6087870;
srom_1(61093) <= 6645354;
srom_1(61094) <= 7211013;
srom_1(61095) <= 7782194;
srom_1(61096) <= 8356218;
srom_1(61097) <= 8930395;
srom_1(61098) <= 9502031;
srom_1(61099) <= 10068445;
srom_1(61100) <= 10626982;
srom_1(61101) <= 11175023;
srom_1(61102) <= 11709997;
srom_1(61103) <= 12229396;
srom_1(61104) <= 12730785;
srom_1(61105) <= 13211811;
srom_1(61106) <= 13670220;
srom_1(61107) <= 14103861;
srom_1(61108) <= 14510702;
srom_1(61109) <= 14888834;
srom_1(61110) <= 15236484;
srom_1(61111) <= 15552022;
srom_1(61112) <= 15833969;
srom_1(61113) <= 16081001;
srom_1(61114) <= 16291961;
srom_1(61115) <= 16465860;
srom_1(61116) <= 16601882;
srom_1(61117) <= 16699389;
srom_1(61118) <= 16757924;
srom_1(61119) <= 16777212;
srom_1(61120) <= 16757163;
srom_1(61121) <= 16697871;
srom_1(61122) <= 16599614;
srom_1(61123) <= 16462853;
srom_1(61124) <= 16288229;
srom_1(61125) <= 16076560;
srom_1(61126) <= 15828841;
srom_1(61127) <= 15546231;
srom_1(61128) <= 15230057;
srom_1(61129) <= 14881802;
srom_1(61130) <= 14503097;
srom_1(61131) <= 14095719;
srom_1(61132) <= 13661579;
srom_1(61133) <= 13202712;
srom_1(61134) <= 12721270;
srom_1(61135) <= 12219510;
srom_1(61136) <= 11699787;
srom_1(61137) <= 11164536;
srom_1(61138) <= 10616267;
srom_1(61139) <= 10057553;
srom_1(61140) <= 9491012;
srom_1(61141) <= 8919301;
srom_1(61142) <= 8345102;
srom_1(61143) <= 7771107;
srom_1(61144) <= 7200008;
srom_1(61145) <= 6634482;
srom_1(61146) <= 6077182;
srom_1(61147) <= 5530721;
srom_1(61148) <= 4997662;
srom_1(61149) <= 4480504;
srom_1(61150) <= 3981673;
srom_1(61151) <= 3503507;
srom_1(61152) <= 3048249;
srom_1(61153) <= 2618033;
srom_1(61154) <= 2214878;
srom_1(61155) <= 1840674;
srom_1(61156) <= 1497175;
srom_1(61157) <= 1185993;
srom_1(61158) <= 908586;
srom_1(61159) <= 666255;
srom_1(61160) <= 460137;
srom_1(61161) <= 291199;
srom_1(61162) <= 160232;
srom_1(61163) <= 67851;
srom_1(61164) <= 14488;
srom_1(61165) <= 395;
srom_1(61166) <= 25637;
srom_1(61167) <= 90096;
srom_1(61168) <= 193469;
srom_1(61169) <= 335272;
srom_1(61170) <= 514840;
srom_1(61171) <= 731331;
srom_1(61172) <= 983729;
srom_1(61173) <= 1270851;
srom_1(61174) <= 1591351;
srom_1(61175) <= 1943726;
srom_1(61176) <= 2326323;
srom_1(61177) <= 2737348;
srom_1(61178) <= 3174874;
srom_1(61179) <= 3636848;
srom_1(61180) <= 4121106;
srom_1(61181) <= 4625375;
srom_1(61182) <= 5147291;
srom_1(61183) <= 5684407;
srom_1(61184) <= 6234204;
srom_1(61185) <= 6794103;
srom_1(61186) <= 7361480;
srom_1(61187) <= 7933673;
srom_1(61188) <= 8508000;
srom_1(61189) <= 9081766;
srom_1(61190) <= 9652283;
srom_1(61191) <= 10216873;
srom_1(61192) <= 10772890;
srom_1(61193) <= 11317726;
srom_1(61194) <= 11848827;
srom_1(61195) <= 12363701;
srom_1(61196) <= 12859935;
srom_1(61197) <= 13335202;
srom_1(61198) <= 13787272;
srom_1(61199) <= 14214026;
srom_1(61200) <= 14613462;
srom_1(61201) <= 14983708;
srom_1(61202) <= 15323027;
srom_1(61203) <= 15629829;
srom_1(61204) <= 15902673;
srom_1(61205) <= 16140282;
srom_1(61206) <= 16341541;
srom_1(61207) <= 16505505;
srom_1(61208) <= 16631407;
srom_1(61209) <= 16718655;
srom_1(61210) <= 16766841;
srom_1(61211) <= 16775738;
srom_1(61212) <= 16745305;
srom_1(61213) <= 16675685;
srom_1(61214) <= 16567204;
srom_1(61215) <= 16420370;
srom_1(61216) <= 16235873;
srom_1(61217) <= 16014577;
srom_1(61218) <= 15757521;
srom_1(61219) <= 15465909;
srom_1(61220) <= 15141109;
srom_1(61221) <= 14784645;
srom_1(61222) <= 14398187;
srom_1(61223) <= 13983548;
srom_1(61224) <= 13542673;
srom_1(61225) <= 13077628;
srom_1(61226) <= 12590595;
srom_1(61227) <= 12083858;
srom_1(61228) <= 11559792;
srom_1(61229) <= 11020855;
srom_1(61230) <= 10469575;
srom_1(61231) <= 9908536;
srom_1(61232) <= 9340370;
srom_1(61233) <= 8767741;
srom_1(61234) <= 8193334;
srom_1(61235) <= 7619843;
srom_1(61236) <= 7049957;
srom_1(61237) <= 6486348;
srom_1(61238) <= 5931659;
srom_1(61239) <= 5388492;
srom_1(61240) <= 4859393;
srom_1(61241) <= 4346844;
srom_1(61242) <= 3853249;
srom_1(61243) <= 3380921;
srom_1(61244) <= 2932076;
srom_1(61245) <= 2508818;
srom_1(61246) <= 2113133;
srom_1(61247) <= 1746876;
srom_1(61248) <= 1411764;
srom_1(61249) <= 1109369;
srom_1(61250) <= 841108;
srom_1(61251) <= 608241;
srom_1(61252) <= 411858;
srom_1(61253) <= 252881;
srom_1(61254) <= 132055;
srom_1(61255) <= 49947;
srom_1(61256) <= 6942;
srom_1(61257) <= 3242;
srom_1(61258) <= 38863;
srom_1(61259) <= 113639;
srom_1(61260) <= 227219;
srom_1(61261) <= 379071;
srom_1(61262) <= 568482;
srom_1(61263) <= 794565;
srom_1(61264) <= 1056258;
srom_1(61265) <= 1352336;
srom_1(61266) <= 1681409;
srom_1(61267) <= 2041934;
srom_1(61268) <= 2432221;
srom_1(61269) <= 2850440;
srom_1(61270) <= 3294629;
srom_1(61271) <= 3762705;
srom_1(61272) <= 4252474;
srom_1(61273) <= 4761638;
srom_1(61274) <= 5287811;
srom_1(61275) <= 5828524;
srom_1(61276) <= 6381243;
srom_1(61277) <= 6943374;
srom_1(61278) <= 7512283;
srom_1(61279) <= 8085301;
srom_1(61280) <= 8659742;
srom_1(61281) <= 9232911;
srom_1(61282) <= 9802121;
srom_1(61283) <= 10364702;
srom_1(61284) <= 10918017;
srom_1(61285) <= 11459471;
srom_1(61286) <= 11986524;
srom_1(61287) <= 12496705;
srom_1(61288) <= 12987622;
srom_1(61289) <= 13456973;
srom_1(61290) <= 13902556;
srom_1(61291) <= 14322283;
srom_1(61292) <= 14714184;
srom_1(61293) <= 15076423;
srom_1(61294) <= 15407300;
srom_1(61295) <= 15705264;
srom_1(61296) <= 15968918;
srom_1(61297) <= 16197025;
srom_1(61298) <= 16388516;
srom_1(61299) <= 16542493;
srom_1(61300) <= 16658233;
srom_1(61301) <= 16735194;
srom_1(61302) <= 16773015;
srom_1(61303) <= 16771518;
srom_1(61304) <= 16730712;
srom_1(61305) <= 16650786;
srom_1(61306) <= 16532116;
srom_1(61307) <= 16375258;
srom_1(61308) <= 16180948;
srom_1(61309) <= 15950098;
srom_1(61310) <= 15683788;
srom_1(61311) <= 15383270;
srom_1(61312) <= 15049950;
srom_1(61313) <= 14685394;
srom_1(61314) <= 14291309;
srom_1(61315) <= 13869545;
srom_1(61316) <= 13422079;
srom_1(61317) <= 12951009;
srom_1(61318) <= 12458545;
srom_1(61319) <= 11946995;
srom_1(61320) <= 11418759;
srom_1(61321) <= 10876313;
srom_1(61322) <= 10322201;
srom_1(61323) <= 9759023;
srom_1(61324) <= 9189418;
srom_1(61325) <= 8616057;
srom_1(61326) <= 8041630;
srom_1(61327) <= 7468830;
srom_1(61328) <= 6900344;
srom_1(61329) <= 6338836;
srom_1(61330) <= 5786940;
srom_1(61331) <= 5247244;
srom_1(61332) <= 4722280;
srom_1(61333) <= 4214508;
srom_1(61334) <= 3726310;
srom_1(61335) <= 3259974;
srom_1(61336) <= 2817689;
srom_1(61337) <= 2401528;
srom_1(61338) <= 2013442;
srom_1(61339) <= 1655252;
srom_1(61340) <= 1328636;
srom_1(61341) <= 1035128;
srom_1(61342) <= 776102;
srom_1(61343) <= 552774;
srom_1(61344) <= 366190;
srom_1(61345) <= 217227;
srom_1(61346) <= 106582;
srom_1(61347) <= 34774;
srom_1(61348) <= 2141;
srom_1(61349) <= 8834;
srom_1(61350) <= 54823;
srom_1(61351) <= 139892;
srom_1(61352) <= 263642;
srom_1(61353) <= 425492;
srom_1(61354) <= 624685;
srom_1(61355) <= 860285;
srom_1(61356) <= 1131188;
srom_1(61357) <= 1436124;
srom_1(61358) <= 1773662;
srom_1(61359) <= 2142220;
srom_1(61360) <= 2540069;
srom_1(61361) <= 2965344;
srom_1(61362) <= 3416051;
srom_1(61363) <= 3890076;
srom_1(61364) <= 4385196;
srom_1(61365) <= 4899089;
srom_1(61366) <= 5429346;
srom_1(61367) <= 5973480;
srom_1(61368) <= 6528939;
srom_1(61369) <= 7093118;
srom_1(61370) <= 7663373;
srom_1(61371) <= 8237029;
srom_1(61372) <= 8811395;
srom_1(61373) <= 9383779;
srom_1(61374) <= 9951496;
srom_1(61375) <= 10511885;
srom_1(61376) <= 11062316;
srom_1(61377) <= 11600209;
srom_1(61378) <= 12123043;
srom_1(61379) <= 12628364;
srom_1(61380) <= 13113803;
srom_1(61381) <= 13577085;
srom_1(61382) <= 14016035;
srom_1(61383) <= 14428597;
srom_1(61384) <= 14812835;
srom_1(61385) <= 15166948;
srom_1(61386) <= 15489275;
srom_1(61387) <= 15778305;
srom_1(61388) <= 16032681;
srom_1(61389) <= 16251212;
srom_1(61390) <= 16432872;
srom_1(61391) <= 16576811;
srom_1(61392) <= 16682351;
srom_1(61393) <= 16749000;
srom_1(61394) <= 16776444;
srom_1(61395) <= 16764554;
srom_1(61396) <= 16713387;
srom_1(61397) <= 16623182;
srom_1(61398) <= 16494362;
srom_1(61399) <= 16327531;
srom_1(61400) <= 16123473;
srom_1(61401) <= 15883142;
srom_1(61402) <= 15607667;
srom_1(61403) <= 15298340;
srom_1(61404) <= 14956611;
srom_1(61405) <= 14584081;
srom_1(61406) <= 14182500;
srom_1(61407) <= 13753748;
srom_1(61408) <= 13299838;
srom_1(61409) <= 12822897;
srom_1(61410) <= 12325162;
srom_1(61411) <= 11808967;
srom_1(61412) <= 11276734;
srom_1(61413) <= 10730956;
srom_1(61414) <= 10174195;
srom_1(61415) <= 9609060;
srom_1(61416) <= 9038203;
srom_1(61417) <= 8464299;
srom_1(61418) <= 7890040;
srom_1(61419) <= 7318119;
srom_1(61420) <= 6751218;
srom_1(61421) <= 6191995;
srom_1(61422) <= 5643073;
srom_1(61423) <= 5107026;
srom_1(61424) <= 4586367;
srom_1(61425) <= 4083538;
srom_1(61426) <= 3600897;
srom_1(61427) <= 3140707;
srom_1(61428) <= 2705127;
srom_1(61429) <= 2296198;
srom_1(61430) <= 1915839;
srom_1(61431) <= 1565832;
srom_1(61432) <= 1247820;
srom_1(61433) <= 963294;
srom_1(61434) <= 713588;
srom_1(61435) <= 499872;
srom_1(61436) <= 323149;
srom_1(61437) <= 184248;
srom_1(61438) <= 83820;
srom_1(61439) <= 22336;
srom_1(61440) <= 84;
srom_1(61441) <= 17169;
srom_1(61442) <= 73511;
srom_1(61443) <= 168845;
srom_1(61444) <= 302724;
srom_1(61445) <= 474521;
srom_1(61446) <= 683429;
srom_1(61447) <= 928470;
srom_1(61448) <= 1208494;
srom_1(61449) <= 1522188;
srom_1(61450) <= 1868081;
srom_1(61451) <= 2244551;
srom_1(61452) <= 2649832;
srom_1(61453) <= 3082025;
srom_1(61454) <= 3539102;
srom_1(61455) <= 4018919;
srom_1(61456) <= 4519228;
srom_1(61457) <= 5037682;
srom_1(61458) <= 5571849;
srom_1(61459) <= 6119226;
srom_1(61460) <= 6677244;
srom_1(61461) <= 7243287;
srom_1(61462) <= 7814701;
srom_1(61463) <= 8388806;
srom_1(61464) <= 8962910;
srom_1(61465) <= 9534322;
srom_1(61466) <= 10100360;
srom_1(61467) <= 10658372;
srom_1(61468) <= 11205740;
srom_1(61469) <= 11739897;
srom_1(61470) <= 12258339;
srom_1(61471) <= 12758634;
srom_1(61472) <= 13238437;
srom_1(61473) <= 13695498;
srom_1(61474) <= 14127672;
srom_1(61475) <= 14532934;
srom_1(61476) <= 14909383;
srom_1(61477) <= 15255255;
srom_1(61478) <= 15568926;
srom_1(61479) <= 15848926;
srom_1(61480) <= 16093942;
srom_1(61481) <= 16302825;
srom_1(61482) <= 16474595;
srom_1(61483) <= 16608448;
srom_1(61484) <= 16703755;
srom_1(61485) <= 16760069;
srom_1(61486) <= 16777127;
srom_1(61487) <= 16754848;
srom_1(61488) <= 16693337;
srom_1(61489) <= 16592882;
srom_1(61490) <= 16453954;
srom_1(61491) <= 16277205;
srom_1(61492) <= 16063464;
srom_1(61493) <= 15813733;
srom_1(61494) <= 15529183;
srom_1(61495) <= 15211148;
srom_1(61496) <= 14861120;
srom_1(61497) <= 14480741;
srom_1(61498) <= 14071793;
srom_1(61499) <= 13636194;
srom_1(61500) <= 13175988;
srom_1(61501) <= 12693333;
srom_1(61502) <= 12190490;
srom_1(61503) <= 11669820;
srom_1(61504) <= 11133763;
srom_1(61505) <= 10584833;
srom_1(61506) <= 10025604;
srom_1(61507) <= 9458698;
srom_1(61508) <= 8886775;
srom_1(61509) <= 8312515;
srom_1(61510) <= 7738612;
srom_1(61511) <= 7167758;
srom_1(61512) <= 6602628;
srom_1(61513) <= 6045873;
srom_1(61514) <= 5500105;
srom_1(61515) <= 4967881;
srom_1(61516) <= 4451698;
srom_1(61517) <= 3953977;
srom_1(61518) <= 3477052;
srom_1(61519) <= 3023158;
srom_1(61520) <= 2594425;
srom_1(61521) <= 2192862;
srom_1(61522) <= 1820354;
srom_1(61523) <= 1478647;
srom_1(61524) <= 1169342;
srom_1(61525) <= 893891;
srom_1(61526) <= 653586;
srom_1(61527) <= 449553;
srom_1(61528) <= 282748;
srom_1(61529) <= 153955;
srom_1(61530) <= 63777;
srom_1(61531) <= 12637;
srom_1(61532) <= 775;
srom_1(61533) <= 28246;
srom_1(61534) <= 94921;
srom_1(61535) <= 200489;
srom_1(61536) <= 344454;
srom_1(61537) <= 526140;
srom_1(61538) <= 744696;
srom_1(61539) <= 999097;
srom_1(61540) <= 1288150;
srom_1(61541) <= 1610500;
srom_1(61542) <= 1964634;
srom_1(61543) <= 2348893;
srom_1(61544) <= 2761474;
srom_1(61545) <= 3200442;
srom_1(61546) <= 3663740;
srom_1(61547) <= 4149194;
srom_1(61548) <= 4654528;
srom_1(61549) <= 5177372;
srom_1(61550) <= 5715275;
srom_1(61551) <= 6265715;
srom_1(61552) <= 6826109;
srom_1(61553) <= 7393830;
srom_1(61554) <= 7966216;
srom_1(61555) <= 8540583;
srom_1(61556) <= 9114237;
srom_1(61557) <= 9684489;
srom_1(61558) <= 10248664;
srom_1(61559) <= 10804116;
srom_1(61560) <= 11348241;
srom_1(61561) <= 11878487;
srom_1(61562) <= 12392368;
srom_1(61563) <= 12887474;
srom_1(61564) <= 13361483;
srom_1(61565) <= 13812173;
srom_1(61566) <= 14237430;
srom_1(61567) <= 14635260;
srom_1(61568) <= 15003797;
srom_1(61569) <= 15341313;
srom_1(61570) <= 15646225;
srom_1(61571) <= 15917104;
srom_1(61572) <= 16152679;
srom_1(61573) <= 16351846;
srom_1(61574) <= 16513671;
srom_1(61575) <= 16637394;
srom_1(61576) <= 16722436;
srom_1(61577) <= 16768397;
srom_1(61578) <= 16775063;
srom_1(61579) <= 16742402;
srom_1(61580) <= 16670568;
srom_1(61581) <= 16559896;
srom_1(61582) <= 16410906;
srom_1(61583) <= 16224297;
srom_1(61584) <= 16000944;
srom_1(61585) <= 15741893;
srom_1(61586) <= 15448361;
srom_1(61587) <= 15121723;
srom_1(61588) <= 14763511;
srom_1(61589) <= 14375405;
srom_1(61590) <= 13959225;
srom_1(61591) <= 13516923;
srom_1(61592) <= 13050572;
srom_1(61593) <= 12562359;
srom_1(61594) <= 12054574;
srom_1(61595) <= 11529598;
srom_1(61596) <= 10989893;
srom_1(61597) <= 10437990;
srom_1(61598) <= 9876477;
srom_1(61599) <= 9307986;
srom_1(61600) <= 8735184;
srom_1(61601) <= 8160757;
srom_1(61602) <= 7587398;
srom_1(61603) <= 7017796;
srom_1(61604) <= 6454623;
srom_1(61605) <= 5900519;
srom_1(61606) <= 5358082;
srom_1(61607) <= 4829856;
srom_1(61608) <= 4318319;
srom_1(61609) <= 3825869;
srom_1(61610) <= 3354814;
srom_1(61611) <= 2907365;
srom_1(61612) <= 2485620;
srom_1(61613) <= 2091555;
srom_1(61614) <= 1727020;
srom_1(61615) <= 1393723;
srom_1(61616) <= 1093228;
srom_1(61617) <= 826943;
srom_1(61618) <= 596117;
srom_1(61619) <= 401833;
srom_1(61620) <= 245001;
srom_1(61621) <= 126358;
srom_1(61622) <= 46460;
srom_1(61623) <= 5680;
srom_1(61624) <= 4211;
srom_1(61625) <= 42059;
srom_1(61626) <= 119047;
srom_1(61627) <= 234814;
srom_1(61628) <= 388817;
srom_1(61629) <= 580334;
srom_1(61630) <= 808466;
srom_1(61631) <= 1072144;
srom_1(61632) <= 1370131;
srom_1(61633) <= 1701031;
srom_1(61634) <= 2063291;
srom_1(61635) <= 2455212;
srom_1(61636) <= 2874958;
srom_1(61637) <= 3320558;
srom_1(61638) <= 3789925;
srom_1(61639) <= 4280856;
srom_1(61640) <= 4791050;
srom_1(61641) <= 5318114;
srom_1(61642) <= 5859577;
srom_1(61643) <= 6412899;
srom_1(61644) <= 6975486;
srom_1(61645) <= 7544699;
srom_1(61646) <= 8117870;
srom_1(61647) <= 8692311;
srom_1(61648) <= 9265327;
srom_1(61649) <= 9834232;
srom_1(61650) <= 10396358;
srom_1(61651) <= 10949069;
srom_1(61652) <= 11489773;
srom_1(61653) <= 12015935;
srom_1(61654) <= 12525087;
srom_1(61655) <= 13014841;
srom_1(61656) <= 13482902;
srom_1(61657) <= 13927073;
srom_1(61658) <= 14345273;
srom_1(61659) <= 14735540;
srom_1(61660) <= 15096044;
srom_1(61661) <= 15425095;
srom_1(61662) <= 15721149;
srom_1(61663) <= 15982818;
srom_1(61664) <= 16208875;
srom_1(61665) <= 16398261;
srom_1(61666) <= 16550086;
srom_1(61667) <= 16663639;
srom_1(61668) <= 16738388;
srom_1(61669) <= 16773982;
srom_1(61670) <= 16770254;
srom_1(61671) <= 16727222;
srom_1(61672) <= 16645087;
srom_1(61673) <= 16524235;
srom_1(61674) <= 16365231;
srom_1(61675) <= 16168823;
srom_1(61676) <= 15935930;
srom_1(61677) <= 15667646;
srom_1(61678) <= 15365228;
srom_1(61679) <= 15030093;
srom_1(61680) <= 14663815;
srom_1(61681) <= 14268110;
srom_1(61682) <= 13844834;
srom_1(61683) <= 13395972;
srom_1(61684) <= 12923629;
srom_1(61685) <= 12430019;
srom_1(61686) <= 11917458;
srom_1(61687) <= 11388348;
srom_1(61688) <= 10845172;
srom_1(61689) <= 10290477;
srom_1(61690) <= 9726862;
srom_1(61691) <= 9156973;
srom_1(61692) <= 8583480;
srom_1(61693) <= 8009073;
srom_1(61694) <= 7436446;
srom_1(61695) <= 6868284;
srom_1(61696) <= 6307251;
srom_1(61697) <= 5755979;
srom_1(61698) <= 5217052;
srom_1(61699) <= 4692997;
srom_1(61700) <= 4186272;
srom_1(61701) <= 3699254;
srom_1(61702) <= 3234225;
srom_1(61703) <= 2793367;
srom_1(61704) <= 2378748;
srom_1(61705) <= 1992310;
srom_1(61706) <= 1635867;
srom_1(61707) <= 1311090;
srom_1(61708) <= 1019501;
srom_1(61709) <= 762469;
srom_1(61710) <= 541199;
srom_1(61711) <= 356728;
srom_1(61712) <= 209921;
srom_1(61713) <= 101466;
srom_1(61714) <= 31873;
srom_1(61715) <= 1468;
srom_1(61716) <= 10392;
srom_1(61717) <= 58605;
srom_1(61718) <= 145880;
srom_1(61719) <= 271809;
srom_1(61720) <= 435799;
srom_1(61721) <= 637083;
srom_1(61722) <= 874717;
srom_1(61723) <= 1147586;
srom_1(61724) <= 1454410;
srom_1(61725) <= 1793752;
srom_1(61726) <= 2164019;
srom_1(61727) <= 2563475;
srom_1(61728) <= 2990247;
srom_1(61729) <= 3442334;
srom_1(61730) <= 3917615;
srom_1(61731) <= 4413863;
srom_1(61732) <= 4928750;
srom_1(61733) <= 5459861;
srom_1(61734) <= 6004706;
srom_1(61735) <= 6560730;
srom_1(61736) <= 7125325;
srom_1(61737) <= 7695844;
srom_1(61738) <= 8269612;
srom_1(61739) <= 8843938;
srom_1(61740) <= 9416129;
srom_1(61741) <= 9983502;
srom_1(61742) <= 10543395;
srom_1(61743) <= 11093184;
srom_1(61744) <= 11630290;
srom_1(61745) <= 12152195;
srom_1(61746) <= 12656451;
srom_1(61747) <= 13140693;
srom_1(61748) <= 13602652;
srom_1(61749) <= 14040160;
srom_1(61750) <= 14451166;
srom_1(61751) <= 14833742;
srom_1(61752) <= 15186095;
srom_1(61753) <= 15506573;
srom_1(61754) <= 15793671;
srom_1(61755) <= 16046045;
srom_1(61756) <= 16262511;
srom_1(61757) <= 16442053;
srom_1(61758) <= 16583829;
srom_1(61759) <= 16687176;
srom_1(61760) <= 16751607;
srom_1(61761) <= 16776822;
srom_1(61762) <= 16762701;
srom_1(61763) <= 16709312;
srom_1(61764) <= 16616903;
srom_1(61765) <= 16485910;
srom_1(61766) <= 16316945;
srom_1(61767) <= 16110802;
srom_1(61768) <= 15868446;
srom_1(61769) <= 15591016;
srom_1(61770) <= 15279810;
srom_1(61771) <= 14936289;
srom_1(61772) <= 14562064;
srom_1(61773) <= 14158890;
srom_1(61774) <= 13728656;
srom_1(61775) <= 13273382;
srom_1(61776) <= 12795201;
srom_1(61777) <= 12296356;
srom_1(61778) <= 11779186;
srom_1(61779) <= 11246116;
srom_1(61780) <= 10699647;
srom_1(61781) <= 10142340;
srom_1(61782) <= 9576810;
srom_1(61783) <= 9005708;
srom_1(61784) <= 8431712;
srom_1(61785) <= 7857513;
srom_1(61786) <= 7285806;
srom_1(61787) <= 6719269;
srom_1(61788) <= 6160561;
srom_1(61789) <= 5612301;
srom_1(61790) <= 5077060;
srom_1(61791) <= 4557347;
srom_1(61792) <= 4055601;
srom_1(61793) <= 3574174;
srom_1(61794) <= 3115324;
srom_1(61795) <= 2681201;
srom_1(61796) <= 2273843;
srom_1(61797) <= 1895159;
srom_1(61798) <= 1546925;
srom_1(61799) <= 1230773;
srom_1(61800) <= 948188;
srom_1(61801) <= 700493;
srom_1(61802) <= 488850;
srom_1(61803) <= 314252;
srom_1(61804) <= 177517;
srom_1(61805) <= 79287;
srom_1(61806) <= 20023;
srom_1(61807) <= 1;
srom_1(61808) <= 19317;
srom_1(61809) <= 77878;
srom_1(61810) <= 175412;
srom_1(61811) <= 311461;
srom_1(61812) <= 485385;
srom_1(61813) <= 696371;
srom_1(61814) <= 943428;
srom_1(61815) <= 1225399;
srom_1(61816) <= 1540960;
srom_1(61817) <= 1888631;
srom_1(61818) <= 2266784;
srom_1(61819) <= 2673644;
srom_1(61820) <= 3107303;
srom_1(61821) <= 3565728;
srom_1(61822) <= 4046770;
srom_1(61823) <= 4548171;
srom_1(61824) <= 5067582;
srom_1(61825) <= 5602566;
srom_1(61826) <= 6150615;
srom_1(61827) <= 6709159;
srom_1(61828) <= 7275578;
srom_1(61829) <= 7847217;
srom_1(61830) <= 8421394;
srom_1(61831) <= 8995417;
srom_1(61832) <= 9566595;
srom_1(61833) <= 10132249;
srom_1(61834) <= 10689727;
srom_1(61835) <= 11236413;
srom_1(61836) <= 11769746;
srom_1(61837) <= 12287223;
srom_1(61838) <= 12786418;
srom_1(61839) <= 13264990;
srom_1(61840) <= 13720695;
srom_1(61841) <= 14151396;
srom_1(61842) <= 14555074;
srom_1(61843) <= 14929835;
srom_1(61844) <= 15273921;
srom_1(61845) <= 15585721;
srom_1(61846) <= 15863770;
srom_1(61847) <= 16106766;
srom_1(61848) <= 16313568;
srom_1(61849) <= 16483208;
srom_1(61850) <= 16614890;
srom_1(61851) <= 16707995;
srom_1(61852) <= 16762088;
srom_1(61853) <= 16776915;
srom_1(61854) <= 16752407;
srom_1(61855) <= 16688677;
srom_1(61856) <= 16586026;
srom_1(61857) <= 16444934;
srom_1(61858) <= 16266063;
srom_1(61859) <= 16050252;
srom_1(61860) <= 15798514;
srom_1(61861) <= 15512027;
srom_1(61862) <= 15192136;
srom_1(61863) <= 14840342;
srom_1(61864) <= 14458292;
srom_1(61865) <= 14047780;
srom_1(61866) <= 13610731;
srom_1(61867) <= 13149192;
srom_1(61868) <= 12665330;
srom_1(61869) <= 12161413;
srom_1(61870) <= 11639804;
srom_1(61871) <= 11102949;
srom_1(61872) <= 10553365;
srom_1(61873) <= 9993630;
srom_1(61874) <= 9426369;
srom_1(61875) <= 8854241;
srom_1(61876) <= 8279929;
srom_1(61877) <= 7706128;
srom_1(61878) <= 7135526;
srom_1(61879) <= 6570801;
srom_1(61880) <= 6014600;
srom_1(61881) <= 5469532;
srom_1(61882) <= 4938152;
srom_1(61883) <= 4422952;
srom_1(61884) <= 3926349;
srom_1(61885) <= 3450671;
srom_1(61886) <= 2998148;
srom_1(61887) <= 2570904;
srom_1(61888) <= 2170940;
srom_1(61889) <= 1800133;
srom_1(61890) <= 1460222;
srom_1(61891) <= 1152801;
srom_1(61892) <= 879310;
srom_1(61893) <= 641033;
srom_1(61894) <= 439088;
srom_1(61895) <= 274420;
srom_1(61896) <= 147803;
srom_1(61897) <= 59829;
srom_1(61898) <= 10912;
srom_1(61899) <= 1281;
srom_1(61900) <= 30981;
srom_1(61901) <= 99873;
srom_1(61902) <= 207633;
srom_1(61903) <= 353757;
srom_1(61904) <= 537559;
srom_1(61905) <= 758177;
srom_1(61906) <= 1014577;
srom_1(61907) <= 1305556;
srom_1(61908) <= 1629751;
srom_1(61909) <= 1985639;
srom_1(61910) <= 2371554;
srom_1(61911) <= 2785684;
srom_1(61912) <= 3226089;
srom_1(61913) <= 3690702;
srom_1(61914) <= 4177346;
srom_1(61915) <= 4683737;
srom_1(61916) <= 5207502;
srom_1(61917) <= 5746184;
srom_1(61918) <= 6297258;
srom_1(61919) <= 6858138;
srom_1(61920) <= 7426195;
srom_1(61921) <= 7998766;
srom_1(61922) <= 8573164;
srom_1(61923) <= 9146698;
srom_1(61924) <= 9716676;
srom_1(61925) <= 10280426;
srom_1(61926) <= 10835305;
srom_1(61927) <= 11378711;
srom_1(61928) <= 11908094;
srom_1(61929) <= 12420974;
srom_1(61930) <= 12914945;
srom_1(61931) <= 13387690;
srom_1(61932) <= 13836993;
srom_1(61933) <= 14260746;
srom_1(61934) <= 14656963;
srom_1(61935) <= 15023785;
srom_1(61936) <= 15359493;
srom_1(61937) <= 15662512;
srom_1(61938) <= 15931421;
srom_1(61939) <= 16164959;
srom_1(61940) <= 16362032;
srom_1(61941) <= 16521714;
srom_1(61942) <= 16643257;
srom_1(61943) <= 16726091;
srom_1(61944) <= 16769828;
srom_1(61945) <= 16774262;
srom_1(61946) <= 16739374;
srom_1(61947) <= 16665325;
srom_1(61948) <= 16552465;
srom_1(61949) <= 16401321;
srom_1(61950) <= 16212602;
srom_1(61951) <= 15987195;
srom_1(61952) <= 15726155;
srom_1(61953) <= 15430706;
srom_1(61954) <= 15102235;
srom_1(61955) <= 14742282;
srom_1(61956) <= 14352533;
srom_1(61957) <= 13934818;
srom_1(61958) <= 13491095;
srom_1(61959) <= 13023445;
srom_1(61960) <= 12534060;
srom_1(61961) <= 12025235;
srom_1(61962) <= 11499358;
srom_1(61963) <= 10958893;
srom_1(61964) <= 10406374;
srom_1(61965) <= 9844394;
srom_1(61966) <= 9275588;
srom_1(61967) <= 8702621;
srom_1(61968) <= 8128183;
srom_1(61969) <= 7554965;
srom_1(61970) <= 6985657;
srom_1(61971) <= 6422928;
srom_1(61972) <= 5869416;
srom_1(61973) <= 5327718;
srom_1(61974) <= 4800373;
srom_1(61975) <= 4289855;
srom_1(61976) <= 3798558;
srom_1(61977) <= 3328784;
srom_1(61978) <= 2882738;
srom_1(61979) <= 2462511;
srom_1(61980) <= 2070073;
srom_1(61981) <= 1707265;
srom_1(61982) <= 1375788;
srom_1(61983) <= 1077197;
srom_1(61984) <= 812891;
srom_1(61985) <= 584110;
srom_1(61986) <= 391928;
srom_1(61987) <= 237244;
srom_1(61988) <= 120786;
srom_1(61989) <= 43097;
srom_1(61990) <= 4544;
srom_1(61991) <= 5307;
srom_1(61992) <= 45381;
srom_1(61993) <= 124580;
srom_1(61994) <= 242532;
srom_1(61995) <= 398684;
srom_1(61996) <= 592303;
srom_1(61997) <= 822481;
srom_1(61998) <= 1088140;
srom_1(61999) <= 1388033;
srom_1(62000) <= 1720754;
srom_1(62001) <= 2084743;
srom_1(62002) <= 2478293;
srom_1(62003) <= 2899559;
srom_1(62004) <= 3346565;
srom_1(62005) <= 3817214;
srom_1(62006) <= 4309300;
srom_1(62007) <= 4820516;
srom_1(62008) <= 5348463;
srom_1(62009) <= 5890667;
srom_1(62010) <= 6444585;
srom_1(62011) <= 7007618;
srom_1(62012) <= 7577128;
srom_1(62013) <= 8150443;
srom_1(62014) <= 8724875;
srom_1(62015) <= 9297730;
srom_1(62016) <= 9866321;
srom_1(62017) <= 10427983;
srom_1(62018) <= 10980082;
srom_1(62019) <= 11520029;
srom_1(62020) <= 12045291;
srom_1(62021) <= 12553406;
srom_1(62022) <= 13041990;
srom_1(62023) <= 13508754;
srom_1(62024) <= 13951507;
srom_1(62025) <= 14368173;
srom_1(62026) <= 14756800;
srom_1(62027) <= 15115564;
srom_1(62028) <= 15442783;
srom_1(62029) <= 15736922;
srom_1(62030) <= 15996603;
srom_1(62031) <= 16220607;
srom_1(62032) <= 16407884;
srom_1(62033) <= 16557556;
srom_1(62034) <= 16668921;
srom_1(62035) <= 16741457;
srom_1(62036) <= 16774823;
srom_1(62037) <= 16768864;
srom_1(62038) <= 16723607;
srom_1(62039) <= 16639264;
srom_1(62040) <= 16516230;
srom_1(62041) <= 16355084;
srom_1(62042) <= 16156580;
srom_1(62043) <= 15921649;
srom_1(62044) <= 15651394;
srom_1(62045) <= 15347080;
srom_1(62046) <= 15010136;
srom_1(62047) <= 14642142;
srom_1(62048) <= 14244822;
srom_1(62049) <= 13820040;
srom_1(62050) <= 13369789;
srom_1(62051) <= 12896179;
srom_1(62052) <= 12401432;
srom_1(62053) <= 11887867;
srom_1(62054) <= 11357893;
srom_1(62055) <= 10813995;
srom_1(62056) <= 10258723;
srom_1(62057) <= 9694682;
srom_1(62058) <= 9124516;
srom_1(62059) <= 8550899;
srom_1(62060) <= 7976521;
srom_1(62061) <= 7404076;
srom_1(62062) <= 6836247;
srom_1(62063) <= 6275698;
srom_1(62064) <= 5725057;
srom_1(62065) <= 5186907;
srom_1(62066) <= 4663770;
srom_1(62067) <= 4158100;
srom_1(62068) <= 3672269;
srom_1(62069) <= 3208554;
srom_1(62070) <= 2769130;
srom_1(62071) <= 2356058;
srom_1(62072) <= 1971274;
srom_1(62073) <= 1616584;
srom_1(62074) <= 1293650;
srom_1(62075) <= 1003986;
srom_1(62076) <= 748952;
srom_1(62077) <= 529743;
srom_1(62078) <= 347386;
srom_1(62079) <= 202738;
srom_1(62080) <= 96476;
srom_1(62081) <= 29098;
srom_1(62082) <= 921;
srom_1(62083) <= 12077;
srom_1(62084) <= 62513;
srom_1(62085) <= 151994;
srom_1(62086) <= 280098;
srom_1(62087) <= 446226;
srom_1(62088) <= 649599;
srom_1(62089) <= 889263;
srom_1(62090) <= 1164093;
srom_1(62091) <= 1472802;
srom_1(62092) <= 1813941;
srom_1(62093) <= 2185911;
srom_1(62094) <= 2586968;
srom_1(62095) <= 3015231;
srom_1(62096) <= 3468691;
srom_1(62097) <= 3945222;
srom_1(62098) <= 4442590;
srom_1(62099) <= 4958463;
srom_1(62100) <= 5490420;
srom_1(62101) <= 6035968;
srom_1(62102) <= 6592548;
srom_1(62103) <= 7157551;
srom_1(62104) <= 7728326;
srom_1(62105) <= 8302198;
srom_1(62106) <= 8876475;
srom_1(62107) <= 9448464;
srom_1(62108) <= 10015483;
srom_1(62109) <= 10574873;
srom_1(62110) <= 11124011;
srom_1(62111) <= 11660322;
srom_1(62112) <= 12181290;
srom_1(62113) <= 12684474;
srom_1(62114) <= 13167512;
srom_1(62115) <= 13628141;
srom_1(62116) <= 14064199;
srom_1(62117) <= 14473643;
srom_1(62118) <= 14854552;
srom_1(62119) <= 15205140;
srom_1(62120) <= 15523763;
srom_1(62121) <= 15808927;
srom_1(62122) <= 16059294;
srom_1(62123) <= 16273691;
srom_1(62124) <= 16451111;
srom_1(62125) <= 16590724;
srom_1(62126) <= 16691875;
srom_1(62127) <= 16754089;
srom_1(62128) <= 16777074;
srom_1(62129) <= 16760722;
srom_1(62130) <= 16705111;
srom_1(62131) <= 16610501;
srom_1(62132) <= 16477335;
srom_1(62133) <= 16306239;
srom_1(62134) <= 16098015;
srom_1(62135) <= 15853638;
srom_1(62136) <= 15574255;
srom_1(62137) <= 15261176;
srom_1(62138) <= 14915869;
srom_1(62139) <= 14539954;
srom_1(62140) <= 14135193;
srom_1(62141) <= 13703484;
srom_1(62142) <= 13246852;
srom_1(62143) <= 12767438;
srom_1(62144) <= 12267490;
srom_1(62145) <= 11749353;
srom_1(62146) <= 11215456;
srom_1(62147) <= 10668303;
srom_1(62148) <= 10110460;
srom_1(62149) <= 9544542;
srom_1(62150) <= 8973204;
srom_1(62151) <= 8399124;
srom_1(62152) <= 7824995;
srom_1(62153) <= 7253509;
srom_1(62154) <= 6687346;
srom_1(62155) <= 6129160;
srom_1(62156) <= 5581570;
srom_1(62157) <= 5047144;
srom_1(62158) <= 4528386;
srom_1(62159) <= 4027730;
srom_1(62160) <= 3547524;
srom_1(62161) <= 3090020;
srom_1(62162) <= 2657362;
srom_1(62163) <= 2251580;
srom_1(62164) <= 1874577;
srom_1(62165) <= 1528120;
srom_1(62166) <= 1213834;
srom_1(62167) <= 933194;
srom_1(62168) <= 687514;
srom_1(62169) <= 477948;
srom_1(62170) <= 305477;
srom_1(62171) <= 170911;
srom_1(62172) <= 74880;
srom_1(62173) <= 17836;
srom_1(62174) <= 44;
srom_1(62175) <= 21590;
srom_1(62176) <= 82371;
srom_1(62177) <= 182104;
srom_1(62178) <= 320319;
srom_1(62179) <= 496369;
srom_1(62180) <= 709429;
srom_1(62181) <= 958499;
srom_1(62182) <= 1242411;
srom_1(62183) <= 1559835;
srom_1(62184) <= 1909280;
srom_1(62185) <= 2289110;
srom_1(62186) <= 2697542;
srom_1(62187) <= 3132662;
srom_1(62188) <= 3592428;
srom_1(62189) <= 4074686;
srom_1(62190) <= 4577172;
srom_1(62191) <= 5097532;
srom_1(62192) <= 5633325;
srom_1(62193) <= 6182039;
srom_1(62194) <= 6741100;
srom_1(62195) <= 7307886;
srom_1(62196) <= 7879740;
srom_1(62197) <= 8453981;
srom_1(62198) <= 9027915;
srom_1(62199) <= 9598851;
srom_1(62200) <= 10164112;
srom_1(62201) <= 10721047;
srom_1(62202) <= 11267044;
srom_1(62203) <= 11799544;
srom_1(62204) <= 12316048;
srom_1(62205) <= 12814135;
srom_1(62206) <= 13291469;
srom_1(62207) <= 13745812;
srom_1(62208) <= 14175034;
srom_1(62209) <= 14577121;
srom_1(62210) <= 14950187;
srom_1(62211) <= 15292484;
srom_1(62212) <= 15602407;
srom_1(62213) <= 15878502;
srom_1(62214) <= 16119473;
srom_1(62215) <= 16324193;
srom_1(62216) <= 16491699;
srom_1(62217) <= 16621207;
srom_1(62218) <= 16712110;
srom_1(62219) <= 16763981;
srom_1(62220) <= 16776577;
srom_1(62221) <= 16749839;
srom_1(62222) <= 16683892;
srom_1(62223) <= 16579046;
srom_1(62224) <= 16435792;
srom_1(62225) <= 16254802;
srom_1(62226) <= 16036925;
srom_1(62227) <= 15783182;
srom_1(62228) <= 15494764;
srom_1(62229) <= 15173022;
srom_1(62230) <= 14819465;
srom_1(62231) <= 14435753;
srom_1(62232) <= 14023683;
srom_1(62233) <= 13585188;
srom_1(62234) <= 13122325;
srom_1(62235) <= 12637264;
srom_1(62236) <= 12132279;
srom_1(62237) <= 11609739;
srom_1(62238) <= 11072094;
srom_1(62239) <= 10521865;
srom_1(62240) <= 9961632;
srom_1(62241) <= 9394023;
srom_1(62242) <= 8821700;
srom_1(62243) <= 8247345;
srom_1(62244) <= 7673653;
srom_1(62245) <= 7103314;
srom_1(62246) <= 6539001;
srom_1(62247) <= 5983362;
srom_1(62248) <= 5439003;
srom_1(62249) <= 4908474;
srom_1(62250) <= 4394266;
srom_1(62251) <= 3898788;
srom_1(62252) <= 3424364;
srom_1(62253) <= 2973220;
srom_1(62254) <= 2547470;
srom_1(62255) <= 2149111;
srom_1(62256) <= 1780012;
srom_1(62257) <= 1441902;
srom_1(62258) <= 1136368;
srom_1(62259) <= 864842;
srom_1(62260) <= 628598;
srom_1(62261) <= 428743;
srom_1(62262) <= 266214;
srom_1(62263) <= 141774;
srom_1(62264) <= 56007;
srom_1(62265) <= 9314;
srom_1(62266) <= 1914;
srom_1(62267) <= 33842;
srom_1(62268) <= 104949;
srom_1(62269) <= 214900;
srom_1(62270) <= 363181;
srom_1(62271) <= 549096;
srom_1(62272) <= 771773;
srom_1(62273) <= 1030168;
srom_1(62274) <= 1323069;
srom_1(62275) <= 1649103;
srom_1(62276) <= 2006741;
srom_1(62277) <= 2394306;
srom_1(62278) <= 2809979;
srom_1(62279) <= 3251813;
srom_1(62280) <= 3717736;
srom_1(62281) <= 4205561;
srom_1(62282) <= 4713002;
srom_1(62283) <= 5237680;
srom_1(62284) <= 5777133;
srom_1(62285) <= 6328832;
srom_1(62286) <= 6890190;
srom_1(62287) <= 7458575;
srom_1(62288) <= 8031321;
srom_1(62289) <= 8605743;
srom_1(62290) <= 9179146;
srom_1(62291) <= 9748842;
srom_1(62292) <= 10312160;
srom_1(62293) <= 10866457;
srom_1(62294) <= 11409135;
srom_1(62295) <= 11937649;
srom_1(62296) <= 12449520;
srom_1(62297) <= 12942348;
srom_1(62298) <= 13413821;
srom_1(62299) <= 13861730;
srom_1(62300) <= 14283974;
srom_1(62301) <= 14678572;
srom_1(62302) <= 15043674;
srom_1(62303) <= 15377569;
srom_1(62304) <= 15678689;
srom_1(62305) <= 15945624;
srom_1(62306) <= 16177122;
srom_1(62307) <= 16372097;
srom_1(62308) <= 16529634;
srom_1(62309) <= 16648995;
srom_1(62310) <= 16729620;
srom_1(62311) <= 16771132;
srom_1(62312) <= 16773335;
srom_1(62313) <= 16736219;
srom_1(62314) <= 16659958;
srom_1(62315) <= 16544910;
srom_1(62316) <= 16391614;
srom_1(62317) <= 16200790;
srom_1(62318) <= 15973331;
srom_1(62319) <= 15710306;
srom_1(62320) <= 15412946;
srom_1(62321) <= 15082646;
srom_1(62322) <= 14720956;
srom_1(62323) <= 14329572;
srom_1(62324) <= 13910328;
srom_1(62325) <= 13465191;
srom_1(62326) <= 12996248;
srom_1(62327) <= 12505698;
srom_1(62328) <= 11995842;
srom_1(62329) <= 11469070;
srom_1(62330) <= 10927853;
srom_1(62331) <= 10374728;
srom_1(62332) <= 9812290;
srom_1(62333) <= 9243176;
srom_1(62334) <= 8670054;
srom_1(62335) <= 8095613;
srom_1(62336) <= 7522545;
srom_1(62337) <= 6953539;
srom_1(62338) <= 6391262;
srom_1(62339) <= 5838352;
srom_1(62340) <= 5297400;
srom_1(62341) <= 4770945;
srom_1(62342) <= 4261453;
srom_1(62343) <= 3771316;
srom_1(62344) <= 3302830;
srom_1(62345) <= 2858193;
srom_1(62346) <= 2439491;
srom_1(62347) <= 2048686;
srom_1(62348) <= 1687611;
srom_1(62349) <= 1357959;
srom_1(62350) <= 1061276;
srom_1(62351) <= 798954;
srom_1(62352) <= 572222;
srom_1(62353) <= 382144;
srom_1(62354) <= 229611;
srom_1(62355) <= 115338;
srom_1(62356) <= 39861;
srom_1(62357) <= 3535;
srom_1(62358) <= 6529;
srom_1(62359) <= 48830;
srom_1(62360) <= 130238;
srom_1(62361) <= 250373;
srom_1(62362) <= 408671;
srom_1(62363) <= 604389;
srom_1(62364) <= 836611;
srom_1(62365) <= 1104246;
srom_1(62366) <= 1406040;
srom_1(62367) <= 1740578;
srom_1(62368) <= 2106291;
srom_1(62369) <= 2501464;
srom_1(62370) <= 2924243;
srom_1(62371) <= 3372647;
srom_1(62372) <= 3844572;
srom_1(62373) <= 4337806;
srom_1(62374) <= 4850036;
srom_1(62375) <= 5378859;
srom_1(62376) <= 5921795;
srom_1(62377) <= 6476300;
srom_1(62378) <= 7039772;
srom_1(62379) <= 7609569;
srom_1(62380) <= 8183019;
srom_1(62381) <= 8757434;
srom_1(62382) <= 9330118;
srom_1(62383) <= 9898388;
srom_1(62384) <= 10459578;
srom_1(62385) <= 11011056;
srom_1(62386) <= 11550237;
srom_1(62387) <= 12074592;
srom_1(62388) <= 12581662;
srom_1(62389) <= 13069069;
srom_1(62390) <= 13534528;
srom_1(62391) <= 13975856;
srom_1(62392) <= 14390984;
srom_1(62393) <= 14777964;
srom_1(62394) <= 15134982;
srom_1(62395) <= 15460365;
srom_1(62396) <= 15752585;
srom_1(62397) <= 16010273;
srom_1(62398) <= 16232221;
srom_1(62399) <= 16417387;
srom_1(62400) <= 16564903;
srom_1(62401) <= 16674078;
srom_1(62402) <= 16744400;
srom_1(62403) <= 16775538;
srom_1(62404) <= 16767347;
srom_1(62405) <= 16719866;
srom_1(62406) <= 16633316;
srom_1(62407) <= 16508104;
srom_1(62408) <= 16344817;
srom_1(62409) <= 16144220;
srom_1(62410) <= 15907255;
srom_1(62411) <= 15635032;
srom_1(62412) <= 15328828;
srom_1(62413) <= 14990079;
srom_1(62414) <= 14620374;
srom_1(62415) <= 14221445;
srom_1(62416) <= 13795165;
srom_1(62417) <= 13343531;
srom_1(62418) <= 12868662;
srom_1(62419) <= 12372784;
srom_1(62420) <= 11858224;
srom_1(62421) <= 11327393;
srom_1(62422) <= 10782781;
srom_1(62423) <= 10226941;
srom_1(62424) <= 9662482;
srom_1(62425) <= 9092048;
srom_1(62426) <= 8518316;
srom_1(62427) <= 7943976;
srom_1(62428) <= 7371721;
srom_1(62429) <= 6804234;
srom_1(62430) <= 6244177;
srom_1(62431) <= 5694176;
srom_1(62432) <= 5156810;
srom_1(62433) <= 4634599;
srom_1(62434) <= 4129992;
srom_1(62435) <= 3645355;
srom_1(62436) <= 3182961;
srom_1(62437) <= 2744977;
srom_1(62438) <= 2333459;
srom_1(62439) <= 1950335;
srom_1(62440) <= 1597403;
srom_1(62441) <= 1276317;
srom_1(62442) <= 988583;
srom_1(62443) <= 735550;
srom_1(62444) <= 518405;
srom_1(62445) <= 338166;
srom_1(62446) <= 195678;
srom_1(62447) <= 91610;
srom_1(62448) <= 26449;
srom_1(62449) <= 501;
srom_1(62450) <= 13888;
srom_1(62451) <= 66547;
srom_1(62452) <= 158231;
srom_1(62453) <= 288510;
srom_1(62454) <= 456773;
srom_1(62455) <= 662231;
srom_1(62456) <= 903921;
srom_1(62457) <= 1180709;
srom_1(62458) <= 1491298;
srom_1(62459) <= 1834230;
srom_1(62460) <= 2207898;
srom_1(62461) <= 2610549;
srom_1(62462) <= 3040296;
srom_1(62463) <= 3495123;
srom_1(62464) <= 3972897;
srom_1(62465) <= 4471377;
srom_1(62466) <= 4988227;
srom_1(62467) <= 5521023;
srom_1(62468) <= 6067266;
srom_1(62469) <= 6624394;
srom_1(62470) <= 7189795;
srom_1(62471) <= 7760818;
srom_1(62472) <= 8334785;
srom_1(62473) <= 8909004;
srom_1(62474) <= 9480782;
srom_1(62475) <= 10047440;
srom_1(62476) <= 10606318;
srom_1(62477) <= 11154797;
srom_1(62478) <= 11690304;
srom_1(62479) <= 12210328;
srom_1(62480) <= 12712431;
srom_1(62481) <= 13194259;
srom_1(62482) <= 13653550;
srom_1(62483) <= 14088153;
srom_1(62484) <= 14496028;
srom_1(62485) <= 14875264;
srom_1(62486) <= 15224082;
srom_1(62487) <= 15540845;
srom_1(62488) <= 15824070;
srom_1(62489) <= 16072427;
srom_1(62490) <= 16284751;
srom_1(62491) <= 16460048;
srom_1(62492) <= 16597496;
srom_1(62493) <= 16696449;
srom_1(62494) <= 16756443;
srom_1(62495) <= 16777198;
srom_1(62496) <= 16758617;
srom_1(62497) <= 16700785;
srom_1(62498) <= 16603974;
srom_1(62499) <= 16468639;
srom_1(62500) <= 16295414;
srom_1(62501) <= 16085111;
srom_1(62502) <= 15838716;
srom_1(62503) <= 15557386;
srom_1(62504) <= 15242438;
srom_1(62505) <= 14895351;
srom_1(62506) <= 14517751;
srom_1(62507) <= 14111410;
srom_1(62508) <= 13678232;
srom_1(62509) <= 13220249;
srom_1(62510) <= 12739610;
srom_1(62511) <= 12238566;
srom_1(62512) <= 11719469;
srom_1(62513) <= 11184753;
srom_1(62514) <= 10636924;
srom_1(62515) <= 10078553;
srom_1(62516) <= 9512256;
srom_1(62517) <= 8940691;
srom_1(62518) <= 8366536;
srom_1(62519) <= 7792485;
srom_1(62520) <= 7221230;
srom_1(62521) <= 6655448;
srom_1(62522) <= 6097794;
srom_1(62523) <= 5550883;
srom_1(62524) <= 5017278;
srom_1(62525) <= 4499483;
srom_1(62526) <= 3999925;
srom_1(62527) <= 3520947;
srom_1(62528) <= 3064796;
srom_1(62529) <= 2633609;
srom_1(62530) <= 2229410;
srom_1(62531) <= 1854093;
srom_1(62532) <= 1509419;
srom_1(62533) <= 1197004;
srom_1(62534) <= 918312;
srom_1(62535) <= 674652;
srom_1(62536) <= 467165;
srom_1(62537) <= 296824;
srom_1(62538) <= 164428;
srom_1(62539) <= 70598;
srom_1(62540) <= 15775;
srom_1(62541) <= 214;
srom_1(62542) <= 23990;
srom_1(62543) <= 86990;
srom_1(62544) <= 188919;
srom_1(62545) <= 329299;
srom_1(62546) <= 507472;
srom_1(62547) <= 722603;
srom_1(62548) <= 973682;
srom_1(62549) <= 1259532;
srom_1(62550) <= 1578813;
srom_1(62551) <= 1930027;
srom_1(62552) <= 2311528;
srom_1(62553) <= 2721526;
srom_1(62554) <= 3158099;
srom_1(62555) <= 3619200;
srom_1(62556) <= 4102667;
srom_1(62557) <= 4606231;
srom_1(62558) <= 5127532;
srom_1(62559) <= 5664126;
srom_1(62560) <= 6213496;
srom_1(62561) <= 6773065;
srom_1(62562) <= 7340210;
srom_1(62563) <= 7912272;
srom_1(62564) <= 8486567;
srom_1(62565) <= 9060403;
srom_1(62566) <= 9631089;
srom_1(62567) <= 10195948;
srom_1(62568) <= 10752332;
srom_1(62569) <= 11297632;
srom_1(62570) <= 11829290;
srom_1(62571) <= 12344814;
srom_1(62572) <= 12841785;
srom_1(62573) <= 13317875;
srom_1(62574) <= 13770849;
srom_1(62575) <= 14198584;
srom_1(62576) <= 14599074;
srom_1(62577) <= 14970441;
srom_1(62578) <= 15310943;
srom_1(62579) <= 15618984;
srom_1(62580) <= 15893120;
srom_1(62581) <= 16132064;
srom_1(62582) <= 16334697;
srom_1(62583) <= 16500068;
srom_1(62584) <= 16627401;
srom_1(62585) <= 16716099;
srom_1(62586) <= 16765748;
srom_1(62587) <= 16776113;
srom_1(62588) <= 16747146;
srom_1(62589) <= 16678982;
srom_1(62590) <= 16571943;
srom_1(62591) <= 16426529;
srom_1(62592) <= 16243423;
srom_1(62593) <= 16023482;
srom_1(62594) <= 15767739;
srom_1(62595) <= 15477393;
srom_1(62596) <= 15153805;
srom_1(62597) <= 14798492;
srom_1(62598) <= 14413122;
srom_1(62599) <= 13999500;
srom_1(62600) <= 13559567;
srom_1(62601) <= 13095386;
srom_1(62602) <= 12609133;
srom_1(62603) <= 12103088;
srom_1(62604) <= 11579625;
srom_1(62605) <= 11041198;
srom_1(62606) <= 10490332;
srom_1(62607) <= 9929611;
srom_1(62608) <= 9361663;
srom_1(62609) <= 8789152;
srom_1(62610) <= 8214763;
srom_1(62611) <= 7641189;
srom_1(62612) <= 7071120;
srom_1(62613) <= 6507229;
srom_1(62614) <= 5952161;
srom_1(62615) <= 5408518;
srom_1(62616) <= 4878850;
srom_1(62617) <= 4365640;
srom_1(62618) <= 3871295;
srom_1(62619) <= 3398133;
srom_1(62620) <= 2948373;
srom_1(62621) <= 2524125;
srom_1(62622) <= 2127377;
srom_1(62623) <= 1759990;
srom_1(62624) <= 1423687;
srom_1(62625) <= 1120045;
srom_1(62626) <= 850488;
srom_1(62627) <= 616279;
srom_1(62628) <= 418518;
srom_1(62629) <= 258131;
srom_1(62630) <= 135871;
srom_1(62631) <= 52310;
srom_1(62632) <= 7842;
srom_1(62633) <= 2673;
srom_1(62634) <= 36829;
srom_1(62635) <= 110150;
srom_1(62636) <= 222291;
srom_1(62637) <= 372727;
srom_1(62638) <= 560752;
srom_1(62639) <= 785484;
srom_1(62640) <= 1045870;
srom_1(62641) <= 1340689;
srom_1(62642) <= 1668558;
srom_1(62643) <= 2027939;
srom_1(62644) <= 2417148;
srom_1(62645) <= 2834359;
srom_1(62646) <= 3277616;
srom_1(62647) <= 3744840;
srom_1(62648) <= 4233840;
srom_1(62649) <= 4742323;
srom_1(62650) <= 5267905;
srom_1(62651) <= 5808121;
srom_1(62652) <= 6360438;
srom_1(62653) <= 6922265;
srom_1(62654) <= 7490969;
srom_1(62655) <= 8063882;
srom_1(62656) <= 8638318;
srom_1(62657) <= 9211583;
srom_1(62658) <= 9780989;
srom_1(62659) <= 10343865;
srom_1(62660) <= 10897572;
srom_1(62661) <= 11439514;
srom_1(62662) <= 11967150;
srom_1(62663) <= 12478004;
srom_1(62664) <= 12969681;
srom_1(62665) <= 13439877;
srom_1(62666) <= 13886385;
srom_1(62667) <= 14307112;
srom_1(62668) <= 14700086;
srom_1(62669) <= 15063462;
srom_1(62670) <= 15395538;
srom_1(62671) <= 15694756;
srom_1(62672) <= 15959714;
srom_1(62673) <= 16189167;
srom_1(62674) <= 16382041;
srom_1(62675) <= 16537431;
srom_1(62676) <= 16654608;
srom_1(62677) <= 16733024;
srom_1(62678) <= 16772309;
srom_1(62679) <= 16772281;
srom_1(62680) <= 16732938;
srom_1(62681) <= 16654466;
srom_1(62682) <= 16537233;
srom_1(62683) <= 16381787;
srom_1(62684) <= 16188860;
srom_1(62685) <= 15959354;
srom_1(62686) <= 15694346;
srom_1(62687) <= 15395079;
srom_1(62688) <= 15062956;
srom_1(62689) <= 14699535;
srom_1(62690) <= 14306520;
srom_1(62691) <= 13885754;
srom_1(62692) <= 13439209;
srom_1(62693) <= 12968981;
srom_1(62694) <= 12477274;
srom_1(62695) <= 11966394;
srom_1(62696) <= 11438736;
srom_1(62697) <= 10896775;
srom_1(62698) <= 10343052;
srom_1(62699) <= 9780164;
srom_1(62700) <= 9210751;
srom_1(62701) <= 8637483;
srom_1(62702) <= 8063047;
srom_1(62703) <= 7490138;
srom_1(62704) <= 6921442;
srom_1(62705) <= 6359627;
srom_1(62706) <= 5807326;
srom_1(62707) <= 5267129;
srom_1(62708) <= 4741570;
srom_1(62709) <= 4233114;
srom_1(62710) <= 3744143;
srom_1(62711) <= 3276953;
srom_1(62712) <= 2833732;
srom_1(62713) <= 2416561;
srom_1(62714) <= 2027394;
srom_1(62715) <= 1668057;
srom_1(62716) <= 1340236;
srom_1(62717) <= 1045466;
srom_1(62718) <= 785131;
srom_1(62719) <= 560451;
srom_1(62720) <= 372480;
srom_1(62721) <= 222100;
srom_1(62722) <= 110015;
srom_1(62723) <= 36751;
srom_1(62724) <= 2652;
srom_1(62725) <= 7878;
srom_1(62726) <= 52403;
srom_1(62727) <= 136020;
srom_1(62728) <= 258337;
srom_1(62729) <= 418779;
srom_1(62730) <= 616594;
srom_1(62731) <= 850854;
srom_1(62732) <= 1120462;
srom_1(62733) <= 1424153;
srom_1(62734) <= 1760502;
srom_1(62735) <= 2127933;
srom_1(62736) <= 2524723;
srom_1(62737) <= 2949010;
srom_1(62738) <= 3398805;
srom_1(62739) <= 3871999;
srom_1(62740) <= 4366373;
srom_1(62741) <= 4879609;
srom_1(62742) <= 5409299;
srom_1(62743) <= 5952961;
srom_1(62744) <= 6508044;
srom_1(62745) <= 7071946;
srom_1(62746) <= 7642022;
srom_1(62747) <= 8215599;
srom_1(62748) <= 8789987;
srom_1(62749) <= 9362493;
srom_1(62750) <= 9930432;
srom_1(62751) <= 10491141;
srom_1(62752) <= 11041991;
srom_1(62753) <= 11580398;
srom_1(62754) <= 12103837;
srom_1(62755) <= 12609855;
srom_1(62756) <= 13096078;
srom_1(62757) <= 13560225;
srom_1(62758) <= 14000121;
srom_1(62759) <= 14413703;
srom_1(62760) <= 14799031;
srom_1(62761) <= 15154299;
srom_1(62762) <= 15477840;
srom_1(62763) <= 15768137;
srom_1(62764) <= 16023828;
srom_1(62765) <= 16243716;
srom_1(62766) <= 16426768;
srom_1(62767) <= 16572127;
srom_1(62768) <= 16679110;
srom_1(62769) <= 16747216;
srom_1(62770) <= 16776126;
srom_1(62771) <= 16765704;
srom_1(62772) <= 16715999;
srom_1(62773) <= 16627243;
srom_1(62774) <= 16499854;
srom_1(62775) <= 16334429;
srom_1(62776) <= 16131743;
srom_1(62777) <= 15892747;
srom_1(62778) <= 15618561;
srom_1(62779) <= 15310471;
srom_1(62780) <= 14969922;
srom_1(62781) <= 14598512;
srom_1(62782) <= 14197981;
srom_1(62783) <= 13770208;
srom_1(62784) <= 13317198;
srom_1(62785) <= 12841077;
srom_1(62786) <= 12344077;
srom_1(62787) <= 11828528;
srom_1(62788) <= 11296848;
srom_1(62789) <= 10751530;
srom_1(62790) <= 10195132;
srom_1(62791) <= 9630262;
srom_1(62792) <= 9059570;
srom_1(62793) <= 8485732;
srom_1(62794) <= 7911438;
srom_1(62795) <= 7339381;
srom_1(62796) <= 6772245;
srom_1(62797) <= 6212688;
srom_1(62798) <= 5663335;
srom_1(62799) <= 5126762;
srom_1(62800) <= 4605485;
srom_1(62801) <= 4101948;
srom_1(62802) <= 3618513;
srom_1(62803) <= 3157446;
srom_1(62804) <= 2720910;
srom_1(62805) <= 2310952;
srom_1(62806) <= 1929494;
srom_1(62807) <= 1578325;
srom_1(62808) <= 1259092;
srom_1(62809) <= 973291;
srom_1(62810) <= 722263;
srom_1(62811) <= 507186;
srom_1(62812) <= 329067;
srom_1(62813) <= 188742;
srom_1(62814) <= 86870;
srom_1(62815) <= 23927;
srom_1(62816) <= 208;
srom_1(62817) <= 15826;
srom_1(62818) <= 70707;
srom_1(62819) <= 164593;
srom_1(62820) <= 297044;
srom_1(62821) <= 467440;
srom_1(62822) <= 674980;
srom_1(62823) <= 918693;
srom_1(62824) <= 1197434;
srom_1(62825) <= 1509897;
srom_1(62826) <= 1854617;
srom_1(62827) <= 2229977;
srom_1(62828) <= 2634217;
srom_1(62829) <= 3065442;
srom_1(62830) <= 3521628;
srom_1(62831) <= 4000637;
srom_1(62832) <= 4500223;
srom_1(62833) <= 5018043;
srom_1(62834) <= 5551669;
srom_1(62835) <= 6098598;
srom_1(62836) <= 6656266;
srom_1(62837) <= 7222057;
srom_1(62838) <= 7793319;
srom_1(62839) <= 8367372;
srom_1(62840) <= 8941525;
srom_1(62841) <= 9513085;
srom_1(62842) <= 10079371;
srom_1(62843) <= 10637730;
srom_1(62844) <= 11185541;
srom_1(62845) <= 11720237;
srom_1(62846) <= 12239309;
srom_1(62847) <= 12740324;
srom_1(62848) <= 13220933;
srom_1(62849) <= 13678881;
srom_1(62850) <= 14112021;
srom_1(62851) <= 14518322;
srom_1(62852) <= 14895878;
srom_1(62853) <= 15242920;
srom_1(62854) <= 15557820;
srom_1(62855) <= 15839101;
srom_1(62856) <= 16085443;
srom_1(62857) <= 16295693;
srom_1(62858) <= 16468864;
srom_1(62859) <= 16604143;
srom_1(62860) <= 16700897;
srom_1(62861) <= 16758672;
srom_1(62862) <= 16777197;
srom_1(62863) <= 16756385;
srom_1(62864) <= 16696333;
srom_1(62865) <= 16597324;
srom_1(62866) <= 16459821;
srom_1(62867) <= 16284469;
srom_1(62868) <= 16072091;
srom_1(62869) <= 15823683;
srom_1(62870) <= 15540409;
srom_1(62871) <= 15223597;
srom_1(62872) <= 14874734;
srom_1(62873) <= 14495455;
srom_1(62874) <= 14087540;
srom_1(62875) <= 13652900;
srom_1(62876) <= 13193573;
srom_1(62877) <= 12711715;
srom_1(62878) <= 12209584;
srom_1(62879) <= 11689536;
srom_1(62880) <= 11154008;
srom_1(62881) <= 10605512;
srom_1(62882) <= 10046620;
srom_1(62883) <= 9479954;
srom_1(62884) <= 8908169;
srom_1(62885) <= 8333949;
srom_1(62886) <= 7759984;
srom_1(62887) <= 7188968;
srom_1(62888) <= 6623577;
srom_1(62889) <= 6066462;
srom_1(62890) <= 5520237;
srom_1(62891) <= 4987463;
srom_1(62892) <= 4470638;
srom_1(62893) <= 3972186;
srom_1(62894) <= 3494444;
srom_1(62895) <= 3039652;
srom_1(62896) <= 2609943;
srom_1(62897) <= 2207333;
srom_1(62898) <= 1833708;
srom_1(62899) <= 1490822;
srom_1(62900) <= 1180282;
srom_1(62901) <= 903544;
srom_1(62902) <= 661906;
srom_1(62903) <= 456501;
srom_1(62904) <= 288293;
srom_1(62905) <= 158070;
srom_1(62906) <= 66442;
srom_1(62907) <= 13840;
srom_1(62908) <= 511;
srom_1(62909) <= 26516;
srom_1(62910) <= 91733;
srom_1(62911) <= 195858;
srom_1(62912) <= 338401;
srom_1(62913) <= 518694;
srom_1(62914) <= 735892;
srom_1(62915) <= 988977;
srom_1(62916) <= 1276760;
srom_1(62917) <= 1597894;
srom_1(62918) <= 1950871;
srom_1(62919) <= 2334038;
srom_1(62920) <= 2745596;
srom_1(62921) <= 3183616;
srom_1(62922) <= 3646044;
srom_1(62923) <= 4130712;
srom_1(62924) <= 4635347;
srom_1(62925) <= 5157581;
srom_1(62926) <= 5694968;
srom_1(62927) <= 6244985;
srom_1(62928) <= 6805055;
srom_1(62929) <= 7372551;
srom_1(62930) <= 7944811;
srom_1(62931) <= 8519152;
srom_1(62932) <= 9092881;
srom_1(62933) <= 9663308;
srom_1(62934) <= 10227757;
srom_1(62935) <= 10783582;
srom_1(62936) <= 11328175;
srom_1(62937) <= 11858985;
srom_1(62938) <= 12373520;
srom_1(62939) <= 12869369;
srom_1(62940) <= 13344205;
srom_1(62941) <= 13795804;
srom_1(62942) <= 14222046;
srom_1(62943) <= 14620933;
srom_1(62944) <= 14990595;
srom_1(62945) <= 15329298;
srom_1(62946) <= 15635453;
srom_1(62947) <= 15907625;
srom_1(62948) <= 16144538;
srom_1(62949) <= 16345081;
srom_1(62950) <= 16508314;
srom_1(62951) <= 16633470;
srom_1(62952) <= 16719963;
srom_1(62953) <= 16767388;
srom_1(62954) <= 16775521;
srom_1(62955) <= 16744326;
srom_1(62956) <= 16673947;
srom_1(62957) <= 16564716;
srom_1(62958) <= 16417145;
srom_1(62959) <= 16231924;
srom_1(62960) <= 16009924;
srom_1(62961) <= 15752185;
srom_1(62962) <= 15459915;
srom_1(62963) <= 15134485;
srom_1(62964) <= 14777422;
srom_1(62965) <= 14390400;
srom_1(62966) <= 13975233;
srom_1(62967) <= 13533868;
srom_1(62968) <= 13068376;
srom_1(62969) <= 12580938;
srom_1(62970) <= 12073841;
srom_1(62971) <= 11549463;
srom_1(62972) <= 11010262;
srom_1(62973) <= 10458768;
srom_1(62974) <= 9897566;
srom_1(62975) <= 9329288;
srom_1(62976) <= 8756599;
srom_1(62977) <= 8182184;
srom_1(62978) <= 7608737;
srom_1(62979) <= 7038947;
srom_1(62980) <= 6475486;
srom_1(62981) <= 5920997;
srom_1(62982) <= 5378078;
srom_1(62983) <= 4849278;
srom_1(62984) <= 4337074;
srom_1(62985) <= 3843870;
srom_1(62986) <= 3371977;
srom_1(62987) <= 2923609;
srom_1(62988) <= 2500868;
srom_1(62989) <= 2105737;
srom_1(62990) <= 1740069;
srom_1(62991) <= 1405577;
srom_1(62992) <= 1103832;
srom_1(62993) <= 836247;
srom_1(62994) <= 604078;
srom_1(62995) <= 408413;
srom_1(62996) <= 250170;
srom_1(62997) <= 130091;
srom_1(62998) <= 48739;
srom_1(62999) <= 6496;
srom_1(63000) <= 3559;
srom_1(63001) <= 39943;
srom_1(63002) <= 115476;
srom_1(63003) <= 229805;
srom_1(63004) <= 382393;
srom_1(63005) <= 572525;
srom_1(63006) <= 799310;
srom_1(63007) <= 1061683;
srom_1(63008) <= 1358415;
srom_1(63009) <= 1688113;
srom_1(63010) <= 2049233;
srom_1(63011) <= 2440080;
srom_1(63012) <= 2858822;
srom_1(63013) <= 3303495;
srom_1(63014) <= 3772013;
srom_1(63015) <= 4262181;
srom_1(63016) <= 4771699;
srom_1(63017) <= 5298177;
srom_1(63018) <= 5839148;
srom_1(63019) <= 6392074;
srom_1(63020) <= 6954362;
srom_1(63021) <= 7523377;
srom_1(63022) <= 8096448;
srom_1(63023) <= 8670890;
srom_1(63024) <= 9244007;
srom_1(63025) <= 9813114;
srom_1(63026) <= 10375540;
srom_1(63027) <= 10928649;
srom_1(63028) <= 11469847;
srom_1(63029) <= 11996596;
srom_1(63030) <= 12506426;
srom_1(63031) <= 12996946;
srom_1(63032) <= 13465856;
srom_1(63033) <= 13910957;
srom_1(63034) <= 14330162;
srom_1(63035) <= 14721504;
srom_1(63036) <= 15083150;
srom_1(63037) <= 15413403;
srom_1(63038) <= 15710713;
srom_1(63039) <= 15973688;
srom_1(63040) <= 16201094;
srom_1(63041) <= 16391865;
srom_1(63042) <= 16545105;
srom_1(63043) <= 16660097;
srom_1(63044) <= 16736301;
srom_1(63045) <= 16773360;
srom_1(63046) <= 16771100;
srom_1(63047) <= 16729531;
srom_1(63048) <= 16648849;
srom_1(63049) <= 16529432;
srom_1(63050) <= 16371840;
srom_1(63051) <= 16176811;
srom_1(63052) <= 15945261;
srom_1(63053) <= 15678276;
srom_1(63054) <= 15377106;
srom_1(63055) <= 15043165;
srom_1(63056) <= 14678019;
srom_1(63057) <= 14283379;
srom_1(63058) <= 13861097;
srom_1(63059) <= 13413152;
srom_1(63060) <= 12941646;
srom_1(63061) <= 12448788;
srom_1(63062) <= 11936891;
srom_1(63063) <= 11408355;
srom_1(63064) <= 10865659;
srom_1(63065) <= 10311346;
srom_1(63066) <= 9748018;
srom_1(63067) <= 9178314;
srom_1(63068) <= 8604907;
srom_1(63069) <= 8030486;
srom_1(63070) <= 7457745;
srom_1(63071) <= 6889368;
srom_1(63072) <= 6328022;
srom_1(63073) <= 5776339;
srom_1(63074) <= 5236905;
srom_1(63075) <= 4712251;
srom_1(63076) <= 4204837;
srom_1(63077) <= 3717041;
srom_1(63078) <= 3251153;
srom_1(63079) <= 2809355;
srom_1(63080) <= 2393721;
srom_1(63081) <= 2006199;
srom_1(63082) <= 1648606;
srom_1(63083) <= 1322619;
srom_1(63084) <= 1029767;
srom_1(63085) <= 771423;
srom_1(63086) <= 548799;
srom_1(63087) <= 362938;
srom_1(63088) <= 214712;
srom_1(63089) <= 104817;
srom_1(63090) <= 33767;
srom_1(63091) <= 1896;
srom_1(63092) <= 9353;
srom_1(63093) <= 56103;
srom_1(63094) <= 141927;
srom_1(63095) <= 266423;
srom_1(63096) <= 429007;
srom_1(63097) <= 628915;
srom_1(63098) <= 865212;
srom_1(63099) <= 1136788;
srom_1(63100) <= 1442371;
srom_1(63101) <= 1780527;
srom_1(63102) <= 2149670;
srom_1(63103) <= 2548070;
srom_1(63104) <= 2973858;
srom_1(63105) <= 3425038;
srom_1(63106) <= 3899494;
srom_1(63107) <= 4395001;
srom_1(63108) <= 4909235;
srom_1(63109) <= 5439785;
srom_1(63110) <= 5984163;
srom_1(63111) <= 6539817;
srom_1(63112) <= 7104140;
srom_1(63113) <= 7674486;
srom_1(63114) <= 8248181;
srom_1(63115) <= 8822535;
srom_1(63116) <= 9394853;
srom_1(63117) <= 9962453;
srom_1(63118) <= 10522673;
srom_1(63119) <= 11072886;
srom_1(63120) <= 11610510;
srom_1(63121) <= 12133027;
srom_1(63122) <= 12637984;
srom_1(63123) <= 13123015;
srom_1(63124) <= 13585844;
srom_1(63125) <= 14024302;
srom_1(63126) <= 14436332;
srom_1(63127) <= 14820002;
srom_1(63128) <= 15173513;
srom_1(63129) <= 15495208;
srom_1(63130) <= 15783577;
srom_1(63131) <= 16037268;
srom_1(63132) <= 16255093;
srom_1(63133) <= 16436028;
srom_1(63134) <= 16579227;
srom_1(63135) <= 16684017;
srom_1(63136) <= 16749907;
srom_1(63137) <= 16776587;
srom_1(63138) <= 16763934;
srom_1(63139) <= 16712006;
srom_1(63140) <= 16621047;
srom_1(63141) <= 16491483;
srom_1(63142) <= 16323922;
srom_1(63143) <= 16119149;
srom_1(63144) <= 15878125;
srom_1(63145) <= 15601980;
srom_1(63146) <= 15292010;
srom_1(63147) <= 14949666;
srom_1(63148) <= 14576556;
srom_1(63149) <= 14174429;
srom_1(63150) <= 13745169;
srom_1(63151) <= 13290791;
srom_1(63152) <= 12813425;
srom_1(63153) <= 12315309;
srom_1(63154) <= 11798780;
srom_1(63155) <= 11266259;
srom_1(63156) <= 10720244;
srom_1(63157) <= 10163295;
srom_1(63158) <= 9598024;
srom_1(63159) <= 9027082;
srom_1(63160) <= 8453145;
srom_1(63161) <= 7878906;
srom_1(63162) <= 7307057;
srom_1(63163) <= 6740280;
srom_1(63164) <= 6181232;
srom_1(63165) <= 5632536;
srom_1(63166) <= 5096764;
srom_1(63167) <= 4576428;
srom_1(63168) <= 4073969;
srom_1(63169) <= 3591742;
srom_1(63170) <= 3132010;
srom_1(63171) <= 2696928;
srom_1(63172) <= 2288536;
srom_1(63173) <= 1908750;
srom_1(63174) <= 1559349;
srom_1(63175) <= 1241974;
srom_1(63176) <= 958111;
srom_1(63177) <= 709093;
srom_1(63178) <= 496086;
srom_1(63179) <= 320090;
srom_1(63180) <= 181930;
srom_1(63181) <= 82255;
srom_1(63182) <= 21530;
srom_1(63183) <= 42;
srom_1(63184) <= 17890;
srom_1(63185) <= 74992;
srom_1(63186) <= 171079;
srom_1(63187) <= 305701;
srom_1(63188) <= 478226;
srom_1(63189) <= 687846;
srom_1(63190) <= 933577;
srom_1(63191) <= 1214268;
srom_1(63192) <= 1528601;
srom_1(63193) <= 1875103;
srom_1(63194) <= 2252150;
srom_1(63195) <= 2657972;
srom_1(63196) <= 3090668;
srom_1(63197) <= 3548207;
srom_1(63198) <= 4028444;
srom_1(63199) <= 4529128;
srom_1(63200) <= 5047910;
srom_1(63201) <= 5582358;
srom_1(63202) <= 6129965;
srom_1(63203) <= 6688164;
srom_1(63204) <= 7254337;
srom_1(63205) <= 7825829;
srom_1(63206) <= 8399960;
srom_1(63207) <= 8974037;
srom_1(63208) <= 9545370;
srom_1(63209) <= 10111278;
srom_1(63210) <= 10669107;
srom_1(63211) <= 11216243;
srom_1(63212) <= 11750119;
srom_1(63213) <= 12268231;
srom_1(63214) <= 12768151;
srom_1(63215) <= 13247534;
srom_1(63216) <= 13704131;
srom_1(63217) <= 14135802;
srom_1(63218) <= 14540522;
srom_1(63219) <= 14916394;
srom_1(63220) <= 15261655;
srom_1(63221) <= 15574686;
srom_1(63222) <= 15854019;
srom_1(63223) <= 16098344;
srom_1(63224) <= 16306515;
srom_1(63225) <= 16477557;
srom_1(63226) <= 16610667;
srom_1(63227) <= 16705220;
srom_1(63228) <= 16760774;
srom_1(63229) <= 16777069;
srom_1(63230) <= 16754026;
srom_1(63231) <= 16691756;
srom_1(63232) <= 16590549;
srom_1(63233) <= 16450881;
srom_1(63234) <= 16273405;
srom_1(63235) <= 16058955;
srom_1(63236) <= 15808537;
srom_1(63237) <= 15523323;
srom_1(63238) <= 15204653;
srom_1(63239) <= 14854020;
srom_1(63240) <= 14473068;
srom_1(63241) <= 14063584;
srom_1(63242) <= 13627488;
srom_1(63243) <= 13166825;
srom_1(63244) <= 12683756;
srom_1(63245) <= 12180545;
srom_1(63246) <= 11659552;
srom_1(63247) <= 11123221;
srom_1(63248) <= 10574066;
srom_1(63249) <= 10014663;
srom_1(63250) <= 9447635;
srom_1(63251) <= 8875640;
srom_1(63252) <= 8301362;
srom_1(63253) <= 7727493;
srom_1(63254) <= 7156724;
srom_1(63255) <= 6591732;
srom_1(63256) <= 6035166;
srom_1(63257) <= 5489636;
srom_1(63258) <= 4957700;
srom_1(63259) <= 4441853;
srom_1(63260) <= 3944513;
srom_1(63261) <= 3468014;
srom_1(63262) <= 3014589;
srom_1(63263) <= 2586364;
srom_1(63264) <= 2185349;
srom_1(63265) <= 1813422;
srom_1(63266) <= 1472329;
srom_1(63267) <= 1163668;
srom_1(63268) <= 888888;
srom_1(63269) <= 649277;
srom_1(63270) <= 445957;
srom_1(63271) <= 279884;
srom_1(63272) <= 151835;
srom_1(63273) <= 62412;
srom_1(63274) <= 12032;
srom_1(63275) <= 934;
srom_1(63276) <= 29168;
srom_1(63277) <= 96602;
srom_1(63278) <= 202920;
srom_1(63279) <= 347624;
srom_1(63280) <= 530035;
srom_1(63281) <= 749297;
srom_1(63282) <= 1004383;
srom_1(63283) <= 1294096;
srom_1(63284) <= 1617077;
srom_1(63285) <= 1971813;
srom_1(63286) <= 2356639;
srom_1(63287) <= 2769751;
srom_1(63288) <= 3209211;
srom_1(63289) <= 3672960;
srom_1(63290) <= 4158822;
srom_1(63291) <= 4664519;
srom_1(63292) <= 5187679;
srom_1(63293) <= 5725850;
srom_1(63294) <= 6276507;
srom_1(63295) <= 6837069;
srom_1(63296) <= 7404906;
srom_1(63297) <= 7977356;
srom_1(63298) <= 8551735;
srom_1(63299) <= 9125349;
srom_1(63300) <= 9695508;
srom_1(63301) <= 10259538;
srom_1(63302) <= 10814795;
srom_1(63303) <= 11358675;
srom_1(63304) <= 11888627;
srom_1(63305) <= 12402166;
srom_1(63306) <= 12896884;
srom_1(63307) <= 13370462;
srom_1(63308) <= 13820677;
srom_1(63309) <= 14245420;
srom_1(63310) <= 14642699;
srom_1(63311) <= 15010649;
srom_1(63312) <= 15347547;
srom_1(63313) <= 15651812;
srom_1(63314) <= 15922017;
srom_1(63315) <= 16156896;
srom_1(63316) <= 16355346;
srom_1(63317) <= 16516437;
srom_1(63318) <= 16639415;
srom_1(63319) <= 16723701;
srom_1(63320) <= 16768901;
srom_1(63321) <= 16774803;
srom_1(63322) <= 16741380;
srom_1(63323) <= 16668787;
srom_1(63324) <= 16557366;
srom_1(63325) <= 16407639;
srom_1(63326) <= 16220308;
srom_1(63327) <= 15996251;
srom_1(63328) <= 15736519;
srom_1(63329) <= 15442330;
srom_1(63330) <= 15115065;
srom_1(63331) <= 14756256;
srom_1(63332) <= 14367587;
srom_1(63333) <= 13950881;
srom_1(63334) <= 13508091;
srom_1(63335) <= 13041295;
srom_1(63336) <= 12552680;
srom_1(63337) <= 12044539;
srom_1(63338) <= 11519253;
srom_1(63339) <= 10979287;
srom_1(63340) <= 10427173;
srom_1(63341) <= 9865498;
srom_1(63342) <= 9296899;
srom_1(63343) <= 8724039;
srom_1(63344) <= 8149607;
srom_1(63345) <= 7576296;
srom_1(63346) <= 7006794;
srom_1(63347) <= 6443772;
srom_1(63348) <= 5889869;
srom_1(63349) <= 5347684;
srom_1(63350) <= 4819759;
srom_1(63351) <= 4308570;
srom_1(63352) <= 3816513;
srom_1(63353) <= 3345897;
srom_1(63354) <= 2898927;
srom_1(63355) <= 2477700;
srom_1(63356) <= 2084192;
srom_1(63357) <= 1720247;
srom_1(63358) <= 1387573;
srom_1(63359) <= 1087728;
srom_1(63360) <= 822120;
srom_1(63361) <= 591994;
srom_1(63362) <= 398429;
srom_1(63363) <= 242333;
srom_1(63364) <= 124437;
srom_1(63365) <= 45295;
srom_1(63366) <= 5277;
srom_1(63367) <= 4572;
srom_1(63368) <= 43182;
srom_1(63369) <= 120927;
srom_1(63370) <= 237442;
srom_1(63371) <= 392180;
srom_1(63372) <= 584417;
srom_1(63373) <= 813250;
srom_1(63374) <= 1077606;
srom_1(63375) <= 1376247;
srom_1(63376) <= 1707770;
srom_1(63377) <= 2070623;
srom_1(63378) <= 2463102;
srom_1(63379) <= 2883369;
srom_1(63380) <= 3329451;
srom_1(63381) <= 3799257;
srom_1(63382) <= 4290585;
srom_1(63383) <= 4801129;
srom_1(63384) <= 5328496;
srom_1(63385) <= 5870214;
srom_1(63386) <= 6423740;
srom_1(63387) <= 6986481;
srom_1(63388) <= 7555797;
srom_1(63389) <= 8129018;
srom_1(63390) <= 8703457;
srom_1(63391) <= 9276419;
srom_1(63392) <= 9845217;
srom_1(63393) <= 10407186;
srom_1(63394) <= 10959688;
srom_1(63395) <= 11500134;
srom_1(63396) <= 12025989;
srom_1(63397) <= 12534786;
srom_1(63398) <= 13024141;
srom_1(63399) <= 13491759;
srom_1(63400) <= 13935445;
srom_1(63401) <= 14353121;
srom_1(63402) <= 14742827;
srom_1(63403) <= 15102736;
srom_1(63404) <= 15431161;
srom_1(63405) <= 15726560;
srom_1(63406) <= 15987549;
srom_1(63407) <= 16212904;
srom_1(63408) <= 16401568;
srom_1(63409) <= 16552657;
srom_1(63410) <= 16665461;
srom_1(63411) <= 16739453;
srom_1(63412) <= 16774284;
srom_1(63413) <= 16769793;
srom_1(63414) <= 16725999;
srom_1(63415) <= 16643108;
srom_1(63416) <= 16521509;
srom_1(63417) <= 16361772;
srom_1(63418) <= 16164646;
srom_1(63419) <= 15931055;
srom_1(63420) <= 15662096;
srom_1(63421) <= 15359028;
srom_1(63422) <= 15023274;
srom_1(63423) <= 14656408;
srom_1(63424) <= 14260149;
srom_1(63425) <= 13836357;
srom_1(63426) <= 13387019;
srom_1(63427) <= 12914241;
srom_1(63428) <= 12420241;
srom_1(63429) <= 11907336;
srom_1(63430) <= 11377930;
srom_1(63431) <= 10834505;
srom_1(63432) <= 10279612;
srom_1(63433) <= 9715850;
srom_1(63434) <= 9145865;
srom_1(63435) <= 8572329;
srom_1(63436) <= 7997931;
srom_1(63437) <= 7425365;
srom_1(63438) <= 6857316;
srom_1(63439) <= 6296448;
srom_1(63440) <= 5745391;
srom_1(63441) <= 5206729;
srom_1(63442) <= 4682987;
srom_1(63443) <= 4176623;
srom_1(63444) <= 3690010;
srom_1(63445) <= 3225430;
srom_1(63446) <= 2785062;
srom_1(63447) <= 2370971;
srom_1(63448) <= 1985099;
srom_1(63449) <= 1629255;
srom_1(63450) <= 1305109;
srom_1(63451) <= 1014179;
srom_1(63452) <= 757830;
srom_1(63453) <= 537264;
srom_1(63454) <= 353517;
srom_1(63455) <= 207448;
srom_1(63456) <= 99744;
srom_1(63457) <= 30909;
srom_1(63458) <= 1266;
srom_1(63459) <= 10955;
srom_1(63460) <= 59929;
srom_1(63461) <= 147959;
srom_1(63462) <= 274632;
srom_1(63463) <= 439355;
srom_1(63464) <= 641354;
srom_1(63465) <= 879683;
srom_1(63466) <= 1153223;
srom_1(63467) <= 1460693;
srom_1(63468) <= 1800651;
srom_1(63469) <= 2171501;
srom_1(63470) <= 2571506;
srom_1(63471) <= 2998789;
srom_1(63472) <= 3451347;
srom_1(63473) <= 3927057;
srom_1(63474) <= 4423689;
srom_1(63475) <= 4938914;
srom_1(63476) <= 5470315;
srom_1(63477) <= 6015402;
srom_1(63478) <= 6571617;
srom_1(63479) <= 7136353;
srom_1(63480) <= 7706961;
srom_1(63481) <= 8280765;
srom_1(63482) <= 8855075;
srom_1(63483) <= 9427198;
srom_1(63484) <= 9994451;
srom_1(63485) <= 10554173;
srom_1(63486) <= 11103740;
srom_1(63487) <= 11640574;
srom_1(63488) <= 12162160;
srom_1(63489) <= 12666049;
srom_1(63490) <= 13149881;
srom_1(63491) <= 13611385;
srom_1(63492) <= 14048397;
srom_1(63493) <= 14458869;
srom_1(63494) <= 14840876;
srom_1(63495) <= 15192625;
srom_1(63496) <= 15512468;
srom_1(63497) <= 15798905;
srom_1(63498) <= 16050593;
srom_1(63499) <= 16266351;
srom_1(63500) <= 16445167;
srom_1(63501) <= 16586203;
srom_1(63502) <= 16688798;
srom_1(63503) <= 16752471;
srom_1(63504) <= 16776922;
srom_1(63505) <= 16762038;
srom_1(63506) <= 16707888;
srom_1(63507) <= 16614726;
srom_1(63508) <= 16482989;
srom_1(63509) <= 16313294;
srom_1(63510) <= 16106438;
srom_1(63511) <= 15863391;
srom_1(63512) <= 15585291;
srom_1(63513) <= 15273444;
srom_1(63514) <= 14929311;
srom_1(63515) <= 14554507;
srom_1(63516) <= 14150789;
srom_1(63517) <= 13720050;
srom_1(63518) <= 13264310;
srom_1(63519) <= 12785706;
srom_1(63520) <= 12286483;
srom_1(63521) <= 11768981;
srom_1(63522) <= 11235627;
srom_1(63523) <= 10688923;
srom_1(63524) <= 10131432;
srom_1(63525) <= 9565768;
srom_1(63526) <= 8994584;
srom_1(63527) <= 8420558;
srom_1(63528) <= 7846382;
srom_1(63529) <= 7274750;
srom_1(63530) <= 6708340;
srom_1(63531) <= 6149810;
srom_1(63532) <= 5601778;
srom_1(63533) <= 5066815;
srom_1(63534) <= 4547428;
srom_1(63535) <= 4046055;
srom_1(63536) <= 3565045;
srom_1(63537) <= 3106654;
srom_1(63538) <= 2673032;
srom_1(63539) <= 2266213;
srom_1(63540) <= 1888103;
srom_1(63541) <= 1540477;
srom_1(63542) <= 1224964;
srom_1(63543) <= 943043;
srom_1(63544) <= 696038;
srom_1(63545) <= 485105;
srom_1(63546) <= 311235;
srom_1(63547) <= 175242;
srom_1(63548) <= 77765;
srom_1(63549) <= 19260;
srom_1(63550) <= 2;
srom_1(63551) <= 20080;
srom_1(63552) <= 79402;
srom_1(63553) <= 177689;
srom_1(63554) <= 314479;
srom_1(63555) <= 489131;
srom_1(63556) <= 700827;
srom_1(63557) <= 948574;
srom_1(63558) <= 1231209;
srom_1(63559) <= 1547408;
srom_1(63560) <= 1895688;
srom_1(63561) <= 2274415;
srom_1(63562) <= 2681814;
srom_1(63563) <= 3115974;
srom_1(63564) <= 3574859;
srom_1(63565) <= 4056317;
srom_1(63566) <= 4558091;
srom_1(63567) <= 5077828;
srom_1(63568) <= 5613089;
srom_1(63569) <= 6161367;
srom_1(63570) <= 6720088;
srom_1(63571) <= 7286634;
srom_1(63572) <= 7858348;
srom_1(63573) <= 8432547;
srom_1(63574) <= 9006541;
srom_1(63575) <= 9577637;
srom_1(63576) <= 10143158;
srom_1(63577) <= 10700451;
srom_1(63578) <= 11246902;
srom_1(63579) <= 11779950;
srom_1(63580) <= 12297095;
srom_1(63581) <= 12795912;
srom_1(63582) <= 13274061;
srom_1(63583) <= 13729301;
srom_1(63584) <= 14159496;
srom_1(63585) <= 14562630;
srom_1(63586) <= 14936812;
srom_1(63587) <= 15280287;
srom_1(63588) <= 15591444;
srom_1(63589) <= 15868825;
srom_1(63590) <= 16111128;
srom_1(63591) <= 16317218;
srom_1(63592) <= 16486128;
srom_1(63593) <= 16617066;
srom_1(63594) <= 16709418;
srom_1(63595) <= 16762750;
srom_1(63596) <= 16776814;
srom_1(63597) <= 16751542;
srom_1(63598) <= 16687054;
srom_1(63599) <= 16583651;
srom_1(63600) <= 16441819;
srom_1(63601) <= 16262222;
srom_1(63602) <= 16045704;
srom_1(63603) <= 15793279;
srom_1(63604) <= 15506130;
srom_1(63605) <= 15185606;
srom_1(63606) <= 14833207;
srom_1(63607) <= 14450588;
srom_1(63608) <= 14039542;
srom_1(63609) <= 13601997;
srom_1(63610) <= 13140005;
srom_1(63611) <= 12655731;
srom_1(63612) <= 12151448;
srom_1(63613) <= 11629519;
srom_1(63614) <= 11092393;
srom_1(63615) <= 10542587;
srom_1(63616) <= 9982681;
srom_1(63617) <= 9415300;
srom_1(63618) <= 8843104;
srom_1(63619) <= 8268777;
srom_1(63620) <= 7695011;
srom_1(63621) <= 7124499;
srom_1(63622) <= 6559914;
srom_1(63623) <= 6003904;
srom_1(63624) <= 5459078;
srom_1(63625) <= 4927988;
srom_1(63626) <= 4413127;
srom_1(63627) <= 3916908;
srom_1(63628) <= 3441659;
srom_1(63629) <= 2989607;
srom_1(63630) <= 2562873;
srom_1(63631) <= 2163458;
srom_1(63632) <= 1793235;
srom_1(63633) <= 1453940;
srom_1(63634) <= 1147164;
srom_1(63635) <= 874345;
srom_1(63636) <= 636764;
srom_1(63637) <= 435533;
srom_1(63638) <= 271598;
srom_1(63639) <= 145725;
srom_1(63640) <= 58507;
srom_1(63641) <= 10351;
srom_1(63642) <= 1483;
srom_1(63643) <= 31946;
srom_1(63644) <= 101596;
srom_1(63645) <= 210106;
srom_1(63646) <= 356969;
srom_1(63647) <= 541494;
srom_1(63648) <= 762818;
srom_1(63649) <= 1019901;
srom_1(63650) <= 1311538;
srom_1(63651) <= 1636363;
srom_1(63652) <= 1992851;
srom_1(63653) <= 2379331;
srom_1(63654) <= 2793990;
srom_1(63655) <= 3234885;
srom_1(63656) <= 3699947;
srom_1(63657) <= 4186996;
srom_1(63658) <= 4693747;
srom_1(63659) <= 5217825;
srom_1(63660) <= 5756772;
srom_1(63661) <= 6308061;
srom_1(63662) <= 6869106;
srom_1(63663) <= 7437276;
srom_1(63664) <= 8009908;
srom_1(63665) <= 8584315;
srom_1(63666) <= 9157805;
srom_1(63667) <= 9727688;
srom_1(63668) <= 10291291;
srom_1(63669) <= 10845972;
srom_1(63670) <= 11389129;
srom_1(63671) <= 11918216;
srom_1(63672) <= 12430751;
srom_1(63673) <= 12924332;
srom_1(63674) <= 13396642;
srom_1(63675) <= 13845469;
srom_1(63676) <= 14268706;
srom_1(63677) <= 14664370;
srom_1(63678) <= 15030604;
srom_1(63679) <= 15365692;
srom_1(63680) <= 15668061;
srom_1(63681) <= 15936295;
srom_1(63682) <= 16169135;
srom_1(63683) <= 16365490;
srom_1(63684) <= 16524438;
srom_1(63685) <= 16645235;
srom_1(63686) <= 16727313;
srom_1(63687) <= 16770288;
srom_1(63688) <= 16773959;
srom_1(63689) <= 16738308;
srom_1(63690) <= 16663502;
srom_1(63691) <= 16549893;
srom_1(63692) <= 16398012;
srom_1(63693) <= 16208573;
srom_1(63694) <= 15982463;
srom_1(63695) <= 15720743;
srom_1(63696) <= 15424639;
srom_1(63697) <= 15095542;
srom_1(63698) <= 14734993;
srom_1(63699) <= 14344684;
srom_1(63700) <= 13926445;
srom_1(63701) <= 13482238;
srom_1(63702) <= 13014144;
srom_1(63703) <= 12524359;
srom_1(63704) <= 12015181;
srom_1(63705) <= 11488996;
srom_1(63706) <= 10948273;
srom_1(63707) <= 10395546;
srom_1(63708) <= 9833409;
srom_1(63709) <= 9264496;
srom_1(63710) <= 8691475;
srom_1(63711) <= 8117035;
srom_1(63712) <= 7543868;
srom_1(63713) <= 6974662;
srom_1(63714) <= 6412086;
srom_1(63715) <= 5858780;
srom_1(63716) <= 5317336;
srom_1(63717) <= 4790295;
srom_1(63718) <= 4280127;
srom_1(63719) <= 3789226;
srom_1(63720) <= 3319892;
srom_1(63721) <= 2874328;
srom_1(63722) <= 2454622;
srom_1(63723) <= 2062742;
srom_1(63724) <= 1700526;
srom_1(63725) <= 1369674;
srom_1(63726) <= 1071735;
srom_1(63727) <= 808108;
srom_1(63728) <= 580028;
srom_1(63729) <= 388565;
srom_1(63730) <= 234618;
srom_1(63731) <= 118907;
srom_1(63732) <= 41976;
srom_1(63733) <= 4185;
srom_1(63734) <= 5711;
srom_1(63735) <= 46547;
srom_1(63736) <= 126503;
srom_1(63737) <= 245202;
srom_1(63738) <= 402088;
srom_1(63739) <= 596426;
srom_1(63740) <= 827304;
srom_1(63741) <= 1093640;
srom_1(63742) <= 1394185;
srom_1(63743) <= 1727528;
srom_1(63744) <= 2092108;
srom_1(63745) <= 2486214;
srom_1(63746) <= 2907998;
srom_1(63747) <= 3355483;
srom_1(63748) <= 3826570;
srom_1(63749) <= 4319050;
srom_1(63750) <= 4830613;
srom_1(63751) <= 5358861;
srom_1(63752) <= 5901317;
srom_1(63753) <= 6455436;
srom_1(63754) <= 7018621;
srom_1(63755) <= 7588230;
srom_1(63756) <= 8161592;
srom_1(63757) <= 8736019;
srom_1(63758) <= 9308817;
srom_1(63759) <= 9877299;
srom_1(63760) <= 10438801;
srom_1(63761) <= 10990688;
srom_1(63762) <= 11530373;
srom_1(63763) <= 12055326;
srom_1(63764) <= 12563084;
srom_1(63765) <= 13051266;
srom_1(63766) <= 13517584;
srom_1(63767) <= 13959850;
srom_1(63768) <= 14375991;
srom_1(63769) <= 14764055;
srom_1(63770) <= 15122222;
srom_1(63771) <= 15448812;
srom_1(63772) <= 15742296;
srom_1(63773) <= 16001295;
srom_1(63774) <= 16224595;
srom_1(63775) <= 16411150;
srom_1(63776) <= 16560085;
srom_1(63777) <= 16670700;
srom_1(63778) <= 16742478;
srom_1(63779) <= 16775082;
srom_1(63780) <= 16768359;
srom_1(63781) <= 16722340;
srom_1(63782) <= 16637242;
srom_1(63783) <= 16513463;
srom_1(63784) <= 16351583;
srom_1(63785) <= 16152363;
srom_1(63786) <= 15916735;
srom_1(63787) <= 15645806;
srom_1(63788) <= 15340845;
srom_1(63789) <= 15003283;
srom_1(63790) <= 14634702;
srom_1(63791) <= 14236831;
srom_1(63792) <= 13811536;
srom_1(63793) <= 13360810;
srom_1(63794) <= 12886769;
srom_1(63795) <= 12391634;
srom_1(63796) <= 11877727;
srom_1(63797) <= 11347459;
srom_1(63798) <= 10803315;
srom_1(63799) <= 10247848;
srom_1(63800) <= 9683663;
srom_1(63801) <= 9113405;
srom_1(63802) <= 8539747;
srom_1(63803) <= 7965382;
srom_1(63804) <= 7393000;
srom_1(63805) <= 6825288;
srom_1(63806) <= 6264906;
srom_1(63807) <= 5714483;
srom_1(63808) <= 5176600;
srom_1(63809) <= 4653779;
srom_1(63810) <= 4148473;
srom_1(63811) <= 3663049;
srom_1(63812) <= 3199785;
srom_1(63813) <= 2760854;
srom_1(63814) <= 2348313;
srom_1(63815) <= 1964097;
srom_1(63816) <= 1610007;
srom_1(63817) <= 1287705;
srom_1(63818) <= 998702;
srom_1(63819) <= 744352;
srom_1(63820) <= 525849;
srom_1(63821) <= 344217;
srom_1(63822) <= 200308;
srom_1(63823) <= 94796;
srom_1(63824) <= 28177;
srom_1(63825) <= 763;
srom_1(63826) <= 12683;
srom_1(63827) <= 63880;
srom_1(63828) <= 154115;
srom_1(63829) <= 282964;
srom_1(63830) <= 449823;
srom_1(63831) <= 653909;
srom_1(63832) <= 894267;
srom_1(63833) <= 1169768;
srom_1(63834) <= 1479121;
srom_1(63835) <= 1820874;
srom_1(63836) <= 2193426;
srom_1(63837) <= 2595029;
srom_1(63838) <= 3023801;
srom_1(63839) <= 3477729;
srom_1(63840) <= 3954687;
srom_1(63841) <= 4452437;
srom_1(63842) <= 4968644;
srom_1(63843) <= 5500889;
srom_1(63844) <= 6046676;
srom_1(63845) <= 6603445;
srom_1(63846) <= 7168585;
srom_1(63847) <= 7739446;
srom_1(63848) <= 8313351;
srom_1(63849) <= 8887609;
srom_1(63850) <= 9459527;
srom_1(63851) <= 10026423;
srom_1(63852) <= 10585639;
srom_1(63853) <= 11134553;
srom_1(63854) <= 11670589;
srom_1(63855) <= 12191236;
srom_1(63856) <= 12694050;
srom_1(63857) <= 13176675;
srom_1(63858) <= 13636846;
srom_1(63859) <= 14072407;
srom_1(63860) <= 14481315;
srom_1(63861) <= 14861652;
srom_1(63862) <= 15211635;
srom_1(63863) <= 15529622;
srom_1(63864) <= 15814122;
srom_1(63865) <= 16063802;
srom_1(63866) <= 16277490;
srom_1(63867) <= 16454184;
srom_1(63868) <= 16593056;
srom_1(63869) <= 16693455;
srom_1(63870) <= 16754909;
srom_1(63871) <= 16777131;
srom_1(63872) <= 16760016;
srom_1(63873) <= 16703644;
srom_1(63874) <= 16608281;
srom_1(63875) <= 16474373;
srom_1(63876) <= 16302548;
srom_1(63877) <= 16093611;
srom_1(63878) <= 15848543;
srom_1(63879) <= 15568493;
srom_1(63880) <= 15254774;
srom_1(63881) <= 14908858;
srom_1(63882) <= 14532365;
srom_1(63883) <= 14127062;
srom_1(63884) <= 13694850;
srom_1(63885) <= 13237755;
srom_1(63886) <= 12757921;
srom_1(63887) <= 12257597;
srom_1(63888) <= 11739131;
srom_1(63889) <= 11204952;
srom_1(63890) <= 10657567;
srom_1(63891) <= 10099542;
srom_1(63892) <= 9533494;
srom_1(63893) <= 8962077;
srom_1(63894) <= 8387970;
srom_1(63895) <= 7813867;
srom_1(63896) <= 7242459;
srom_1(63897) <= 6676425;
srom_1(63898) <= 6118421;
srom_1(63899) <= 5571062;
srom_1(63900) <= 5036916;
srom_1(63901) <= 4518487;
srom_1(63902) <= 4018206;
srom_1(63903) <= 3538420;
srom_1(63904) <= 3081377;
srom_1(63905) <= 2649222;
srom_1(63906) <= 2243981;
srom_1(63907) <= 1867555;
srom_1(63908) <= 1521708;
srom_1(63909) <= 1208062;
srom_1(63910) <= 928088;
srom_1(63911) <= 683099;
srom_1(63912) <= 474244;
srom_1(63913) <= 302502;
srom_1(63914) <= 168678;
srom_1(63915) <= 73401;
srom_1(63916) <= 17116;
srom_1(63917) <= 88;
srom_1(63918) <= 22397;
srom_1(63919) <= 83938;
srom_1(63920) <= 184422;
srom_1(63921) <= 323379;
srom_1(63922) <= 500156;
srom_1(63923) <= 713925;
srom_1(63924) <= 963683;
srom_1(63925) <= 1248259;
srom_1(63926) <= 1566319;
srom_1(63927) <= 1916370;
srom_1(63928) <= 2296773;
srom_1(63929) <= 2705741;
srom_1(63930) <= 3141359;
srom_1(63931) <= 3601583;
srom_1(63932) <= 4084255;
srom_1(63933) <= 4587112;
srom_1(63934) <= 5107795;
srom_1(63935) <= 5643863;
srom_1(63936) <= 6192802;
srom_1(63937) <= 6752038;
srom_1(63938) <= 7318948;
srom_1(63939) <= 7890874;
srom_1(63940) <= 8465134;
srom_1(63941) <= 9039036;
srom_1(63942) <= 9609887;
srom_1(63943) <= 10175012;
srom_1(63944) <= 10731759;
srom_1(63945) <= 11277518;
srom_1(63946) <= 11809731;
srom_1(63947) <= 12325900;
srom_1(63948) <= 12823606;
srom_1(63949) <= 13300515;
srom_1(63950) <= 13754391;
srom_1(63951) <= 14183104;
srom_1(63952) <= 14584645;
srom_1(63953) <= 14957130;
srom_1(63954) <= 15298814;
srom_1(63955) <= 15608093;
srom_1(63956) <= 15883518;
srom_1(63957) <= 16123796;
srom_1(63958) <= 16327801;
srom_1(63959) <= 16494577;
srom_1(63960) <= 16623341;
srom_1(63961) <= 16713490;
srom_1(63962) <= 16764600;
srom_1(63963) <= 16776432;
srom_1(63964) <= 16748931;
srom_1(63965) <= 16682226;
srom_1(63966) <= 16576629;
srom_1(63967) <= 16432635;
srom_1(63968) <= 16250921;
srom_1(63969) <= 16032337;
srom_1(63970) <= 15777909;
srom_1(63971) <= 15488830;
srom_1(63972) <= 15166456;
srom_1(63973) <= 14812298;
srom_1(63974) <= 14428017;
srom_1(63975) <= 14015415;
srom_1(63976) <= 13576428;
srom_1(63977) <= 13113112;
srom_1(63978) <= 12627642;
srom_1(63979) <= 12122294;
srom_1(63980) <= 11599437;
srom_1(63981) <= 11061524;
srom_1(63982) <= 10511076;
srom_1(63983) <= 9950675;
srom_1(63984) <= 9382949;
srom_1(63985) <= 8810561;
srom_1(63986) <= 8236193;
srom_1(63987) <= 7662541;
srom_1(63988) <= 7092293;
srom_1(63989) <= 6528124;
srom_1(63990) <= 5972679;
srom_1(63991) <= 5428564;
srom_1(63992) <= 4898329;
srom_1(63993) <= 4384461;
srom_1(63994) <= 3889370;
srom_1(63995) <= 3415378;
srom_1(63996) <= 2964707;
srom_1(63997) <= 2539470;
srom_1(63998) <= 2141662;
srom_1(63999) <= 1773148;
srom_1(64000) <= 1435656;
srom_1(64001) <= 1130769;
srom_1(64002) <= 859916;
srom_1(64003) <= 624368;
srom_1(64004) <= 425230;
srom_1(64005) <= 263434;
srom_1(64006) <= 139740;
srom_1(64007) <= 54727;
srom_1(64008) <= 8796;
srom_1(64009) <= 2159;
srom_1(64010) <= 34850;
srom_1(64011) <= 106715;
srom_1(64012) <= 217416;
srom_1(64013) <= 366435;
srom_1(64014) <= 553072;
srom_1(64015) <= 776453;
srom_1(64016) <= 1035530;
srom_1(64017) <= 1329088;
srom_1(64018) <= 1655750;
srom_1(64019) <= 2013986;
srom_1(64020) <= 2402114;
srom_1(64021) <= 2818314;
srom_1(64022) <= 3260636;
srom_1(64023) <= 3727004;
srom_1(64024) <= 4215233;
srom_1(64025) <= 4723032;
srom_1(64026) <= 5248019;
srom_1(64027) <= 5787735;
srom_1(64028) <= 6339646;
srom_1(64029) <= 6901166;
srom_1(64030) <= 7469661;
srom_1(64031) <= 8042465;
srom_1(64032) <= 8616893;
srom_1(64033) <= 9190250;
srom_1(64034) <= 9759847;
srom_1(64035) <= 10323015;
srom_1(64036) <= 10877111;
srom_1(64037) <= 11419538;
srom_1(64038) <= 11947752;
srom_1(64039) <= 12459276;
srom_1(64040) <= 12951711;
srom_1(64041) <= 13422748;
srom_1(64042) <= 13870178;
srom_1(64043) <= 14291903;
srom_1(64044) <= 14685946;
srom_1(64045) <= 15050458;
srom_1(64046) <= 15383731;
srom_1(64047) <= 15684201;
srom_1(64048) <= 15950459;
srom_1(64049) <= 16181258;
srom_1(64050) <= 16375514;
srom_1(64051) <= 16532316;
srom_1(64052) <= 16650930;
srom_1(64053) <= 16730799;
srom_1(64054) <= 16771549;
srom_1(64055) <= 16772988;
srom_1(64056) <= 16735110;
srom_1(64057) <= 16658092;
srom_1(64058) <= 16542296;
srom_1(64059) <= 16388265;
srom_1(64060) <= 16196720;
srom_1(64061) <= 15968560;
srom_1(64062) <= 15704855;
srom_1(64063) <= 15406842;
srom_1(64064) <= 15075918;
srom_1(64065) <= 14713635;
srom_1(64066) <= 14321692;
srom_1(64067) <= 13901926;
srom_1(64068) <= 13456307;
srom_1(64069) <= 12986923;
srom_1(64070) <= 12495976;
srom_1(64071) <= 11985769;
srom_1(64072) <= 11458693;
srom_1(64073) <= 10917220;
srom_1(64074) <= 10363890;
srom_1(64075) <= 9801297;
srom_1(64076) <= 9232079;
srom_1(64077) <= 8658906;
srom_1(64078) <= 8084466;
srom_1(64079) <= 7511452;
srom_1(64080) <= 6942551;
srom_1(64081) <= 6380431;
srom_1(64082) <= 5827728;
srom_1(64083) <= 5287034;
srom_1(64084) <= 4760885;
srom_1(64085) <= 4251747;
srom_1(64086) <= 3762008;
srom_1(64087) <= 3293964;
srom_1(64088) <= 2849812;
srom_1(64089) <= 2431633;
srom_1(64090) <= 2041387;
srom_1(64091) <= 1680907;
srom_1(64092) <= 1351881;
srom_1(64093) <= 1055852;
srom_1(64094) <= 794210;
srom_1(64095) <= 568180;
srom_1(64096) <= 378823;
srom_1(64097) <= 227026;
srom_1(64098) <= 113502;
srom_1(64099) <= 38783;
srom_1(64100) <= 3219;
srom_1(64101) <= 6976;
srom_1(64102) <= 50039;
srom_1(64103) <= 132203;
srom_1(64104) <= 253085;
srom_1(64105) <= 412117;
srom_1(64106) <= 608553;
srom_1(64107) <= 841473;
srom_1(64108) <= 1109784;
srom_1(64109) <= 1412228;
srom_1(64110) <= 1747386;
srom_1(64111) <= 2113688;
srom_1(64112) <= 2509414;
srom_1(64113) <= 2932711;
srom_1(64114) <= 3381591;
srom_1(64115) <= 3853952;
srom_1(64116) <= 4347577;
srom_1(64117) <= 4860151;
srom_1(64118) <= 5389272;
srom_1(64119) <= 5932458;
srom_1(64120) <= 6487162;
srom_1(64121) <= 7050782;
srom_1(64122) <= 7620675;
srom_1(64123) <= 8194170;
srom_1(64124) <= 8768576;
srom_1(64125) <= 9341201;
srom_1(64126) <= 9909358;
srom_1(64127) <= 10470385;
srom_1(64128) <= 11021649;
srom_1(64129) <= 11560566;
srom_1(64130) <= 12084608;
srom_1(64131) <= 12591319;
srom_1(64132) <= 13078321;
srom_1(64133) <= 13543332;
srom_1(64134) <= 13984171;
srom_1(64135) <= 14398770;
srom_1(64136) <= 14785185;
srom_1(64137) <= 15141605;
srom_1(64138) <= 15466358;
srom_1(64139) <= 15757920;
srom_1(64140) <= 16014926;
srom_1(64141) <= 16236168;
srom_1(64142) <= 16420611;
srom_1(64143) <= 16567389;
srom_1(64144) <= 16675814;
srom_1(64145) <= 16745378;
srom_1(64146) <= 16775754;
srom_1(64147) <= 16766799;
srom_1(64148) <= 16718556;
srom_1(64149) <= 16631251;
srom_1(64150) <= 16505294;
srom_1(64151) <= 16341275;
srom_1(64152) <= 16139963;
srom_1(64153) <= 15902302;
srom_1(64154) <= 15629407;
srom_1(64155) <= 15322557;
srom_1(64156) <= 14983191;
srom_1(64157) <= 14612902;
srom_1(64158) <= 14213424;
srom_1(64159) <= 13786632;
srom_1(64160) <= 13334527;
srom_1(64161) <= 12859228;
srom_1(64162) <= 12362965;
srom_1(64163) <= 11848066;
srom_1(64164) <= 11316943;
srom_1(64165) <= 10772089;
srom_1(64166) <= 10216057;
srom_1(64167) <= 9651456;
srom_1(64168) <= 9080933;
srom_1(64169) <= 8507164;
srom_1(64170) <= 7932838;
srom_1(64171) <= 7360650;
srom_1(64172) <= 6793283;
srom_1(64173) <= 6233396;
srom_1(64174) <= 5683616;
srom_1(64175) <= 5146520;
srom_1(64176) <= 4624628;
srom_1(64177) <= 4120386;
srom_1(64178) <= 3636160;
srom_1(64179) <= 3174219;
srom_1(64180) <= 2736730;
srom_1(64181) <= 2325745;
srom_1(64182) <= 1943191;
srom_1(64183) <= 1590862;
srom_1(64184) <= 1270409;
srom_1(64185) <= 983336;
srom_1(64186) <= 730989;
srom_1(64187) <= 514552;
srom_1(64188) <= 335038;
srom_1(64189) <= 193290;
srom_1(64190) <= 89973;
srom_1(64191) <= 25572;
srom_1(64192) <= 387;
srom_1(64193) <= 14537;
srom_1(64194) <= 67957;
srom_1(64195) <= 160395;
srom_1(64196) <= 291417;
srom_1(64197) <= 460411;
srom_1(64198) <= 666582;
srom_1(64199) <= 908964;
srom_1(64200) <= 1186421;
srom_1(64201) <= 1497652;
srom_1(64202) <= 1841197;
srom_1(64203) <= 2215444;
srom_1(64204) <= 2618640;
srom_1(64205) <= 3048893;
srom_1(64206) <= 3504186;
srom_1(64207) <= 3982384;
srom_1(64208) <= 4481244;
srom_1(64209) <= 4998427;
srom_1(64210) <= 5531507;
srom_1(64211) <= 6077986;
srom_1(64212) <= 6635300;
srom_1(64213) <= 7200835;
srom_1(64214) <= 7771941;
srom_1(64215) <= 8345938;
srom_1(64216) <= 8920135;
srom_1(64217) <= 9491840;
srom_1(64218) <= 10058372;
srom_1(64219) <= 10617073;
srom_1(64220) <= 11165324;
srom_1(64221) <= 11700555;
srom_1(64222) <= 12220254;
srom_1(64223) <= 12721986;
srom_1(64224) <= 13203396;
srom_1(64225) <= 13662229;
srom_1(64226) <= 14096332;
srom_1(64227) <= 14503669;
srom_1(64228) <= 14882331;
srom_1(64229) <= 15230541;
srom_1(64230) <= 15546667;
srom_1(64231) <= 15829227;
srom_1(64232) <= 16076895;
srom_1(64233) <= 16288510;
srom_1(64234) <= 16463079;
srom_1(64235) <= 16599785;
srom_1(64236) <= 16697985;
srom_1(64237) <= 16757220;
srom_1(64238) <= 16777212;
srom_1(64239) <= 16757867;
srom_1(64240) <= 16699275;
srom_1(64241) <= 16601712;
srom_1(64242) <= 16465635;
srom_1(64243) <= 16291681;
srom_1(64244) <= 16080668;
srom_1(64245) <= 15833584;
srom_1(64246) <= 15551587;
srom_1(64247) <= 15236001;
srom_1(64248) <= 14888305;
srom_1(64249) <= 14510130;
srom_1(64250) <= 14103249;
srom_1(64251) <= 13669570;
srom_1(64252) <= 13211127;
srom_1(64253) <= 12730070;
srom_1(64254) <= 12228653;
srom_1(64255) <= 11709230;
srom_1(64256) <= 11174235;
srom_1(64257) <= 10626177;
srom_1(64258) <= 10067626;
srom_1(64259) <= 9501202;
srom_1(64260) <= 8929561;
srom_1(64261) <= 8355383;
srom_1(64262) <= 7781360;
srom_1(64263) <= 7210185;
srom_1(64264) <= 6644537;
srom_1(64265) <= 6087066;
srom_1(64266) <= 5540389;
srom_1(64267) <= 5007068;
srom_1(64268) <= 4489604;
srom_1(64269) <= 3990423;
srom_1(64270) <= 3511868;
srom_1(64271) <= 3056181;
srom_1(64272) <= 2625499;
srom_1(64273) <= 2221843;
srom_1(64274) <= 1847105;
srom_1(64275) <= 1503042;
srom_1(64276) <= 1191268;
srom_1(64277) <= 913245;
srom_1(64278) <= 670276;
srom_1(64279) <= 463501;
srom_1(64280) <= 293890;
srom_1(64281) <= 162238;
srom_1(64282) <= 69162;
srom_1(64283) <= 15098;
srom_1(64284) <= 301;
srom_1(64285) <= 24840;
srom_1(64286) <= 88599;
srom_1(64287) <= 191280;
srom_1(64288) <= 332401;
srom_1(64289) <= 511300;
srom_1(64290) <= 727138;
srom_1(64291) <= 978904;
srom_1(64292) <= 1265417;
srom_1(64293) <= 1585332;
srom_1(64294) <= 1937150;
srom_1(64295) <= 2319222;
srom_1(64296) <= 2729755;
srom_1(64297) <= 3166824;
srom_1(64298) <= 3628380;
srom_1(64299) <= 4112258;
srom_1(64300) <= 4616190;
srom_1(64301) <= 5137812;
srom_1(64302) <= 5674677;
srom_1(64303) <= 6224270;
srom_1(64304) <= 6784011;
srom_1(64305) <= 7351278;
srom_1(64306) <= 7923408;
srom_1(64307) <= 8497720;
srom_1(64308) <= 9071521;
srom_1(64309) <= 9642119;
srom_1(64310) <= 10206838;
srom_1(64311) <= 10763032;
srom_1(64312) <= 11308091;
srom_1(64313) <= 11839459;
srom_1(64314) <= 12354646;
srom_1(64315) <= 12851234;
srom_1(64316) <= 13326895;
srom_1(64317) <= 13779399;
srom_1(64318) <= 14206624;
srom_1(64319) <= 14606566;
srom_1(64320) <= 14977350;
srom_1(64321) <= 15317237;
srom_1(64322) <= 15624633;
srom_1(64323) <= 15898097;
srom_1(64324) <= 16136347;
srom_1(64325) <= 16338265;
srom_1(64326) <= 16502904;
srom_1(64327) <= 16629492;
srom_1(64328) <= 16717436;
srom_1(64329) <= 16766323;
srom_1(64330) <= 16775924;
srom_1(64331) <= 16746195;
srom_1(64332) <= 16677273;
srom_1(64333) <= 16569483;
srom_1(64334) <= 16423331;
srom_1(64335) <= 16239500;
srom_1(64336) <= 16018855;
srom_1(64337) <= 15762428;
srom_1(64338) <= 15471423;
srom_1(64339) <= 15147204;
srom_1(64340) <= 14791292;
srom_1(64341) <= 14405355;
srom_1(64342) <= 13991204;
srom_1(64343) <= 13550780;
srom_1(64344) <= 13086149;
srom_1(64345) <= 12599490;
srom_1(64346) <= 12093084;
srom_1(64347) <= 11569307;
srom_1(64348) <= 11030614;
srom_1(64349) <= 10479532;
srom_1(64350) <= 9918646;
srom_1(64351) <= 9350584;
srom_1(64352) <= 8778011;
srom_1(64353) <= 8203612;
srom_1(64354) <= 7630081;
srom_1(64355) <= 7060106;
srom_1(64356) <= 6496362;
srom_1(64357) <= 5941490;
srom_1(64358) <= 5398094;
srom_1(64359) <= 4868722;
srom_1(64360) <= 4355856;
srom_1(64361) <= 3861900;
srom_1(64362) <= 3389172;
srom_1(64363) <= 2939888;
srom_1(64364) <= 2516155;
srom_1(64365) <= 2119960;
srom_1(64366) <= 1753160;
srom_1(64367) <= 1417477;
srom_1(64368) <= 1114483;
srom_1(64369) <= 845601;
srom_1(64370) <= 612090;
srom_1(64371) <= 415046;
srom_1(64372) <= 255392;
srom_1(64373) <= 133879;
srom_1(64374) <= 51074;
srom_1(64375) <= 7367;
srom_1(64376) <= 2962;
srom_1(64377) <= 37881;
srom_1(64378) <= 111959;
srom_1(64379) <= 224849;
srom_1(64380) <= 376022;
srom_1(64381) <= 564768;
srom_1(64382) <= 790203;
srom_1(64383) <= 1051270;
srom_1(64384) <= 1346744;
srom_1(64385) <= 1675239;
srom_1(64386) <= 2035216;
srom_1(64387) <= 2424987;
srom_1(64388) <= 2842722;
srom_1(64389) <= 3286464;
srom_1(64390) <= 3754132;
srom_1(64391) <= 4243533;
srom_1(64392) <= 4752371;
srom_1(64393) <= 5278261;
srom_1(64394) <= 5818736;
srom_1(64395) <= 6371262;
srom_1(64396) <= 6933249;
srom_1(64397) <= 7502060;
srom_1(64398) <= 8075028;
srom_1(64399) <= 8649467;
srom_1(64400) <= 9222682;
srom_1(64401) <= 9791986;
srom_1(64402) <= 10354710;
srom_1(64403) <= 10908213;
srom_1(64404) <= 11449901;
srom_1(64405) <= 11977234;
srom_1(64406) <= 12487739;
srom_1(64407) <= 12979021;
srom_1(64408) <= 13448777;
srom_1(64409) <= 13894805;
srom_1(64410) <= 14315011;
srom_1(64411) <= 14707427;
srom_1(64412) <= 15070212;
srom_1(64413) <= 15401665;
srom_1(64414) <= 15700230;
srom_1(64415) <= 15964510;
srom_1(64416) <= 16193263;
srom_1(64417) <= 16385417;
srom_1(64418) <= 16540072;
srom_1(64419) <= 16656501;
srom_1(64420) <= 16734160;
srom_1(64421) <= 16772683;
srom_1(64422) <= 16771891;
srom_1(64423) <= 16731786;
srom_1(64424) <= 16652558;
srom_1(64425) <= 16534577;
srom_1(64426) <= 16378396;
srom_1(64427) <= 16184749;
srom_1(64428) <= 15954543;
srom_1(64429) <= 15688858;
srom_1(64430) <= 15388939;
srom_1(64431) <= 15056194;
srom_1(64432) <= 14692182;
srom_1(64433) <= 14298610;
srom_1(64434) <= 13877324;
srom_1(64435) <= 13430299;
srom_1(64436) <= 12959633;
srom_1(64437) <= 12467531;
srom_1(64438) <= 11956302;
srom_1(64439) <= 11428343;
srom_1(64440) <= 10886129;
srom_1(64441) <= 10332204;
srom_1(64442) <= 9769164;
srom_1(64443) <= 9199650;
srom_1(64444) <= 8626334;
srom_1(64445) <= 8051902;
srom_1(64446) <= 7479049;
srom_1(64447) <= 6910462;
srom_1(64448) <= 6348806;
srom_1(64449) <= 5796715;
srom_1(64450) <= 5256779;
srom_1(64451) <= 4731529;
srom_1(64452) <= 4223428;
srom_1(64453) <= 3734859;
srom_1(64454) <= 3268114;
srom_1(64455) <= 2825379;
srom_1(64456) <= 2408733;
srom_1(64457) <= 2020129;
srom_1(64458) <= 1661388;
srom_1(64459) <= 1334194;
srom_1(64460) <= 1040080;
srom_1(64461) <= 780426;
srom_1(64462) <= 556450;
srom_1(64463) <= 369201;
srom_1(64464) <= 219557;
srom_1(64465) <= 108222;
srom_1(64466) <= 35716;
srom_1(64467) <= 2379;
srom_1(64468) <= 8368;
srom_1(64469) <= 53656;
srom_1(64470) <= 138028;
srom_1(64471) <= 261091;
srom_1(64472) <= 422266;
srom_1(64473) <= 620798;
srom_1(64474) <= 855756;
srom_1(64475) <= 1126038;
srom_1(64476) <= 1430377;
srom_1(64477) <= 1767345;
srom_1(64478) <= 2135362;
srom_1(64479) <= 2532704;
srom_1(64480) <= 2957505;
srom_1(64481) <= 3407775;
srom_1(64482) <= 3881402;
srom_1(64483) <= 4376165;
srom_1(64484) <= 4889743;
srom_1(64485) <= 5419729;
srom_1(64486) <= 5963636;
srom_1(64487) <= 6518916;
srom_1(64488) <= 7082962;
srom_1(64489) <= 7653132;
srom_1(64490) <= 8226750;
srom_1(64491) <= 8801128;
srom_1(64492) <= 9373571;
srom_1(64493) <= 9941395;
srom_1(64494) <= 10501937;
srom_1(64495) <= 11052570;
srom_1(64496) <= 11590710;
srom_1(64497) <= 12113834;
srom_1(64498) <= 12619490;
srom_1(64499) <= 13105305;
srom_1(64500) <= 13569003;
srom_1(64501) <= 14008407;
srom_1(64502) <= 14421459;
srom_1(64503) <= 14806220;
srom_1(64504) <= 15160887;
srom_1(64505) <= 15483796;
srom_1(64506) <= 15773434;
srom_1(64507) <= 16028441;
srom_1(64508) <= 16247623;
srom_1(64509) <= 16429951;
srom_1(64510) <= 16574571;
srom_1(64511) <= 16680803;
srom_1(64512) <= 16748151;
srom_1(64513) <= 16776298;
srom_1(64514) <= 16765112;
srom_1(64515) <= 16714646;
srom_1(64516) <= 16625137;
srom_1(64517) <= 16497003;
srom_1(64518) <= 16330846;
srom_1(64519) <= 16127446;
srom_1(64520) <= 15887755;
srom_1(64521) <= 15612898;
srom_1(64522) <= 15304164;
srom_1(64523) <= 14963001;
srom_1(64524) <= 14591008;
srom_1(64525) <= 14189930;
srom_1(64526) <= 13761647;
srom_1(64527) <= 13308168;
srom_1(64528) <= 12831620;
srom_1(64529) <= 12334237;
srom_1(64530) <= 11818352;
srom_1(64531) <= 11286383;
srom_1(64532) <= 10740826;
srom_1(64533) <= 10184238;
srom_1(64534) <= 9619230;
srom_1(64535) <= 9048452;
srom_1(64536) <= 8474579;
srom_1(64537) <= 7900302;
srom_1(64538) <= 7328316;
srom_1(64539) <= 6761302;
srom_1(64540) <= 6201918;
srom_1(64541) <= 5652789;
srom_1(64542) <= 5116489;
srom_1(64543) <= 4595533;
srom_1(64544) <= 4092364;
srom_1(64545) <= 3609342;
srom_1(64546) <= 3148731;
srom_1(64547) <= 2712692;
srom_1(64548) <= 2303269;
srom_1(64549) <= 1922383;
srom_1(64550) <= 1571819;
srom_1(64551) <= 1253221;
srom_1(64552) <= 968083;
srom_1(64553) <= 717742;
srom_1(64554) <= 503373;
srom_1(64555) <= 325981;
srom_1(64556) <= 186397;
srom_1(64557) <= 85276;
srom_1(64558) <= 23092;
srom_1(64559) <= 137;
srom_1(64560) <= 16518;
srom_1(64561) <= 72159;
srom_1(64562) <= 166799;
srom_1(64563) <= 299993;
srom_1(64564) <= 471118;
srom_1(64565) <= 679371;
srom_1(64566) <= 923774;
srom_1(64567) <= 1203183;
srom_1(64568) <= 1516287;
srom_1(64569) <= 1861618;
srom_1(64570) <= 2237556;
srom_1(64571) <= 2642338;
srom_1(64572) <= 3074067;
srom_1(64573) <= 3530717;
srom_1(64574) <= 4010147;
srom_1(64575) <= 4510110;
srom_1(64576) <= 5028260;
srom_1(64577) <= 5562168;
srom_1(64578) <= 6109330;
srom_1(64579) <= 6667181;
srom_1(64580) <= 7233104;
srom_1(64581) <= 7804445;
srom_1(64582) <= 8378526;
srom_1(64583) <= 8952654;
srom_1(64584) <= 9524137;
srom_1(64585) <= 10090295;
srom_1(64586) <= 10648473;
srom_1(64587) <= 11196054;
srom_1(64588) <= 11730470;
srom_1(64589) <= 12249215;
srom_1(64590) <= 12749856;
srom_1(64591) <= 13230045;
srom_1(64592) <= 13687532;
srom_1(64593) <= 14120170;
srom_1(64594) <= 14525931;
srom_1(64595) <= 14902911;
srom_1(64596) <= 15249344;
srom_1(64597) <= 15563605;
srom_1(64598) <= 15844219;
srom_1(64599) <= 16089872;
srom_1(64600) <= 16299411;
srom_1(64601) <= 16471853;
srom_1(64602) <= 16606390;
srom_1(64603) <= 16702391;
srom_1(64604) <= 16759406;
srom_1(64605) <= 16777167;
srom_1(64606) <= 16755592;
srom_1(64607) <= 16694781;
srom_1(64608) <= 16595019;
srom_1(64609) <= 16456775;
srom_1(64610) <= 16280696;
srom_1(64611) <= 16067608;
srom_1(64612) <= 15818511;
srom_1(64613) <= 15534573;
srom_1(64614) <= 15217125;
srom_1(64615) <= 14867655;
srom_1(64616) <= 14487803;
srom_1(64617) <= 14079350;
srom_1(64618) <= 13644211;
srom_1(64619) <= 13184427;
srom_1(64620) <= 12702153;
srom_1(64621) <= 12199652;
srom_1(64622) <= 11679279;
srom_1(64623) <= 11143475;
srom_1(64624) <= 10594753;
srom_1(64625) <= 10035685;
srom_1(64626) <= 9468894;
srom_1(64627) <= 8897037;
srom_1(64628) <= 8322795;
srom_1(64629) <= 7748862;
srom_1(64630) <= 7177930;
srom_1(64631) <= 6612674;
srom_1(64632) <= 6055747;
srom_1(64633) <= 5509759;
srom_1(64634) <= 4977270;
srom_1(64635) <= 4460779;
srom_1(64636) <= 3962707;
srom_1(64637) <= 3485389;
srom_1(64638) <= 3031065;
srom_1(64639) <= 2601863;
srom_1(64640) <= 2199798;
srom_1(64641) <= 1826754;
srom_1(64642) <= 1484481;
srom_1(64643) <= 1174583;
srom_1(64644) <= 898515;
srom_1(64645) <= 657570;
srom_1(64646) <= 452879;
srom_1(64647) <= 285401;
srom_1(64648) <= 155922;
srom_1(64649) <= 65049;
srom_1(64650) <= 13207;
srom_1(64651) <= 641;
srom_1(64652) <= 27409;
srom_1(64653) <= 93386;
srom_1(64654) <= 198261;
srom_1(64655) <= 341544;
srom_1(64656) <= 522562;
srom_1(64657) <= 740467;
srom_1(64658) <= 994237;
srom_1(64659) <= 1282682;
srom_1(64660) <= 1604448;
srom_1(64661) <= 1958028;
srom_1(64662) <= 2341763;
srom_1(64663) <= 2753854;
srom_1(64664) <= 3192368;
srom_1(64665) <= 3655249;
srom_1(64666) <= 4140326;
srom_1(64667) <= 4645325;
srom_1(64668) <= 5167877;
srom_1(64669) <= 5705533;
srom_1(64670) <= 6255771;
srom_1(64671) <= 6816010;
srom_1(64672) <= 7383623;
srom_1(64673) <= 7955949;
srom_1(64674) <= 8530304;
srom_1(64675) <= 9103995;
srom_1(64676) <= 9674331;
srom_1(64677) <= 10238638;
srom_1(64678) <= 10794269;
srom_1(64679) <= 11338619;
srom_1(64680) <= 11869136;
srom_1(64681) <= 12383331;
srom_1(64682) <= 12878794;
srom_1(64683) <= 13353201;
srom_1(64684) <= 13804326;
srom_1(64685) <= 14230056;
srom_1(64686) <= 14628393;
srom_1(64687) <= 14997470;
srom_1(64688) <= 15335556;
srom_1(64689) <= 15641064;
srom_1(64690) <= 15912564;
srom_1(64691) <= 16148781;
srom_1(64692) <= 16348608;
srom_1(64693) <= 16511108;
srom_1(64694) <= 16635519;
srom_1(64695) <= 16721257;
srom_1(64696) <= 16767920;
srom_1(64697) <= 16775290;
srom_1(64698) <= 16743332;
srom_1(64699) <= 16672195;
srom_1(64700) <= 16562214;
srom_1(64701) <= 16413905;
srom_1(64702) <= 16227962;
srom_1(64703) <= 16005257;
srom_1(64704) <= 15746835;
srom_1(64705) <= 15453908;
srom_1(64706) <= 15127850;
srom_1(64707) <= 14770189;
srom_1(64708) <= 14382602;
srom_1(64709) <= 13966907;
srom_1(64710) <= 13525054;
srom_1(64711) <= 13059115;
srom_1(64712) <= 12571273;
srom_1(64713) <= 12063818;
srom_1(64714) <= 11539129;
srom_1(64715) <= 10999665;
srom_1(64716) <= 10447958;
srom_1(64717) <= 9886593;
srom_1(64718) <= 9318204;
srom_1(64719) <= 8745455;
srom_1(64720) <= 8171034;
srom_1(64721) <= 7597632;
srom_1(64722) <= 7027940;
srom_1(64723) <= 6464628;
srom_1(64724) <= 5910338;
srom_1(64725) <= 5367670;
srom_1(64726) <= 4839169;
srom_1(64727) <= 4327311;
srom_1(64728) <= 3834499;
srom_1(64729) <= 3363042;
srom_1(64730) <= 2915152;
srom_1(64731) <= 2492929;
srom_1(64732) <= 2098352;
srom_1(64733) <= 1733273;
srom_1(64734) <= 1399403;
srom_1(64735) <= 1098308;
srom_1(64736) <= 831399;
srom_1(64737) <= 599929;
srom_1(64738) <= 404982;
srom_1(64739) <= 247474;
srom_1(64740) <= 128142;
srom_1(64741) <= 47546;
srom_1(64742) <= 6065;
srom_1(64743) <= 3892;
srom_1(64744) <= 41037;
srom_1(64745) <= 117328;
srom_1(64746) <= 232405;
srom_1(64747) <= 385729;
srom_1(64748) <= 576582;
srom_1(64749) <= 804068;
srom_1(64750) <= 1067121;
srom_1(64751) <= 1364506;
srom_1(64752) <= 1694830;
srom_1(64753) <= 2056543;
srom_1(64754) <= 2447950;
srom_1(64755) <= 2867214;
srom_1(64756) <= 3312370;
srom_1(64757) <= 3781330;
srom_1(64758) <= 4271896;
srom_1(64759) <= 4781766;
srom_1(64760) <= 5308549;
srom_1(64761) <= 5849776;
srom_1(64762) <= 6402909;
srom_1(64763) <= 6965353;
srom_1(64764) <= 7534472;
srom_1(64765) <= 8107595;
srom_1(64766) <= 8682037;
srom_1(64767) <= 9255102;
srom_1(64768) <= 9824104;
srom_1(64769) <= 10386375;
srom_1(64770) <= 10939277;
srom_1(64771) <= 11480219;
srom_1(64772) <= 12006662;
srom_1(64773) <= 12516140;
srom_1(64774) <= 13006262;
srom_1(64775) <= 13474730;
srom_1(64776) <= 13919348;
srom_1(64777) <= 14338030;
srom_1(64778) <= 14728813;
srom_1(64779) <= 15089865;
srom_1(64780) <= 15419492;
srom_1(64781) <= 15716150;
srom_1(64782) <= 15978445;
srom_1(64783) <= 16205150;
srom_1(64784) <= 16395200;
srom_1(64785) <= 16547704;
srom_1(64786) <= 16661947;
srom_1(64787) <= 16737394;
srom_1(64788) <= 16773691;
srom_1(64789) <= 16770667;
srom_1(64790) <= 16728336;
srom_1(64791) <= 16646898;
srom_1(64792) <= 16526734;
srom_1(64793) <= 16368407;
srom_1(64794) <= 16172661;
srom_1(64795) <= 15940412;
srom_1(64796) <= 15672750;
srom_1(64797) <= 15370931;
srom_1(64798) <= 15036368;
srom_1(64799) <= 14670633;
srom_1(64800) <= 14275438;
srom_1(64801) <= 13852639;
srom_1(64802) <= 13404216;
srom_1(64803) <= 12932274;
srom_1(64804) <= 12439025;
srom_1(64805) <= 11926782;
srom_1(64806) <= 11397947;
srom_1(64807) <= 10855000;
srom_1(64808) <= 10300488;
srom_1(64809) <= 9737010;
srom_1(64810) <= 9167209;
srom_1(64811) <= 8593757;
srom_1(64812) <= 8019343;
srom_1(64813) <= 7446661;
srom_1(64814) <= 6878395;
srom_1(64815) <= 6317212;
srom_1(64816) <= 5765742;
srom_1(64817) <= 5226571;
srom_1(64818) <= 4702229;
srom_1(64819) <= 4195173;
srom_1(64820) <= 3707781;
srom_1(64821) <= 3242340;
srom_1(64822) <= 2801031;
srom_1(64823) <= 2385924;
srom_1(64824) <= 1998966;
srom_1(64825) <= 1641971;
srom_1(64826) <= 1316614;
srom_1(64827) <= 1024419;
srom_1(64828) <= 766758;
srom_1(64829) <= 544838;
srom_1(64830) <= 359700;
srom_1(64831) <= 212212;
srom_1(64832) <= 103067;
srom_1(64833) <= 32775;
srom_1(64834) <= 1666;
srom_1(64835) <= 9887;
srom_1(64836) <= 57398;
srom_1(64837) <= 143978;
srom_1(64838) <= 269219;
srom_1(64839) <= 432535;
srom_1(64840) <= 633159;
srom_1(64841) <= 870152;
srom_1(64842) <= 1142401;
srom_1(64843) <= 1448630;
srom_1(64844) <= 1787403;
srom_1(64845) <= 2157132;
srom_1(64846) <= 2556081;
srom_1(64847) <= 2982382;
srom_1(64848) <= 3434034;
srom_1(64849) <= 3908920;
srom_1(64850) <= 4404813;
srom_1(64851) <= 4919387;
srom_1(64852) <= 5450229;
srom_1(64853) <= 5994851;
srom_1(64854) <= 6550698;
srom_1(64855) <= 7115163;
srom_1(64856) <= 7685600;
srom_1(64857) <= 8259333;
srom_1(64858) <= 8833673;
srom_1(64859) <= 9405926;
srom_1(64860) <= 9973408;
srom_1(64861) <= 10533458;
srom_1(64862) <= 11083450;
srom_1(64863) <= 11620806;
srom_1(64864) <= 12143004;
srom_1(64865) <= 12647597;
srom_1(64866) <= 13132218;
srom_1(64867) <= 13594595;
srom_1(64868) <= 14032559;
srom_1(64869) <= 14444056;
srom_1(64870) <= 14827157;
srom_1(64871) <= 15180066;
srom_1(64872) <= 15501128;
srom_1(64873) <= 15788836;
srom_1(64874) <= 16041842;
srom_1(64875) <= 16258959;
srom_1(64876) <= 16439170;
srom_1(64877) <= 16581629;
srom_1(64878) <= 16685667;
srom_1(64879) <= 16750798;
srom_1(64880) <= 16776716;
srom_1(64881) <= 16763299;
srom_1(64882) <= 16710611;
srom_1(64883) <= 16618897;
srom_1(64884) <= 16488589;
srom_1(64885) <= 16320298;
srom_1(64886) <= 16114812;
srom_1(64887) <= 15873095;
srom_1(64888) <= 15596280;
srom_1(64889) <= 15285667;
srom_1(64890) <= 14942711;
srom_1(64891) <= 14569020;
srom_1(64892) <= 14166347;
srom_1(64893) <= 13736581;
srom_1(64894) <= 13281736;
srom_1(64895) <= 12803945;
srom_1(64896) <= 12305450;
srom_1(64897) <= 11788586;
srom_1(64898) <= 11255780;
srom_1(64899) <= 10709528;
srom_1(64900) <= 10152392;
srom_1(64901) <= 9586986;
srom_1(64902) <= 9015960;
srom_1(64903) <= 8441992;
srom_1(64904) <= 7867774;
srom_1(64905) <= 7295998;
srom_1(64906) <= 6729345;
srom_1(64907) <= 6170474;
srom_1(64908) <= 5622004;
srom_1(64909) <= 5086507;
srom_1(64910) <= 4566496;
srom_1(64911) <= 4064407;
srom_1(64912) <= 3582597;
srom_1(64913) <= 3123323;
srom_1(64914) <= 2688740;
srom_1(64915) <= 2280885;
srom_1(64916) <= 1901672;
srom_1(64917) <= 1552878;
srom_1(64918) <= 1236140;
srom_1(64919) <= 952941;
srom_1(64920) <= 704611;
srom_1(64921) <= 492314;
srom_1(64922) <= 317046;
srom_1(64923) <= 179627;
srom_1(64924) <= 80704;
srom_1(64925) <= 20739;
srom_1(64926) <= 14;
srom_1(64927) <= 18626;
srom_1(64928) <= 76487;
srom_1(64929) <= 173327;
srom_1(64930) <= 308691;
srom_1(64931) <= 481945;
srom_1(64932) <= 692276;
srom_1(64933) <= 938697;
srom_1(64934) <= 1220054;
srom_1(64935) <= 1535026;
srom_1(64936) <= 1882138;
srom_1(64937) <= 2259760;
srom_1(64938) <= 2666123;
srom_1(64939) <= 3099320;
srom_1(64940) <= 3557321;
srom_1(64941) <= 4037977;
srom_1(64942) <= 4539035;
srom_1(64943) <= 5058144;
srom_1(64944) <= 5592872;
srom_1(64945) <= 6140709;
srom_1(64946) <= 6699088;
srom_1(64947) <= 7265389;
srom_1(64948) <= 7836958;
srom_1(64949) <= 8411114;
srom_1(64950) <= 8985163;
srom_1(64951) <= 9556416;
srom_1(64952) <= 10122192;
srom_1(64953) <= 10679839;
srom_1(64954) <= 11226741;
srom_1(64955) <= 11760335;
srom_1(64956) <= 12278117;
srom_1(64957) <= 12777660;
srom_1(64958) <= 13256621;
srom_1(64959) <= 13712755;
srom_1(64960) <= 14143922;
srom_1(64961) <= 14548100;
srom_1(64962) <= 14923394;
srom_1(64963) <= 15268044;
srom_1(64964) <= 15580434;
srom_1(64965) <= 15859099;
srom_1(64966) <= 16102733;
srom_1(64967) <= 16310192;
srom_1(64968) <= 16480504;
srom_1(64969) <= 16612871;
srom_1(64970) <= 16706671;
srom_1(64971) <= 16761465;
srom_1(64972) <= 16776996;
srom_1(64973) <= 16753190;
srom_1(64974) <= 16690161;
srom_1(64975) <= 16588202;
srom_1(64976) <= 16447793;
srom_1(64977) <= 16269591;
srom_1(64978) <= 16054433;
srom_1(64979) <= 15803327;
srom_1(64980) <= 15517451;
srom_1(64981) <= 15198145;
srom_1(64982) <= 14846907;
srom_1(64983) <= 14465384;
srom_1(64984) <= 14055365;
srom_1(64985) <= 13618772;
srom_1(64986) <= 13157653;
srom_1(64987) <= 12674171;
srom_1(64988) <= 12170592;
srom_1(64989) <= 11649278;
srom_1(64990) <= 11112674;
srom_1(64991) <= 10563296;
srom_1(64992) <= 10003719;
srom_1(64993) <= 9436569;
srom_1(64994) <= 8864505;
srom_1(64995) <= 8290209;
srom_1(64996) <= 7716374;
srom_1(64997) <= 7145692;
srom_1(64998) <= 6580838;
srom_1(64999) <= 6024462;
srom_1(65000) <= 5479172;
srom_1(65001) <= 4947525;
srom_1(65002) <= 4432014;
srom_1(65003) <= 3935058;
srom_1(65004) <= 3458985;
srom_1(65005) <= 3006029;
srom_1(65006) <= 2578314;
srom_1(65007) <= 2177846;
srom_1(65008) <= 1806502;
srom_1(65009) <= 1466023;
srom_1(65010) <= 1158007;
srom_1(65011) <= 883898;
srom_1(65012) <= 644981;
srom_1(65013) <= 442376;
srom_1(65014) <= 277034;
srom_1(65015) <= 149730;
srom_1(65016) <= 61061;
srom_1(65017) <= 11443;
srom_1(65018) <= 1108;
srom_1(65019) <= 30104;
srom_1(65020) <= 98297;
srom_1(65021) <= 205366;
srom_1(65022) <= 350809;
srom_1(65023) <= 533944;
srom_1(65024) <= 753912;
srom_1(65025) <= 1009682;
srom_1(65026) <= 1300054;
srom_1(65027) <= 1623667;
srom_1(65028) <= 1979002;
srom_1(65029) <= 2364395;
srom_1(65030) <= 2778038;
srom_1(65031) <= 3217990;
srom_1(65032) <= 3682189;
srom_1(65033) <= 4168458;
srom_1(65034) <= 4674517;
srom_1(65035) <= 5197992;
srom_1(65036) <= 5736429;
srom_1(65037) <= 6287303;
srom_1(65038) <= 6848031;
srom_1(65039) <= 7415984;
srom_1(65040) <= 7988497;
srom_1(65041) <= 8562886;
srom_1(65042) <= 9136459;
srom_1(65043) <= 9706524;
srom_1(65044) <= 10270409;
srom_1(65045) <= 10825470;
srom_1(65046) <= 11369103;
srom_1(65047) <= 11898760;
srom_1(65048) <= 12411957;
srom_1(65049) <= 12906286;
srom_1(65050) <= 13379431;
srom_1(65051) <= 13829172;
srom_1(65052) <= 14253400;
srom_1(65053) <= 14650127;
srom_1(65054) <= 15017490;
srom_1(65055) <= 15353769;
srom_1(65056) <= 15657386;
srom_1(65057) <= 15926917;
srom_1(65058) <= 16161098;
srom_1(65059) <= 16358831;
srom_1(65060) <= 16519190;
srom_1(65061) <= 16641421;
srom_1(65062) <= 16724951;
srom_1(65063) <= 16769390;
srom_1(65064) <= 16774529;
srom_1(65065) <= 16740343;
srom_1(65066) <= 16666993;
srom_1(65067) <= 16554822;
srom_1(65068) <= 16404358;
srom_1(65069) <= 16216304;
srom_1(65070) <= 15991544;
srom_1(65071) <= 15731132;
srom_1(65072) <= 15436287;
srom_1(65073) <= 15108394;
srom_1(65074) <= 14748989;
srom_1(65075) <= 14359759;
srom_1(65076) <= 13942527;
srom_1(65077) <= 13499251;
srom_1(65078) <= 13032010;
srom_1(65079) <= 12542994;
srom_1(65080) <= 12034497;
srom_1(65081) <= 11508903;
srom_1(65082) <= 10968676;
srom_1(65083) <= 10416351;
srom_1(65084) <= 9854518;
srom_1(65085) <= 9285810;
srom_1(65086) <= 8712894;
srom_1(65087) <= 8138458;
srom_1(65088) <= 7565195;
srom_1(65089) <= 6995794;
srom_1(65090) <= 6432923;
srom_1(65091) <= 5879224;
srom_1(65092) <= 5337292;
srom_1(65093) <= 4809669;
srom_1(65094) <= 4298828;
srom_1(65095) <= 3807166;
srom_1(65096) <= 3336988;
srom_1(65097) <= 2890498;
srom_1(65098) <= 2469791;
srom_1(65099) <= 2076840;
srom_1(65100) <= 1713486;
srom_1(65101) <= 1381435;
srom_1(65102) <= 1082242;
srom_1(65103) <= 817311;
srom_1(65104) <= 587885;
srom_1(65105) <= 395040;
srom_1(65106) <= 239678;
srom_1(65107) <= 122530;
srom_1(65108) <= 44144;
srom_1(65109) <= 4889;
srom_1(65110) <= 4947;
srom_1(65111) <= 44320;
srom_1(65112) <= 122821;
srom_1(65113) <= 240084;
srom_1(65114) <= 395558;
srom_1(65115) <= 588514;
srom_1(65116) <= 818047;
srom_1(65117) <= 1083082;
srom_1(65118) <= 1382374;
srom_1(65119) <= 1714521;
srom_1(65120) <= 2077966;
srom_1(65121) <= 2471003;
srom_1(65122) <= 2891789;
srom_1(65123) <= 3338352;
srom_1(65124) <= 3808598;
srom_1(65125) <= 4300320;
srom_1(65126) <= 4811214;
srom_1(65127) <= 5338884;
srom_1(65128) <= 5880855;
srom_1(65129) <= 6434586;
srom_1(65130) <= 6997479;
srom_1(65131) <= 7566896;
srom_1(65132) <= 8140167;
srom_1(65133) <= 8714602;
srom_1(65134) <= 9287509;
srom_1(65135) <= 9856200;
srom_1(65136) <= 10418010;
srom_1(65137) <= 10970303;
srom_1(65138) <= 11510489;
srom_1(65139) <= 12036036;
srom_1(65140) <= 12544479;
srom_1(65141) <= 13033433;
srom_1(65142) <= 13500606;
srom_1(65143) <= 13943808;
srom_1(65144) <= 14360959;
srom_1(65145) <= 14750104;
srom_1(65146) <= 15109417;
srom_1(65147) <= 15437214;
srom_1(65148) <= 15731958;
srom_1(65149) <= 15992267;
srom_1(65150) <= 16216919;
srom_1(65151) <= 16404861;
srom_1(65152) <= 16555213;
srom_1(65153) <= 16667269;
srom_1(65154) <= 16740503;
srom_1(65155) <= 16774572;
srom_1(65156) <= 16769316;
srom_1(65157) <= 16724761;
srom_1(65158) <= 16641114;
srom_1(65159) <= 16518769;
srom_1(65160) <= 16358298;
srom_1(65161) <= 16160455;
srom_1(65162) <= 15926167;
srom_1(65163) <= 15656533;
srom_1(65164) <= 15352817;
srom_1(65165) <= 15016443;
srom_1(65166) <= 14648989;
srom_1(65167) <= 14252178;
srom_1(65168) <= 13827871;
srom_1(65169) <= 13378057;
srom_1(65170) <= 12904846;
srom_1(65171) <= 12410457;
srom_1(65172) <= 11897208;
srom_1(65173) <= 11367505;
srom_1(65174) <= 10823834;
srom_1(65175) <= 10268743;
srom_1(65176) <= 9704836;
srom_1(65177) <= 9134756;
srom_1(65178) <= 8561178;
srom_1(65179) <= 7986790;
srom_1(65180) <= 7414286;
srom_1(65181) <= 6846351;
srom_1(65182) <= 6285649;
srom_1(65183) <= 5734808;
srom_1(65184) <= 5196411;
srom_1(65185) <= 4672984;
srom_1(65186) <= 4166981;
srom_1(65187) <= 3680774;
srom_1(65188) <= 3216644;
srom_1(65189) <= 2776767;
srom_1(65190) <= 2363206;
srom_1(65191) <= 1977900;
srom_1(65192) <= 1622656;
srom_1(65193) <= 1299140;
srom_1(65194) <= 1008869;
srom_1(65195) <= 753204;
srom_1(65196) <= 533344;
srom_1(65197) <= 350320;
srom_1(65198) <= 204990;
srom_1(65199) <= 98036;
srom_1(65200) <= 29960;
srom_1(65201) <= 1080;
srom_1(65202) <= 11532;
srom_1(65203) <= 61267;
srom_1(65204) <= 150052;
srom_1(65205) <= 277470;
srom_1(65206) <= 442924;
srom_1(65207) <= 645638;
srom_1(65208) <= 884662;
srom_1(65209) <= 1158874;
srom_1(65210) <= 1466989;
srom_1(65211) <= 1807561;
srom_1(65212) <= 2178995;
srom_1(65213) <= 2579547;
srom_1(65214) <= 3007340;
srom_1(65215) <= 3460368;
srom_1(65216) <= 3936506;
srom_1(65217) <= 4433521;
srom_1(65218) <= 4949084;
srom_1(65219) <= 5480775;
srom_1(65220) <= 6026102;
srom_1(65221) <= 6582507;
srom_1(65222) <= 7147383;
srom_1(65223) <= 7718078;
srom_1(65224) <= 8291918;
srom_1(65225) <= 8866211;
srom_1(65226) <= 9438265;
srom_1(65227) <= 10005397;
srom_1(65228) <= 10564946;
srom_1(65229) <= 11114291;
srom_1(65230) <= 11650853;
srom_1(65231) <= 12172118;
srom_1(65232) <= 12675640;
srom_1(65233) <= 13159059;
srom_1(65234) <= 13620108;
srom_1(65235) <= 14056625;
srom_1(65236) <= 14466562;
srom_1(65237) <= 14847998;
srom_1(65238) <= 15199143;
srom_1(65239) <= 15518352;
srom_1(65240) <= 15804126;
srom_1(65241) <= 16055127;
srom_1(65242) <= 16270177;
srom_1(65243) <= 16448267;
srom_1(65244) <= 16588563;
srom_1(65245) <= 16690406;
srom_1(65246) <= 16753319;
srom_1(65247) <= 16777008;
srom_1(65248) <= 16761360;
srom_1(65249) <= 16706450;
srom_1(65250) <= 16612534;
srom_1(65251) <= 16480054;
srom_1(65252) <= 16309630;
srom_1(65253) <= 16102061;
srom_1(65254) <= 15858322;
srom_1(65255) <= 15579554;
srom_1(65256) <= 15267066;
srom_1(65257) <= 14922322;
srom_1(65258) <= 14546939;
srom_1(65259) <= 14142678;
srom_1(65260) <= 13711434;
srom_1(65261) <= 13255229;
srom_1(65262) <= 12776204;
srom_1(65263) <= 12276603;
srom_1(65264) <= 11758770;
srom_1(65265) <= 11225133;
srom_1(65266) <= 10678195;
srom_1(65267) <= 10120520;
srom_1(65268) <= 9554723;
srom_1(65269) <= 8983459;
srom_1(65270) <= 8409404;
srom_1(65271) <= 7835253;
srom_1(65272) <= 7263696;
srom_1(65273) <= 6697414;
srom_1(65274) <= 6139063;
srom_1(65275) <= 5591260;
srom_1(65276) <= 5056576;
srom_1(65277) <= 4537516;
srom_1(65278) <= 4036516;
srom_1(65279) <= 3555924;
srom_1(65280) <= 3097994;
srom_1(65281) <= 2664873;
srom_1(65282) <= 2258593;
srom_1(65283) <= 1881059;
srom_1(65284) <= 1534041;
srom_1(65285) <= 1219166;
srom_1(65286) <= 937912;
srom_1(65287) <= 691596;
srom_1(65288) <= 481374;
srom_1(65289) <= 308232;
srom_1(65290) <= 172982;
srom_1(65291) <= 76257;
srom_1(65292) <= 18512;
srom_1(65293) <= 17;
srom_1(65294) <= 20859;
srom_1(65295) <= 80940;
srom_1(65296) <= 179979;
srom_1(65297) <= 317511;
srom_1(65298) <= 492891;
srom_1(65299) <= 705297;
srom_1(65300) <= 953733;
srom_1(65301) <= 1237033;
srom_1(65302) <= 1553869;
srom_1(65303) <= 1902756;
srom_1(65304) <= 2282057;
srom_1(65305) <= 2689994;
srom_1(65306) <= 3124653;
srom_1(65307) <= 3583997;
srom_1(65308) <= 4065872;
srom_1(65309) <= 4568017;
srom_1(65310) <= 5088079;
srom_1(65311) <= 5623617;
srom_1(65312) <= 6172122;
srom_1(65313) <= 6731021;
srom_1(65314) <= 7297692;
srom_1(65315) <= 7869479;
srom_1(65316) <= 8443701;
srom_1(65317) <= 9017664;
srom_1(65318) <= 9588678;
srom_1(65319) <= 10154063;
srom_1(65320) <= 10711170;
srom_1(65321) <= 11257386;
srom_1(65322) <= 11790149;
srom_1(65323) <= 12306961;
srom_1(65324) <= 12805398;
srom_1(65325) <= 13283124;
srom_1(65326) <= 13737897;
srom_1(65327) <= 14167586;
srom_1(65328) <= 14570176;
srom_1(65329) <= 14943777;
srom_1(65330) <= 15286640;
srom_1(65331) <= 15597155;
srom_1(65332) <= 15873866;
srom_1(65333) <= 16115477;
srom_1(65334) <= 16320854;
srom_1(65335) <= 16489034;
srom_1(65336) <= 16619228;
srom_1(65337) <= 16710826;
srom_1(65338) <= 16763398;
srom_1(65339) <= 16776698;
srom_1(65340) <= 16750663;
srom_1(65341) <= 16685415;
srom_1(65342) <= 16581261;
srom_1(65343) <= 16438689;
srom_1(65344) <= 16258368;
srom_1(65345) <= 16041142;
srom_1(65346) <= 15788031;
srom_1(65347) <= 15500221;
srom_1(65348) <= 15179063;
srom_1(65349) <= 14826062;
srom_1(65350) <= 14442873;
srom_1(65351) <= 14031294;
srom_1(65352) <= 13593254;
srom_1(65353) <= 13130808;
srom_1(65354) <= 12646125;
srom_1(65355) <= 12141476;
srom_1(65356) <= 11619229;
srom_1(65357) <= 11081832;
srom_1(65358) <= 10531806;
srom_1(65359) <= 9971729;
srom_1(65360) <= 9404229;
srom_1(65361) <= 8831966;
srom_1(65362) <= 8257624;
srom_1(65363) <= 7683897;
srom_1(65364) <= 7113474;
srom_1(65365) <= 6549030;
srom_1(65366) <= 5993213;
srom_1(65367) <= 5448629;
srom_1(65368) <= 4917831;
srom_1(65369) <= 4403309;
srom_1(65370) <= 3907475;
srom_1(65371) <= 3432655;
srom_1(65372) <= 2981075;
srom_1(65373) <= 2554853;
srom_1(65374) <= 2155988;
srom_1(65375) <= 1786349;
srom_1(65376) <= 1447670;
srom_1(65377) <= 1141540;
srom_1(65378) <= 869394;
srom_1(65379) <= 632508;
srom_1(65380) <= 431993;
srom_1(65381) <= 268790;
srom_1(65382) <= 143663;
srom_1(65383) <= 57199;
srom_1(65384) <= 9804;
srom_1(65385) <= 1700;
srom_1(65386) <= 32926;
srom_1(65387) <= 103334;
srom_1(65388) <= 212594;
srom_1(65389) <= 360195;
srom_1(65390) <= 545444;
srom_1(65391) <= 767472;
srom_1(65392) <= 1025238;
srom_1(65393) <= 1317533;
srom_1(65394) <= 1642987;
srom_1(65395) <= 2000074;
srom_1(65396) <= 2387118;
srom_1(65397) <= 2802306;
srom_1(65398) <= 3243690;
srom_1(65399) <= 3709200;
srom_1(65400) <= 4196653;
srom_1(65401) <= 4703764;
srom_1(65402) <= 5228155;
srom_1(65403) <= 5767365;
srom_1(65404) <= 6318868;
srom_1(65405) <= 6880077;
srom_1(65406) <= 7448359;
srom_1(65407) <= 8021051;
srom_1(65408) <= 8595466;
srom_1(65409) <= 9168911;
srom_1(65410) <= 9738697;
srom_1(65411) <= 10302152;
srom_1(65412) <= 10856634;
srom_1(65413) <= 11399542;
srom_1(65414) <= 11928331;
srom_1(65415) <= 12440521;
srom_1(65416) <= 12933710;
srom_1(65417) <= 13405586;
srom_1(65418) <= 13853935;
srom_1(65419) <= 14276656;
srom_1(65420) <= 14671765;
srom_1(65421) <= 15037411;
srom_1(65422) <= 15371878;
srom_1(65423) <= 15673598;
srom_1(65424) <= 15941156;
srom_1(65425) <= 16173298;
srom_1(65426) <= 16368934;
srom_1(65427) <= 16527148;
srom_1(65428) <= 16647198;
srom_1(65429) <= 16728521;
srom_1(65430) <= 16770734;
srom_1(65431) <= 16773641;
srom_1(65432) <= 16737228;
srom_1(65433) <= 16661665;
srom_1(65434) <= 16547307;
srom_1(65435) <= 16394690;
srom_1(65436) <= 16204529;
srom_1(65437) <= 15977717;
srom_1(65438) <= 15715317;
srom_1(65439) <= 15418560;
srom_1(65440) <= 15088837;
srom_1(65441) <= 14727694;
srom_1(65442) <= 14336825;
srom_1(65443) <= 13918063;
srom_1(65444) <= 13473371;
srom_1(65445) <= 13004835;
srom_1(65446) <= 12514652;
srom_1(65447) <= 12005120;
srom_1(65448) <= 11478630;
srom_1(65449) <= 10937649;
srom_1(65450) <= 10384715;
srom_1(65451) <= 9822420;
srom_1(65452) <= 9253402;
srom_1(65453) <= 8680329;
srom_1(65454) <= 8105887;
srom_1(65455) <= 7532771;
srom_1(65456) <= 6963669;
srom_1(65457) <= 6401248;
srom_1(65458) <= 5848147;
srom_1(65459) <= 5306960;
srom_1(65460) <= 4780223;
srom_1(65461) <= 4270406;
srom_1(65462) <= 3779902;
srom_1(65463) <= 3311009;
srom_1(65464) <= 2865927;
srom_1(65465) <= 2446743;
srom_1(65466) <= 2055422;
srom_1(65467) <= 1693800;
srom_1(65468) <= 1363572;
srom_1(65469) <= 1066287;
srom_1(65470) <= 803338;
srom_1(65471) <= 575960;
srom_1(65472) <= 385217;
srom_1(65473) <= 232006;
srom_1(65474) <= 117043;
srom_1(65475) <= 40869;
srom_1(65476) <= 3840;
srom_1(65477) <= 6130;
srom_1(65478) <= 47728;
srom_1(65479) <= 128440;
srom_1(65480) <= 247886;
srom_1(65481) <= 405507;
srom_1(65482) <= 600564;
srom_1(65483) <= 832141;
srom_1(65484) <= 1099153;
srom_1(65485) <= 1400348;
srom_1(65486) <= 1734314;
srom_1(65487) <= 2099483;
srom_1(65488) <= 2494145;
srom_1(65489) <= 2916447;
srom_1(65490) <= 3364411;
srom_1(65491) <= 3835934;
srom_1(65492) <= 4328807;
srom_1(65493) <= 4840717;
srom_1(65494) <= 5369265;
srom_1(65495) <= 5911971;
srom_1(65496) <= 6466292;
srom_1(65497) <= 7029626;
srom_1(65498) <= 7599334;
srom_1(65499) <= 8172742;
srom_1(65500) <= 8747163;
srom_1(65501) <= 9319902;
srom_1(65502) <= 9888275;
srom_1(65503) <= 10449614;
srom_1(65504) <= 11001289;
srom_1(65505) <= 11540713;
srom_1(65506) <= 12065354;
srom_1(65507) <= 12572755;
srom_1(65508) <= 13060534;
srom_1(65509) <= 13526406;
srom_1(65510) <= 13968184;
srom_1(65511) <= 14383798;
srom_1(65512) <= 14771298;
srom_1(65513) <= 15128867;
srom_1(65514) <= 15454830;
srom_1(65515) <= 15747656;
srom_1(65516) <= 16005973;
srom_1(65517) <= 16228570;
srom_1(65518) <= 16414402;
srom_1(65519) <= 16562599;
srom_1(65520) <= 16672465;
srom_1(65521) <= 16743485;
srom_1(65522) <= 16775326;
srom_1(65523) <= 16767839;
srom_1(65524) <= 16721059;
srom_1(65525) <= 16635206;
srom_1(65526) <= 16510681;
srom_1(65527) <= 16348069;
srom_1(65528) <= 16148132;
srom_1(65529) <= 15911808;
srom_1(65530) <= 15640205;
srom_1(65531) <= 15334597;
srom_1(65532) <= 14996417;
srom_1(65533) <= 14627251;
srom_1(65534) <= 14228829;
srom_1(65535) <= 13803021;
srom_1(65536) <= 13351823;
srom_1(65537) <= 12877350;
srom_1(65538) <= 12381828;
srom_1(65539) <= 11867581;
srom_1(65540) <= 11337019;
srom_1(65541) <= 10792632;
srom_1(65542) <= 10236971;
srom_1(65543) <= 9672642;
srom_1(65544) <= 9102292;
srom_1(65545) <= 8528595;
srom_1(65546) <= 7954242;
srom_1(65547) <= 7381926;
srom_1(65548) <= 6814331;
srom_1(65549) <= 6254118;
srom_1(65550) <= 5703914;
srom_1(65551) <= 5166299;
srom_1(65552) <= 4643795;
srom_1(65553) <= 4138852;
srom_1(65554) <= 3653838;
srom_1(65555) <= 3191026;
srom_1(65556) <= 2752588;
srom_1(65557) <= 2340578;
srom_1(65558) <= 1956931;
srom_1(65559) <= 1603443;
srom_1(65560) <= 1281773;
srom_1(65561) <= 993430;
srom_1(65562) <= 739765;
srom_1(65563) <= 521969;
srom_1(65564) <= 341061;
srom_1(65565) <= 197892;
srom_1(65566) <= 93131;
srom_1(65567) <= 27271;
srom_1(65568) <= 620;
srom_1(65569) <= 13303;
srom_1(65570) <= 65261;
srom_1(65571) <= 156250;
srom_1(65572) <= 285843;
srom_1(65573) <= 453433;
srom_1(65574) <= 658234;
srom_1(65575) <= 899285;
srom_1(65576) <= 1175456;
srom_1(65577) <= 1485451;
srom_1(65578) <= 1827819;
srom_1(65579) <= 2200952;
srom_1(65580) <= 2603101;
srom_1(65581) <= 3032380;
srom_1(65582) <= 3486776;
srom_1(65583) <= 3964159;
srom_1(65584) <= 4462290;
srom_1(65585) <= 4978832;
srom_1(65586) <= 5511364;
srom_1(65587) <= 6057388;
srom_1(65588) <= 6614345;
srom_1(65589) <= 7179621;
srom_1(65590) <= 7750567;
srom_1(65591) <= 8324504;
srom_1(65592) <= 8898743;
srom_1(65593) <= 9470589;
srom_1(65594) <= 10037361;
srom_1(65595) <= 10596402;
srom_1(65596) <= 11145089;
srom_1(65597) <= 11680851;
srom_1(65598) <= 12201174;
srom_1(65599) <= 12703619;
srom_1(65600) <= 13185829;
srom_1(65601) <= 13645543;
srom_1(65602) <= 14080606;
srom_1(65603) <= 14488977;
srom_1(65604) <= 14868741;
srom_1(65605) <= 15218117;
srom_1(65606) <= 15535468;
srom_1(65607) <= 15819305;
srom_1(65608) <= 16068296;
srom_1(65609) <= 16281275;
srom_1(65610) <= 16457242;
srom_1(65611) <= 16595373;
srom_1(65612) <= 16695019;
srom_1(65613) <= 16755714;
srom_1(65614) <= 16777173;
srom_1(65615) <= 16759294;
srom_1(65616) <= 16702163;
srom_1(65617) <= 16606047;
srom_1(65618) <= 16471396;
srom_1(65619) <= 16298842;
srom_1(65620) <= 16089194;
srom_1(65621) <= 15843436;
srom_1(65622) <= 15562719;
srom_1(65623) <= 15248361;
srom_1(65624) <= 14901834;
srom_1(65625) <= 14524765;
srom_1(65626) <= 14118922;
srom_1(65627) <= 13686207;
srom_1(65628) <= 13228650;
srom_1(65629) <= 12748396;
srom_1(65630) <= 12247697;
srom_1(65631) <= 11728902;
srom_1(65632) <= 11194443;
srom_1(65633) <= 10646827;
srom_1(65634) <= 10088621;
srom_1(65635) <= 9522443;
srom_1(65636) <= 8950948;
srom_1(65637) <= 8376817;
srom_1(65638) <= 7802740;
srom_1(65639) <= 7231411;
srom_1(65640) <= 6665508;
srom_1(65641) <= 6107685;
srom_1(65642) <= 5560559;
srom_1(65643) <= 5026694;
srom_1(65644) <= 4508594;
srom_1(65645) <= 4008689;
srom_1(65646) <= 3529323;
srom_1(65647) <= 3072744;
srom_1(65648) <= 2641093;
srom_1(65649) <= 2236394;
srom_1(65650) <= 1860544;
srom_1(65651) <= 1515307;
srom_1(65652) <= 1202302;
srom_1(65653) <= 922995;
srom_1(65654) <= 678697;
srom_1(65655) <= 470553;
srom_1(65656) <= 299540;
srom_1(65657) <= 166460;
srom_1(65658) <= 71936;
srom_1(65659) <= 16411;
srom_1(65660) <= 147;
srom_1(65661) <= 23219;
srom_1(65662) <= 85519;
srom_1(65663) <= 186755;
srom_1(65664) <= 326453;
srom_1(65665) <= 503957;
srom_1(65666) <= 718434;
srom_1(65667) <= 968880;
srom_1(65668) <= 1254119;
srom_1(65669) <= 1572815;
srom_1(65670) <= 1923472;
srom_1(65671) <= 2304446;
srom_1(65672) <= 2713951;
srom_1(65673) <= 3150066;
srom_1(65674) <= 3610747;
srom_1(65675) <= 4093832;
srom_1(65676) <= 4597058;
srom_1(65677) <= 5118063;
srom_1(65678) <= 5654405;
srom_1(65679) <= 6203568;
srom_1(65680) <= 6762978;
srom_1(65681) <= 7330011;
srom_1(65682) <= 7902009;
srom_1(65683) <= 8476288;
srom_1(65684) <= 9050155;
srom_1(65685) <= 9620921;
srom_1(65686) <= 10185908;
srom_1(65687) <= 10742467;
srom_1(65688) <= 11287987;
srom_1(65689) <= 11819912;
srom_1(65690) <= 12335745;
srom_1(65691) <= 12833070;
srom_1(65692) <= 13309553;
srom_1(65693) <= 13762959;
srom_1(65694) <= 14191164;
srom_1(65695) <= 14592158;
srom_1(65696) <= 14964062;
srom_1(65697) <= 15305131;
srom_1(65698) <= 15613767;
srom_1(65699) <= 15888521;
srom_1(65700) <= 16128105;
srom_1(65701) <= 16331396;
srom_1(65702) <= 16497441;
srom_1(65703) <= 16625460;
srom_1(65704) <= 16714855;
srom_1(65705) <= 16765204;
srom_1(65706) <= 16776273;
srom_1(65707) <= 16748009;
srom_1(65708) <= 16680545;
srom_1(65709) <= 16574197;
srom_1(65710) <= 16429464;
srom_1(65711) <= 16247025;
srom_1(65712) <= 16027735;
srom_1(65713) <= 15772623;
srom_1(65714) <= 15482884;
srom_1(65715) <= 15159878;
srom_1(65716) <= 14805119;
srom_1(65717) <= 14420271;
srom_1(65718) <= 14007138;
srom_1(65719) <= 13567658;
srom_1(65720) <= 13103892;
srom_1(65721) <= 12618014;
srom_1(65722) <= 12112303;
srom_1(65723) <= 11589130;
srom_1(65724) <= 11050949;
srom_1(65725) <= 10500283;
srom_1(65726) <= 9939715;
srom_1(65727) <= 9371873;
srom_1(65728) <= 8799421;
srom_1(65729) <= 8225041;
srom_1(65730) <= 7651429;
srom_1(65731) <= 7081274;
srom_1(65732) <= 6517249;
srom_1(65733) <= 5962000;
srom_1(65734) <= 5418130;
srom_1(65735) <= 4888190;
srom_1(65736) <= 4374664;
srom_1(65737) <= 3879961;
srom_1(65738) <= 3406400;
srom_1(65739) <= 2956203;
srom_1(65740) <= 2531480;
srom_1(65741) <= 2134223;
srom_1(65742) <= 1766296;
srom_1(65743) <= 1429422;
srom_1(65744) <= 1125183;
srom_1(65745) <= 855004;
srom_1(65746) <= 620153;
srom_1(65747) <= 421730;
srom_1(65748) <= 260668;
srom_1(65749) <= 137720;
srom_1(65750) <= 53463;
srom_1(65751) <= 8292;
srom_1(65752) <= 2420;
srom_1(65753) <= 35873;
srom_1(65754) <= 108496;
srom_1(65755) <= 219946;
srom_1(65756) <= 369702;
srom_1(65757) <= 557062;
srom_1(65758) <= 781146;
srom_1(65759) <= 1040905;
srom_1(65760) <= 1335119;
srom_1(65761) <= 1662409;
srom_1(65762) <= 2021241;
srom_1(65763) <= 2409932;
srom_1(65764) <= 2826659;
srom_1(65765) <= 3269467;
srom_1(65766) <= 3736282;
srom_1(65767) <= 4224912;
srom_1(65768) <= 4733067;
srom_1(65769) <= 5258365;
srom_1(65770) <= 5798341;
srom_1(65771) <= 6350464;
srom_1(65772) <= 6912144;
srom_1(65773) <= 7480748;
srom_1(65774) <= 8053610;
srom_1(65775) <= 8628042;
srom_1(65776) <= 9201352;
srom_1(65777) <= 9770850;
srom_1(65778) <= 10333866;
srom_1(65779) <= 10887761;
srom_1(65780) <= 11429936;
srom_1(65781) <= 11957849;
srom_1(65782) <= 12469025;
srom_1(65783) <= 12961066;
srom_1(65784) <= 13431665;
srom_1(65785) <= 13878616;
srom_1(65786) <= 14299823;
srom_1(65787) <= 14693309;
srom_1(65788) <= 15057231;
srom_1(65789) <= 15389881;
srom_1(65790) <= 15689700;
srom_1(65791) <= 15955281;
srom_1(65792) <= 16185380;
srom_1(65793) <= 16378917;
srom_1(65794) <= 16534985;
srom_1(65795) <= 16652851;
srom_1(65796) <= 16731964;
srom_1(65797) <= 16771951;
srom_1(65798) <= 16772627;
srom_1(65799) <= 16733987;
srom_1(65800) <= 16656212;
srom_1(65801) <= 16539668;
srom_1(65802) <= 16384901;
srom_1(65803) <= 16192636;
srom_1(65804) <= 15963775;
srom_1(65805) <= 15699392;
srom_1(65806) <= 15400727;
srom_1(65807) <= 15069179;
srom_1(65808) <= 14706303;
srom_1(65809) <= 14313802;
srom_1(65810) <= 13893515;
srom_1(65811) <= 13447414;
srom_1(65812) <= 12977590;
srom_1(65813) <= 12486247;
srom_1(65814) <= 11975689;
srom_1(65815) <= 11448310;
srom_1(65816) <= 10906583;
srom_1(65817) <= 10353048;
srom_1(65818) <= 9790301;
srom_1(65819) <= 9220981;
srom_1(65820) <= 8647758;
srom_1(65821) <= 8073320;
srom_1(65822) <= 7500360;
srom_1(65823) <= 6931565;
srom_1(65824) <= 6369603;
srom_1(65825) <= 5817109;
srom_1(65826) <= 5276674;
srom_1(65827) <= 4750831;
srom_1(65828) <= 4242047;
srom_1(65829) <= 3752708;
srom_1(65830) <= 3285108;
srom_1(65831) <= 2841440;
srom_1(65832) <= 2423785;
srom_1(65833) <= 2034101;
srom_1(65834) <= 1674215;
srom_1(65835) <= 1345815;
srom_1(65836) <= 1050442;
srom_1(65837) <= 789479;
srom_1(65838) <= 564152;
srom_1(65839) <= 375516;
srom_1(65840) <= 224456;
srom_1(65841) <= 111681;
srom_1(65842) <= 37719;
srom_1(65843) <= 2917;
srom_1(65844) <= 7439;
srom_1(65845) <= 51262;
srom_1(65846) <= 134183;
srom_1(65847) <= 255811;
srom_1(65848) <= 415577;
srom_1(65849) <= 612731;
srom_1(65850) <= 846349;
srom_1(65851) <= 1115335;
srom_1(65852) <= 1418428;
srom_1(65853) <= 1754206;
srom_1(65854) <= 2121096;
srom_1(65855) <= 2517376;
srom_1(65856) <= 2941188;
srom_1(65857) <= 3390545;
srom_1(65858) <= 3863339;
srom_1(65859) <= 4357355;
srom_1(65860) <= 4870274;
srom_1(65861) <= 5399691;
srom_1(65862) <= 5943125;
srom_1(65863) <= 6498027;
srom_1(65864) <= 7061794;
srom_1(65865) <= 7631783;
srom_1(65866) <= 8205321;
srom_1(65867) <= 8779718;
srom_1(65868) <= 9352282;
srom_1(65869) <= 9920326;
srom_1(65870) <= 10481188;
srom_1(65871) <= 11032236;
srom_1(65872) <= 11570888;
srom_1(65873) <= 12094617;
srom_1(65874) <= 12600968;
srom_1(65875) <= 13087565;
srom_1(65876) <= 13552127;
srom_1(65877) <= 13992476;
srom_1(65878) <= 14406546;
srom_1(65879) <= 14792396;
srom_1(65880) <= 15148216;
srom_1(65881) <= 15472338;
srom_1(65882) <= 15763243;
srom_1(65883) <= 16019564;
srom_1(65884) <= 16240102;
srom_1(65885) <= 16423822;
srom_1(65886) <= 16569861;
srom_1(65887) <= 16677536;
srom_1(65888) <= 16746341;
srom_1(65889) <= 16775954;
srom_1(65890) <= 16766236;
srom_1(65891) <= 16717232;
srom_1(65892) <= 16629173;
srom_1(65893) <= 16502470;
srom_1(65894) <= 16337719;
srom_1(65895) <= 16135692;
srom_1(65896) <= 15897336;
srom_1(65897) <= 15623769;
srom_1(65898) <= 15316273;
srom_1(65899) <= 14976292;
srom_1(65900) <= 14605419;
srom_1(65901) <= 14205393;
srom_1(65902) <= 13778090;
srom_1(65903) <= 13325513;
srom_1(65904) <= 12849786;
srom_1(65905) <= 12353139;
srom_1(65906) <= 11837901;
srom_1(65907) <= 11306488;
srom_1(65908) <= 10761392;
srom_1(65909) <= 10205170;
srom_1(65910) <= 9640429;
srom_1(65911) <= 9069817;
srom_1(65912) <= 8496011;
srom_1(65913) <= 7921702;
srom_1(65914) <= 7349582;
srom_1(65915) <= 6782334;
srom_1(65916) <= 6222619;
srom_1(65917) <= 5673060;
srom_1(65918) <= 5136236;
srom_1(65919) <= 4614663;
srom_1(65920) <= 4110788;
srom_1(65921) <= 3626973;
srom_1(65922) <= 3165487;
srom_1(65923) <= 2728493;
srom_1(65924) <= 2318042;
srom_1(65925) <= 1936058;
srom_1(65926) <= 1584332;
srom_1(65927) <= 1264514;
srom_1(65928) <= 978103;
srom_1(65929) <= 726442;
srom_1(65930) <= 510712;
srom_1(65931) <= 331924;
srom_1(65932) <= 190917;
srom_1(65933) <= 88352;
srom_1(65934) <= 24709;
srom_1(65935) <= 287;
srom_1(65936) <= 15201;
srom_1(65937) <= 69381;
srom_1(65938) <= 162573;
srom_1(65939) <= 294339;
srom_1(65940) <= 464062;
srom_1(65941) <= 670946;
srom_1(65942) <= 914021;
srom_1(65943) <= 1192146;
srom_1(65944) <= 1504019;
srom_1(65945) <= 1848175;
srom_1(65946) <= 2223002;
srom_1(65947) <= 2626741;
srom_1(65948) <= 3057500;
srom_1(65949) <= 3513258;
srom_1(65950) <= 3991879;
srom_1(65951) <= 4491117;
srom_1(65952) <= 5008632;
srom_1(65953) <= 5541997;
srom_1(65954) <= 6088710;
srom_1(65955) <= 6646208;
srom_1(65956) <= 7211878;
srom_1(65957) <= 7783065;
srom_1(65958) <= 8357092;
srom_1(65959) <= 8931266;
srom_1(65960) <= 9502896;
srom_1(65961) <= 10069301;
srom_1(65962) <= 10627824;
srom_1(65963) <= 11175847;
srom_1(65964) <= 11710799;
srom_1(65965) <= 12230173;
srom_1(65966) <= 12731532;
srom_1(65967) <= 13212526;
srom_1(65968) <= 13670898;
srom_1(65969) <= 14104500;
srom_1(65970) <= 14511299;
srom_1(65971) <= 14889386;
srom_1(65972) <= 15236988;
srom_1(65973) <= 15552477;
srom_1(65974) <= 15834371;
srom_1(65975) <= 16081349;
srom_1(65976) <= 16292254;
srom_1(65977) <= 16466096;
srom_1(65978) <= 16602060;
srom_1(65979) <= 16699507;
srom_1(65980) <= 16757983;
srom_1(65981) <= 16777211;
srom_1(65982) <= 16757102;
srom_1(65983) <= 16697751;
srom_1(65984) <= 16599435;
srom_1(65985) <= 16462616;
srom_1(65986) <= 16287935;
srom_1(65987) <= 16076211;
srom_1(65988) <= 15828437;
srom_1(65989) <= 15545776;
srom_1(65990) <= 15229552;
srom_1(65991) <= 14881249;
srom_1(65992) <= 14502499;
srom_1(65993) <= 14095079;
srom_1(65994) <= 13660900;
srom_1(65995) <= 13201997;
srom_1(65996) <= 12720522;
srom_1(65997) <= 12218734;
srom_1(65998) <= 11698984;
srom_1(65999) <= 11163711;
srom_1(66000) <= 10615425;
srom_1(66001) <= 10056697;
srom_1(66002) <= 9490146;
srom_1(66003) <= 8918430;
srom_1(66004) <= 8344229;
srom_1(66005) <= 7770236;
srom_1(66006) <= 7199143;
srom_1(66007) <= 6633628;
srom_1(66008) <= 6076343;
srom_1(66009) <= 5529900;
srom_1(66010) <= 4996863;
srom_1(66011) <= 4479731;
srom_1(66012) <= 3980929;
srom_1(66013) <= 3502797;
srom_1(66014) <= 3047575;
srom_1(66015) <= 2617400;
srom_1(66016) <= 2214287;
srom_1(66017) <= 1840128;
srom_1(66018) <= 1496677;
srom_1(66019) <= 1185545;
srom_1(66020) <= 908191;
srom_1(66021) <= 665914;
srom_1(66022) <= 459852;
srom_1(66023) <= 290971;
srom_1(66024) <= 160062;
srom_1(66025) <= 67740;
srom_1(66026) <= 14437;
srom_1(66027) <= 403;
srom_1(66028) <= 25705;
srom_1(66029) <= 90223;
srom_1(66030) <= 193655;
srom_1(66031) <= 335516;
srom_1(66032) <= 515141;
srom_1(66033) <= 731687;
srom_1(66034) <= 984140;
srom_1(66035) <= 1271314;
srom_1(66036) <= 1591863;
srom_1(66037) <= 1944285;
srom_1(66038) <= 2326927;
srom_1(66039) <= 2737993;
srom_1(66040) <= 3175558;
srom_1(66041) <= 3637568;
srom_1(66042) <= 4121858;
srom_1(66043) <= 4626155;
srom_1(66044) <= 5148097;
srom_1(66045) <= 5685234;
srom_1(66046) <= 6235048;
srom_1(66047) <= 6794961;
srom_1(66048) <= 7362347;
srom_1(66049) <= 7934545;
srom_1(66050) <= 8508873;
srom_1(66051) <= 9082637;
srom_1(66052) <= 9653146;
srom_1(66053) <= 10217725;
srom_1(66054) <= 10773727;
srom_1(66055) <= 11318545;
srom_1(66056) <= 11849623;
srom_1(66057) <= 12364471;
srom_1(66058) <= 12860674;
srom_1(66059) <= 13335907;
srom_1(66060) <= 13787940;
srom_1(66061) <= 14214654;
srom_1(66062) <= 14614047;
srom_1(66063) <= 14984248;
srom_1(66064) <= 15323519;
srom_1(66065) <= 15630269;
srom_1(66066) <= 15903062;
srom_1(66067) <= 16140616;
srom_1(66068) <= 16341818;
srom_1(66069) <= 16505726;
srom_1(66070) <= 16631569;
srom_1(66071) <= 16718758;
srom_1(66072) <= 16766884;
srom_1(66073) <= 16775721;
srom_1(66074) <= 16745229;
srom_1(66075) <= 16675549;
srom_1(66076) <= 16567009;
srom_1(66077) <= 16420118;
srom_1(66078) <= 16235564;
srom_1(66079) <= 16014213;
srom_1(66080) <= 15757104;
srom_1(66081) <= 15465440;
srom_1(66082) <= 15140591;
srom_1(66083) <= 14784080;
srom_1(66084) <= 14397578;
srom_1(66085) <= 13982897;
srom_1(66086) <= 13541984;
srom_1(66087) <= 13076904;
srom_1(66088) <= 12589839;
srom_1(66089) <= 12083074;
srom_1(66090) <= 11558983;
srom_1(66091) <= 11020026;
srom_1(66092) <= 10468729;
srom_1(66093) <= 9907678;
srom_1(66094) <= 9339503;
srom_1(66095) <= 8766869;
srom_1(66096) <= 8192461;
srom_1(66097) <= 7618973;
srom_1(66098) <= 7049094;
srom_1(66099) <= 6485497;
srom_1(66100) <= 5930824;
srom_1(66101) <= 5387676;
srom_1(66102) <= 4858601;
srom_1(66103) <= 4346079;
srom_1(66104) <= 3852514;
srom_1(66105) <= 3380220;
srom_1(66106) <= 2931412;
srom_1(66107) <= 2508195;
srom_1(66108) <= 2112554;
srom_1(66109) <= 1746342;
srom_1(66110) <= 1411279;
srom_1(66111) <= 1108935;
srom_1(66112) <= 840727;
srom_1(66113) <= 607914;
srom_1(66114) <= 411588;
srom_1(66115) <= 252668;
srom_1(66116) <= 131901;
srom_1(66117) <= 49852;
srom_1(66118) <= 6907;
srom_1(66119) <= 3266;
srom_1(66120) <= 38947;
srom_1(66121) <= 113782;
srom_1(66122) <= 227421;
srom_1(66123) <= 379331;
srom_1(66124) <= 568798;
srom_1(66125) <= 794936;
srom_1(66126) <= 1056683;
srom_1(66127) <= 1352811;
srom_1(66128) <= 1681933;
srom_1(66129) <= 2042505;
srom_1(66130) <= 2432836;
srom_1(66131) <= 2851096;
srom_1(66132) <= 3295322;
srom_1(66133) <= 3763433;
srom_1(66134) <= 4253233;
srom_1(66135) <= 4762426;
srom_1(66136) <= 5288622;
srom_1(66137) <= 5829356;
srom_1(66138) <= 6382091;
srom_1(66139) <= 6944235;
srom_1(66140) <= 7513152;
srom_1(66141) <= 8086174;
srom_1(66142) <= 8660615;
srom_1(66143) <= 9233780;
srom_1(66144) <= 9802982;
srom_1(66145) <= 10365551;
srom_1(66146) <= 10918850;
srom_1(66147) <= 11460283;
srom_1(66148) <= 11987313;
srom_1(66149) <= 12497466;
srom_1(66150) <= 12988352;
srom_1(66151) <= 13457669;
srom_1(66152) <= 13903214;
srom_1(66153) <= 14322900;
srom_1(66154) <= 14714758;
srom_1(66155) <= 15076950;
srom_1(66156) <= 15407778;
srom_1(66157) <= 15705691;
srom_1(66158) <= 15969292;
srom_1(66159) <= 16197344;
srom_1(66160) <= 16388779;
srom_1(66161) <= 16542698;
srom_1(66162) <= 16658379;
srom_1(66163) <= 16735281;
srom_1(66164) <= 16773042;
srom_1(66165) <= 16771486;
srom_1(66166) <= 16730620;
srom_1(66167) <= 16650635;
srom_1(66168) <= 16531906;
srom_1(66169) <= 16374991;
srom_1(66170) <= 16180625;
srom_1(66171) <= 15949719;
srom_1(66172) <= 15683357;
srom_1(66173) <= 15382787;
srom_1(66174) <= 15049420;
srom_1(66175) <= 14684817;
srom_1(66176) <= 14290689;
srom_1(66177) <= 13868884;
srom_1(66178) <= 13421381;
srom_1(66179) <= 12950276;
srom_1(66180) <= 12457781;
srom_1(66181) <= 11946204;
srom_1(66182) <= 11417944;
srom_1(66183) <= 10875479;
srom_1(66184) <= 10321352;
srom_1(66185) <= 9758161;
srom_1(66186) <= 9188548;
srom_1(66187) <= 8615184;
srom_1(66188) <= 8040758;
srom_1(66189) <= 7467962;
srom_1(66190) <= 6899484;
srom_1(66191) <= 6337989;
srom_1(66192) <= 5786110;
srom_1(66193) <= 5246435;
srom_1(66194) <= 4721494;
srom_1(66195) <= 4213750;
srom_1(66196) <= 3725584;
srom_1(66197) <= 3259283;
srom_1(66198) <= 2817036;
srom_1(66199) <= 2400916;
srom_1(66200) <= 2012875;
srom_1(66201) <= 1654731;
srom_1(66202) <= 1328165;
srom_1(66203) <= 1034707;
srom_1(66204) <= 775735;
srom_1(66205) <= 552462;
srom_1(66206) <= 365935;
srom_1(66207) <= 217030;
srom_1(66208) <= 106443;
srom_1(66209) <= 34695;
srom_1(66210) <= 2121;
srom_1(66211) <= 8874;
srom_1(66212) <= 54922;
srom_1(66213) <= 140051;
srom_1(66214) <= 263859;
srom_1(66215) <= 425767;
srom_1(66216) <= 625016;
srom_1(66217) <= 860670;
srom_1(66218) <= 1131626;
srom_1(66219) <= 1436612;
srom_1(66220) <= 1774199;
srom_1(66221) <= 2142803;
srom_1(66222) <= 2540695;
srom_1(66223) <= 2966011;
srom_1(66224) <= 3416754;
srom_1(66225) <= 3890813;
srom_1(66226) <= 4385963;
srom_1(66227) <= 4899883;
srom_1(66228) <= 5430163;
srom_1(66229) <= 5974316;
srom_1(66230) <= 6529790;
srom_1(66231) <= 7093981;
srom_1(66232) <= 7664243;
srom_1(66233) <= 8237902;
srom_1(66234) <= 8812268;
srom_1(66235) <= 9384646;
srom_1(66236) <= 9952354;
srom_1(66237) <= 10512729;
srom_1(66238) <= 11063144;
srom_1(66239) <= 11601016;
srom_1(66240) <= 12123825;
srom_1(66241) <= 12629117;
srom_1(66242) <= 13114525;
srom_1(66243) <= 13577771;
srom_1(66244) <= 14016683;
srom_1(66245) <= 14429203;
srom_1(66246) <= 14813397;
srom_1(66247) <= 15167463;
srom_1(66248) <= 15489740;
srom_1(66249) <= 15778718;
srom_1(66250) <= 16033041;
srom_1(66251) <= 16251516;
srom_1(66252) <= 16433120;
srom_1(66253) <= 16577000;
srom_1(66254) <= 16682482;
srom_1(66255) <= 16749071;
srom_1(66256) <= 16776456;
srom_1(66257) <= 16764506;
srom_1(66258) <= 16713279;
srom_1(66259) <= 16623015;
srom_1(66260) <= 16494137;
srom_1(66261) <= 16327249;
srom_1(66262) <= 16123134;
srom_1(66263) <= 15882750;
srom_1(66264) <= 15607223;
srom_1(66265) <= 15297845;
srom_1(66266) <= 14956067;
srom_1(66267) <= 14583493;
srom_1(66268) <= 14181868;
srom_1(66269) <= 13753077;
srom_1(66270) <= 13299130;
srom_1(66271) <= 12822155;
srom_1(66272) <= 12324391;
srom_1(66273) <= 11808170;
srom_1(66274) <= 11275914;
srom_1(66275) <= 10730118;
srom_1(66276) <= 10173342;
srom_1(66277) <= 9608196;
srom_1(66278) <= 9037332;
srom_1(66279) <= 8463425;
srom_1(66280) <= 7889168;
srom_1(66281) <= 7317253;
srom_1(66282) <= 6750361;
srom_1(66283) <= 6191152;
srom_1(66284) <= 5642248;
srom_1(66285) <= 5106222;
srom_1(66286) <= 4585588;
srom_1(66287) <= 4082788;
srom_1(66288) <= 3600180;
srom_1(66289) <= 3140026;
srom_1(66290) <= 2704484;
srom_1(66291) <= 2295598;
srom_1(66292) <= 1915283;
srom_1(66293) <= 1565324;
srom_1(66294) <= 1247362;
srom_1(66295) <= 962888;
srom_1(66296) <= 713235;
srom_1(66297) <= 499575;
srom_1(66298) <= 322909;
srom_1(66299) <= 184066;
srom_1(66300) <= 83697;
srom_1(66301) <= 22272;
srom_1(66302) <= 81;
srom_1(66303) <= 17225;
srom_1(66304) <= 73626;
srom_1(66305) <= 169019;
srom_1(66306) <= 302957;
srom_1(66307) <= 474810;
srom_1(66308) <= 683775;
srom_1(66309) <= 928869;
srom_1(66310) <= 1208945;
srom_1(66311) <= 1522689;
srom_1(66312) <= 1868630;
srom_1(66313) <= 2245145;
srom_1(66314) <= 2650469;
srom_1(66315) <= 3082701;
srom_1(66316) <= 3539814;
srom_1(66317) <= 4019665;
srom_1(66318) <= 4520003;
srom_1(66319) <= 5038483;
srom_1(66320) <= 5572672;
srom_1(66321) <= 6120066;
srom_1(66322) <= 6678099;
srom_1(66323) <= 7244152;
srom_1(66324) <= 7815572;
srom_1(66325) <= 8389679;
srom_1(66326) <= 8963782;
srom_1(66327) <= 9535187;
srom_1(66328) <= 10101215;
srom_1(66329) <= 10659212;
srom_1(66330) <= 11206562;
srom_1(66331) <= 11740697;
srom_1(66332) <= 12259114;
srom_1(66333) <= 12759380;
srom_1(66334) <= 13239150;
srom_1(66335) <= 13696174;
srom_1(66336) <= 14128309;
srom_1(66337) <= 14533529;
srom_1(66338) <= 14909933;
srom_1(66339) <= 15255756;
srom_1(66340) <= 15569377;
srom_1(66341) <= 15849325;
srom_1(66342) <= 16094287;
srom_1(66343) <= 16303114;
srom_1(66344) <= 16474828;
srom_1(66345) <= 16608622;
srom_1(66346) <= 16703870;
srom_1(66347) <= 16760125;
srom_1(66348) <= 16777123;
srom_1(66349) <= 16754784;
srom_1(66350) <= 16693213;
srom_1(66351) <= 16592700;
srom_1(66352) <= 16453714;
srom_1(66353) <= 16276908;
srom_1(66354) <= 16063112;
srom_1(66355) <= 15813327;
srom_1(66356) <= 15528725;
srom_1(66357) <= 15210640;
srom_1(66358) <= 14860565;
srom_1(66359) <= 14480140;
srom_1(66360) <= 14071150;
srom_1(66361) <= 13635513;
srom_1(66362) <= 13175271;
srom_1(66363) <= 12692583;
srom_1(66364) <= 12189712;
srom_1(66365) <= 11669016;
srom_1(66366) <= 11132938;
srom_1(66367) <= 10583990;
srom_1(66368) <= 10024747;
srom_1(66369) <= 9457832;
srom_1(66370) <= 8885903;
srom_1(66371) <= 8311642;
srom_1(66372) <= 7737742;
srom_1(66373) <= 7166894;
srom_1(66374) <= 6601775;
srom_1(66375) <= 6045035;
srom_1(66376) <= 5499285;
srom_1(66377) <= 4967084;
srom_1(66378) <= 4450927;
srom_1(66379) <= 3953236;
srom_1(66380) <= 3476344;
srom_1(66381) <= 3022487;
srom_1(66382) <= 2593793;
srom_1(66383) <= 2192274;
srom_1(66384) <= 1819811;
srom_1(66385) <= 1478151;
srom_1(66386) <= 1168897;
srom_1(66387) <= 893499;
srom_1(66388) <= 653248;
srom_1(66389) <= 449271;
srom_1(66390) <= 282524;
srom_1(66391) <= 153789;
srom_1(66392) <= 63670;
srom_1(66393) <= 12589;
srom_1(66394) <= 787;
srom_1(66395) <= 28317;
srom_1(66396) <= 95053;
srom_1(66397) <= 200679;
srom_1(66398) <= 344701;
srom_1(66399) <= 526445;
srom_1(66400) <= 745056;
srom_1(66401) <= 999511;
srom_1(66402) <= 1288615;
srom_1(66403) <= 1611014;
srom_1(66404) <= 1965196;
srom_1(66405) <= 2349499;
srom_1(66406) <= 2762121;
srom_1(66407) <= 3201128;
srom_1(66408) <= 3664461;
srom_1(66409) <= 4149947;
srom_1(66410) <= 4655310;
srom_1(66411) <= 5178179;
srom_1(66412) <= 5716103;
srom_1(66413) <= 6266560;
srom_1(66414) <= 6826967;
srom_1(66415) <= 7394697;
srom_1(66416) <= 7967089;
srom_1(66417) <= 8541456;
srom_1(66418) <= 9115107;
srom_1(66419) <= 9685352;
srom_1(66420) <= 10249515;
srom_1(66421) <= 10804952;
srom_1(66422) <= 11349058;
srom_1(66423) <= 11879281;
srom_1(66424) <= 12393136;
srom_1(66425) <= 12888211;
srom_1(66426) <= 13362187;
srom_1(66427) <= 13812839;
srom_1(66428) <= 14238056;
srom_1(66429) <= 14635843;
srom_1(66430) <= 15004334;
srom_1(66431) <= 15341801;
srom_1(66432) <= 15646663;
srom_1(66433) <= 15917489;
srom_1(66434) <= 16153010;
srom_1(66435) <= 16352121;
srom_1(66436) <= 16513888;
srom_1(66437) <= 16637553;
srom_1(66438) <= 16722535;
srom_1(66439) <= 16768437;
srom_1(66440) <= 16775044;
srom_1(66441) <= 16742323;
srom_1(66442) <= 16670429;
srom_1(66443) <= 16559698;
srom_1(66444) <= 16410651;
srom_1(66445) <= 16223985;
srom_1(66446) <= 16000577;
srom_1(66447) <= 15741473;
srom_1(66448) <= 15447889;
srom_1(66449) <= 15121202;
srom_1(66450) <= 14762944;
srom_1(66451) <= 14374794;
srom_1(66452) <= 13958572;
srom_1(66453) <= 13516231;
srom_1(66454) <= 13049846;
srom_1(66455) <= 12561601;
srom_1(66456) <= 12053789;
srom_1(66457) <= 11528789;
srom_1(66458) <= 10989063;
srom_1(66459) <= 10437143;
srom_1(66460) <= 9875617;
srom_1(66461) <= 9307118;
srom_1(66462) <= 8734311;
srom_1(66463) <= 8159884;
srom_1(66464) <= 7586529;
srom_1(66465) <= 7016935;
srom_1(66466) <= 6453773;
srom_1(66467) <= 5899685;
srom_1(66468) <= 5357268;
srom_1(66469) <= 4829066;
srom_1(66470) <= 4317555;
srom_1(66471) <= 3825136;
srom_1(66472) <= 3354116;
srom_1(66473) <= 2906704;
srom_1(66474) <= 2484999;
srom_1(66475) <= 2090978;
srom_1(66476) <= 1726489;
srom_1(66477) <= 1393241;
srom_1(66478) <= 1092797;
srom_1(66479) <= 826565;
srom_1(66480) <= 595794;
srom_1(66481) <= 401566;
srom_1(66482) <= 244792;
srom_1(66483) <= 126207;
srom_1(66484) <= 46368;
srom_1(66485) <= 5648;
srom_1(66486) <= 4239;
srom_1(66487) <= 42147;
srom_1(66488) <= 119194;
srom_1(66489) <= 235019;
srom_1(66490) <= 389080;
srom_1(66491) <= 580653;
srom_1(66492) <= 808840;
srom_1(66493) <= 1072571;
srom_1(66494) <= 1370610;
srom_1(66495) <= 1701558;
srom_1(66496) <= 2063865;
srom_1(66497) <= 2455830;
srom_1(66498) <= 2875616;
srom_1(66499) <= 3321254;
srom_1(66500) <= 3790655;
srom_1(66501) <= 4281617;
srom_1(66502) <= 4791839;
srom_1(66503) <= 5318927;
srom_1(66504) <= 5860409;
srom_1(66505) <= 6413748;
srom_1(66506) <= 6976347;
srom_1(66507) <= 7545568;
srom_1(66508) <= 8118743;
srom_1(66509) <= 8693183;
srom_1(66510) <= 9266195;
srom_1(66511) <= 9835092;
srom_1(66512) <= 10397206;
srom_1(66513) <= 10949901;
srom_1(66514) <= 11490584;
srom_1(66515) <= 12016722;
srom_1(66516) <= 12525846;
srom_1(66517) <= 13015570;
srom_1(66518) <= 13483595;
srom_1(66519) <= 13927729;
srom_1(66520) <= 14345888;
srom_1(66521) <= 14736111;
srom_1(66522) <= 15096568;
srom_1(66523) <= 15425570;
srom_1(66524) <= 15721573;
srom_1(66525) <= 15983189;
srom_1(66526) <= 16209191;
srom_1(66527) <= 16398520;
srom_1(66528) <= 16550288;
srom_1(66529) <= 16663783;
srom_1(66530) <= 16738472;
srom_1(66531) <= 16774007;
srom_1(66532) <= 16770219;
srom_1(66533) <= 16727127;
srom_1(66534) <= 16644933;
srom_1(66535) <= 16524022;
srom_1(66536) <= 16364961;
srom_1(66537) <= 16168496;
srom_1(66538) <= 15935549;
srom_1(66539) <= 15667212;
srom_1(66540) <= 15364743;
srom_1(66541) <= 15029560;
srom_1(66542) <= 14663235;
srom_1(66543) <= 14267487;
srom_1(66544) <= 13844171;
srom_1(66545) <= 13395271;
srom_1(66546) <= 12922894;
srom_1(66547) <= 12429254;
srom_1(66548) <= 11916665;
srom_1(66549) <= 11387533;
srom_1(66550) <= 10844337;
srom_1(66551) <= 10289626;
srom_1(66552) <= 9726000;
srom_1(66553) <= 9156103;
srom_1(66554) <= 8582607;
srom_1(66555) <= 8008201;
srom_1(66556) <= 7435578;
srom_1(66557) <= 6867425;
srom_1(66558) <= 6306405;
srom_1(66559) <= 5755150;
srom_1(66560) <= 5216243;
srom_1(66561) <= 4692213;
srom_1(66562) <= 4185516;
srom_1(66563) <= 3698530;
srom_1(66564) <= 3233536;
srom_1(66565) <= 2792717;
srom_1(66566) <= 2378138;
srom_1(66567) <= 1991745;
srom_1(66568) <= 1635349;
srom_1(66569) <= 1310621;
srom_1(66570) <= 1019084;
srom_1(66571) <= 762106;
srom_1(66572) <= 540890;
srom_1(66573) <= 356476;
srom_1(66574) <= 209726;
srom_1(66575) <= 101331;
srom_1(66576) <= 31797;
srom_1(66577) <= 1451;
srom_1(66578) <= 10436;
srom_1(66579) <= 58708;
srom_1(66580) <= 146043;
srom_1(66581) <= 272029;
srom_1(66582) <= 436077;
srom_1(66583) <= 637417;
srom_1(66584) <= 875105;
srom_1(66585) <= 1148027;
srom_1(66586) <= 1454902;
srom_1(66587) <= 1794291;
srom_1(66588) <= 2164604;
srom_1(66589) <= 2564103;
srom_1(66590) <= 2990915;
srom_1(66591) <= 3443039;
srom_1(66592) <= 3918354;
srom_1(66593) <= 4414632;
srom_1(66594) <= 4929545;
srom_1(66595) <= 5460679;
srom_1(66596) <= 6005543;
srom_1(66597) <= 6561582;
srom_1(66598) <= 7126188;
srom_1(66599) <= 7696715;
srom_1(66600) <= 8270486;
srom_1(66601) <= 8844811;
srom_1(66602) <= 9416996;
srom_1(66603) <= 9984359;
srom_1(66604) <= 10544239;
srom_1(66605) <= 11094011;
srom_1(66606) <= 11631096;
srom_1(66607) <= 12152975;
srom_1(66608) <= 12657203;
srom_1(66609) <= 13141413;
srom_1(66610) <= 13603336;
srom_1(66611) <= 14040805;
srom_1(66612) <= 14451769;
srom_1(66613) <= 14834301;
srom_1(66614) <= 15186607;
srom_1(66615) <= 15507035;
srom_1(66616) <= 15794082;
srom_1(66617) <= 16046402;
srom_1(66618) <= 16262812;
srom_1(66619) <= 16442297;
srom_1(66620) <= 16584016;
srom_1(66621) <= 16687303;
srom_1(66622) <= 16751675;
srom_1(66623) <= 16776830;
srom_1(66624) <= 16762650;
srom_1(66625) <= 16709201;
srom_1(66626) <= 16616733;
srom_1(66627) <= 16485682;
srom_1(66628) <= 16316660;
srom_1(66629) <= 16110461;
srom_1(66630) <= 15868051;
srom_1(66631) <= 15590568;
srom_1(66632) <= 15279312;
srom_1(66633) <= 14935743;
srom_1(66634) <= 14561473;
srom_1(66635) <= 14158256;
srom_1(66636) <= 13727983;
srom_1(66637) <= 13272672;
srom_1(66638) <= 12794458;
srom_1(66639) <= 12295583;
srom_1(66640) <= 11778387;
srom_1(66641) <= 11245295;
srom_1(66642) <= 10698808;
srom_1(66643) <= 10141486;
srom_1(66644) <= 9575946;
srom_1(66645) <= 9004837;
srom_1(66646) <= 8430838;
srom_1(66647) <= 7856642;
srom_1(66648) <= 7284940;
srom_1(66649) <= 6718413;
srom_1(66650) <= 6159719;
srom_1(66651) <= 5611477;
srom_1(66652) <= 5076257;
srom_1(66653) <= 4556571;
srom_1(66654) <= 4054854;
srom_1(66655) <= 3573459;
srom_1(66656) <= 3114644;
srom_1(66657) <= 2680561;
srom_1(66658) <= 2273245;
srom_1(66659) <= 1894606;
srom_1(66660) <= 1546419;
srom_1(66661) <= 1230318;
srom_1(66662) <= 947785;
srom_1(66663) <= 700144;
srom_1(66664) <= 488556;
srom_1(66665) <= 314015;
srom_1(66666) <= 177339;
srom_1(66667) <= 79168;
srom_1(66668) <= 19962;
srom_1(66669) <= 1;
srom_1(66670) <= 19376;
srom_1(66671) <= 77997;
srom_1(66672) <= 175590;
srom_1(66673) <= 311696;
srom_1(66674) <= 485678;
srom_1(66675) <= 696719;
srom_1(66676) <= 943831;
srom_1(66677) <= 1225853;
srom_1(66678) <= 1541464;
srom_1(66679) <= 1889184;
srom_1(66680) <= 2267381;
srom_1(66681) <= 2674283;
srom_1(66682) <= 3107982;
srom_1(66683) <= 3566443;
srom_1(66684) <= 4047517;
srom_1(66685) <= 4548948;
srom_1(66686) <= 5068384;
srom_1(66687) <= 5603390;
srom_1(66688) <= 6151457;
srom_1(66689) <= 6710015;
srom_1(66690) <= 7276444;
srom_1(66691) <= 7848088;
srom_1(66692) <= 8422267;
srom_1(66693) <= 8996288;
srom_1(66694) <= 9567460;
srom_1(66695) <= 10133104;
srom_1(66696) <= 10690567;
srom_1(66697) <= 11237235;
srom_1(66698) <= 11770545;
srom_1(66699) <= 12287996;
srom_1(66700) <= 12787162;
srom_1(66701) <= 13265701;
srom_1(66702) <= 13721369;
srom_1(66703) <= 14152031;
srom_1(66704) <= 14555666;
srom_1(66705) <= 14930381;
srom_1(66706) <= 15274420;
srom_1(66707) <= 15586169;
srom_1(66708) <= 15864166;
srom_1(66709) <= 16107108;
srom_1(66710) <= 16313855;
srom_1(66711) <= 16483437;
srom_1(66712) <= 16615061;
srom_1(66713) <= 16708107;
srom_1(66714) <= 16762141;
srom_1(66715) <= 16776908;
srom_1(66716) <= 16752339;
srom_1(66717) <= 16688551;
srom_1(66718) <= 16585840;
srom_1(66719) <= 16444691;
srom_1(66720) <= 16265763;
srom_1(66721) <= 16049897;
srom_1(66722) <= 15798104;
srom_1(66723) <= 15511566;
srom_1(66724) <= 15191625;
srom_1(66725) <= 14839783;
srom_1(66726) <= 14457690;
srom_1(66727) <= 14047136;
srom_1(66728) <= 13610047;
srom_1(66729) <= 13148473;
srom_1(66730) <= 12664579;
srom_1(66731) <= 12160633;
srom_1(66732) <= 11638999;
srom_1(66733) <= 11102122;
srom_1(66734) <= 10552521;
srom_1(66735) <= 9992773;
srom_1(66736) <= 9425502;
srom_1(66737) <= 8853369;
srom_1(66738) <= 8279056;
srom_1(66739) <= 7705257;
srom_1(66740) <= 7134663;
srom_1(66741) <= 6569948;
srom_1(66742) <= 6013762;
srom_1(66743) <= 5468713;
srom_1(66744) <= 4937356;
srom_1(66745) <= 4422183;
srom_1(66746) <= 3925609;
srom_1(66747) <= 3449965;
srom_1(66748) <= 2997479;
srom_1(66749) <= 2570274;
srom_1(66750) <= 2170354;
srom_1(66751) <= 1799593;
srom_1(66752) <= 1459730;
srom_1(66753) <= 1152359;
srom_1(66754) <= 878921;
srom_1(66755) <= 640699;
srom_1(66756) <= 438809;
srom_1(66757) <= 274199;
srom_1(66758) <= 147639;
srom_1(66759) <= 59725;
srom_1(66760) <= 10868;
srom_1(66761) <= 1296;
srom_1(66762) <= 31056;
srom_1(66763) <= 100007;
srom_1(66764) <= 207826;
srom_1(66765) <= 354008;
srom_1(66766) <= 537866;
srom_1(66767) <= 758540;
srom_1(66768) <= 1014993;
srom_1(66769) <= 1306024;
srom_1(66770) <= 1630268;
srom_1(66771) <= 1986204;
srom_1(66772) <= 2372162;
srom_1(66773) <= 2786334;
srom_1(66774) <= 3226777;
srom_1(66775) <= 3691426;
srom_1(66776) <= 4178101;
srom_1(66777) <= 4684521;
srom_1(66778) <= 5208310;
srom_1(66779) <= 5747013;
srom_1(66780) <= 6298103;
srom_1(66781) <= 6858997;
srom_1(66782) <= 7427063;
srom_1(66783) <= 7999638;
srom_1(66784) <= 8574038;
srom_1(66785) <= 9147567;
srom_1(66786) <= 9717538;
srom_1(66787) <= 10281277;
srom_1(66788) <= 10836140;
srom_1(66789) <= 11379526;
srom_1(66790) <= 11908887;
srom_1(66791) <= 12421740;
srom_1(66792) <= 12915680;
srom_1(66793) <= 13388391;
srom_1(66794) <= 13837657;
srom_1(66795) <= 14261370;
srom_1(66796) <= 14657543;
srom_1(66797) <= 15024320;
srom_1(66798) <= 15359979;
srom_1(66799) <= 15662947;
srom_1(66800) <= 15931803;
srom_1(66801) <= 16165287;
srom_1(66802) <= 16362303;
srom_1(66803) <= 16521927;
srom_1(66804) <= 16643412;
srom_1(66805) <= 16726187;
srom_1(66806) <= 16769864;
srom_1(66807) <= 16774239;
srom_1(66808) <= 16739291;
srom_1(66809) <= 16665183;
srom_1(66810) <= 16552264;
srom_1(66811) <= 16401062;
srom_1(66812) <= 16212287;
srom_1(66813) <= 15986825;
srom_1(66814) <= 15725731;
srom_1(66815) <= 15430232;
srom_1(66816) <= 15101712;
srom_1(66817) <= 14741711;
srom_1(66818) <= 14351919;
srom_1(66819) <= 13934163;
srom_1(66820) <= 13490402;
srom_1(66821) <= 13022717;
srom_1(66822) <= 12533300;
srom_1(66823) <= 12024448;
srom_1(66824) <= 11498547;
srom_1(66825) <= 10958061;
srom_1(66826) <= 10405527;
srom_1(66827) <= 9843534;
srom_1(66828) <= 9274719;
srom_1(66829) <= 8701749;
srom_1(66830) <= 8127310;
srom_1(66831) <= 7554096;
srom_1(66832) <= 6984796;
srom_1(66833) <= 6422079;
srom_1(66834) <= 5868583;
srom_1(66835) <= 5326905;
srom_1(66836) <= 4799584;
srom_1(66837) <= 4289093;
srom_1(66838) <= 3797827;
srom_1(66839) <= 3328088;
srom_1(66840) <= 2882079;
srom_1(66841) <= 2461893;
srom_1(66842) <= 2069498;
srom_1(66843) <= 1706737;
srom_1(66844) <= 1375309;
srom_1(66845) <= 1076769;
srom_1(66846) <= 812516;
srom_1(66847) <= 583790;
srom_1(66848) <= 391664;
srom_1(66849) <= 237038;
srom_1(66850) <= 120638;
srom_1(66851) <= 43009;
srom_1(66852) <= 4516;
srom_1(66853) <= 5338;
srom_1(66854) <= 45472;
srom_1(66855) <= 124730;
srom_1(66856) <= 242741;
srom_1(66857) <= 398950;
srom_1(66858) <= 592625;
srom_1(66859) <= 822858;
srom_1(66860) <= 1088570;
srom_1(66861) <= 1388514;
srom_1(66862) <= 1721284;
srom_1(66863) <= 2085320;
srom_1(66864) <= 2478913;
srom_1(66865) <= 2900219;
srom_1(66866) <= 3347263;
srom_1(66867) <= 3817946;
srom_1(66868) <= 4310063;
srom_1(66869) <= 4821306;
srom_1(66870) <= 5349277;
srom_1(66871) <= 5891501;
srom_1(66872) <= 6445434;
srom_1(66873) <= 7008480;
srom_1(66874) <= 7577997;
srom_1(66875) <= 8151316;
srom_1(66876) <= 8725747;
srom_1(66877) <= 9298598;
srom_1(66878) <= 9867181;
srom_1(66879) <= 10428831;
srom_1(66880) <= 10980913;
srom_1(66881) <= 11520839;
srom_1(66882) <= 12046077;
srom_1(66883) <= 12554164;
srom_1(66884) <= 13042717;
srom_1(66885) <= 13509445;
srom_1(66886) <= 13952160;
srom_1(66887) <= 14368786;
srom_1(66888) <= 14757368;
srom_1(66889) <= 15116086;
srom_1(66890) <= 15443255;
srom_1(66891) <= 15737343;
srom_1(66892) <= 15996971;
srom_1(66893) <= 16220920;
srom_1(66894) <= 16408140;
srom_1(66895) <= 16557755;
srom_1(66896) <= 16669061;
srom_1(66897) <= 16741538;
srom_1(66898) <= 16774844;
srom_1(66899) <= 16768825;
srom_1(66900) <= 16723508;
srom_1(66901) <= 16639106;
srom_1(66902) <= 16516014;
srom_1(66903) <= 16354810;
srom_1(66904) <= 16156250;
srom_1(66905) <= 15921265;
srom_1(66906) <= 15650957;
srom_1(66907) <= 15346593;
srom_1(66908) <= 15009600;
srom_1(66909) <= 14641559;
srom_1(66910) <= 14244197;
srom_1(66911) <= 13819375;
srom_1(66912) <= 13369086;
srom_1(66913) <= 12895443;
srom_1(66914) <= 12400665;
srom_1(66915) <= 11887073;
srom_1(66916) <= 11357076;
srom_1(66917) <= 10813159;
srom_1(66918) <= 10257872;
srom_1(66919) <= 9693819;
srom_1(66920) <= 9123646;
srom_1(66921) <= 8550026;
srom_1(66922) <= 7975649;
srom_1(66923) <= 7403209;
srom_1(66924) <= 6835389;
srom_1(66925) <= 6274853;
srom_1(66926) <= 5724229;
srom_1(66927) <= 5186100;
srom_1(66928) <= 4662987;
srom_1(66929) <= 4157346;
srom_1(66930) <= 3671547;
srom_1(66931) <= 3207867;
srom_1(66932) <= 2768482;
srom_1(66933) <= 2355451;
srom_1(66934) <= 1970712;
srom_1(66935) <= 1616069;
srom_1(66936) <= 1293184;
srom_1(66937) <= 1003572;
srom_1(66938) <= 748591;
srom_1(66939) <= 529437;
srom_1(66940) <= 347137;
srom_1(66941) <= 202547;
srom_1(66942) <= 96344;
srom_1(66943) <= 29025;
srom_1(66944) <= 908;
srom_1(66945) <= 12124;
srom_1(66946) <= 62620;
srom_1(66947) <= 152159;
srom_1(66948) <= 280322;
srom_1(66949) <= 446507;
srom_1(66950) <= 649936;
srom_1(66951) <= 889654;
srom_1(66952) <= 1164537;
srom_1(66953) <= 1473296;
srom_1(66954) <= 1814484;
srom_1(66955) <= 2186499;
srom_1(66956) <= 2587599;
srom_1(66957) <= 3015901;
srom_1(66958) <= 3469398;
srom_1(66959) <= 3945963;
srom_1(66960) <= 4443361;
srom_1(66961) <= 4959260;
srom_1(66962) <= 5491240;
srom_1(66963) <= 6036806;
srom_1(66964) <= 6593401;
srom_1(66965) <= 7158415;
srom_1(66966) <= 7729197;
srom_1(66967) <= 8303071;
srom_1(66968) <= 8877347;
srom_1(66969) <= 9449330;
srom_1(66970) <= 10016340;
srom_1(66971) <= 10575716;
srom_1(66972) <= 11124837;
srom_1(66973) <= 11661126;
srom_1(66974) <= 12182069;
srom_1(66975) <= 12685224;
srom_1(66976) <= 13168230;
srom_1(66977) <= 13628823;
srom_1(66978) <= 14064842;
srom_1(66979) <= 14474244;
srom_1(66980) <= 14855108;
srom_1(66981) <= 15205649;
srom_1(66982) <= 15524222;
srom_1(66983) <= 15809334;
srom_1(66984) <= 16059647;
srom_1(66985) <= 16273989;
srom_1(66986) <= 16451353;
srom_1(66987) <= 16590908;
srom_1(66988) <= 16691999;
srom_1(66989) <= 16754153;
srom_1(66990) <= 16777079;
srom_1(66991) <= 16760667;
srom_1(66992) <= 16704997;
srom_1(66993) <= 16610328;
srom_1(66994) <= 16477104;
srom_1(66995) <= 16305951;
srom_1(66996) <= 16097670;
srom_1(66997) <= 15853239;
srom_1(66998) <= 15573804;
srom_1(66999) <= 15260675;
srom_1(67000) <= 14915321;
srom_1(67001) <= 14539360;
srom_1(67002) <= 14134557;
srom_1(67003) <= 13702809;
srom_1(67004) <= 13246140;
srom_1(67005) <= 12766693;
srom_1(67006) <= 12266716;
srom_1(67007) <= 11748553;
srom_1(67008) <= 11214634;
srom_1(67009) <= 10667462;
srom_1(67010) <= 10109605;
srom_1(67011) <= 9543677;
srom_1(67012) <= 8972332;
srom_1(67013) <= 8398251;
srom_1(67014) <= 7824124;
srom_1(67015) <= 7252644;
srom_1(67016) <= 6686491;
srom_1(67017) <= 6128319;
srom_1(67018) <= 5580747;
srom_1(67019) <= 5046343;
srom_1(67020) <= 4527611;
srom_1(67021) <= 4026984;
srom_1(67022) <= 3546811;
srom_1(67023) <= 3089343;
srom_1(67024) <= 2656724;
srom_1(67025) <= 2250985;
srom_1(67026) <= 1874027;
srom_1(67027) <= 1527617;
srom_1(67028) <= 1213382;
srom_1(67029) <= 932794;
srom_1(67030) <= 687168;
srom_1(67031) <= 477657;
srom_1(67032) <= 305243;
srom_1(67033) <= 170735;
srom_1(67034) <= 74764;
srom_1(67035) <= 17779;
srom_1(67036) <= 47;
srom_1(67037) <= 21653;
srom_1(67038) <= 82494;
srom_1(67039) <= 182285;
srom_1(67040) <= 320558;
srom_1(67041) <= 496665;
srom_1(67042) <= 709781;
srom_1(67043) <= 958904;
srom_1(67044) <= 1242869;
srom_1(67045) <= 1560342;
srom_1(67046) <= 1909835;
srom_1(67047) <= 2289710;
srom_1(67048) <= 2698184;
srom_1(67049) <= 3133342;
srom_1(67050) <= 3593145;
srom_1(67051) <= 4075435;
srom_1(67052) <= 4577950;
srom_1(67053) <= 5098336;
srom_1(67054) <= 5634150;
srom_1(67055) <= 6182881;
srom_1(67056) <= 6741956;
srom_1(67057) <= 7308752;
srom_1(67058) <= 7880612;
srom_1(67059) <= 8454854;
srom_1(67060) <= 9028786;
srom_1(67061) <= 9599715;
srom_1(67062) <= 10164966;
srom_1(67063) <= 10721886;
srom_1(67064) <= 11267865;
srom_1(67065) <= 11800341;
srom_1(67066) <= 12316820;
srom_1(67067) <= 12814877;
srom_1(67068) <= 13292178;
srom_1(67069) <= 13746484;
srom_1(67070) <= 14175666;
srom_1(67071) <= 14577710;
srom_1(67072) <= 14950731;
srom_1(67073) <= 15292980;
srom_1(67074) <= 15602853;
srom_1(67075) <= 15878895;
srom_1(67076) <= 16119812;
srom_1(67077) <= 16324476;
srom_1(67078) <= 16491925;
srom_1(67079) <= 16621375;
srom_1(67080) <= 16712219;
srom_1(67081) <= 16764030;
srom_1(67082) <= 16776566;
srom_1(67083) <= 16749769;
srom_1(67084) <= 16683762;
srom_1(67085) <= 16578857;
srom_1(67086) <= 16435546;
srom_1(67087) <= 16254499;
srom_1(67088) <= 16036566;
srom_1(67089) <= 15782770;
srom_1(67090) <= 15494299;
srom_1(67091) <= 15172508;
srom_1(67092) <= 14818905;
srom_1(67093) <= 14435147;
srom_1(67094) <= 14023036;
srom_1(67095) <= 13584502;
srom_1(67096) <= 13121604;
srom_1(67097) <= 12636510;
srom_1(67098) <= 12131497;
srom_1(67099) <= 11608932;
srom_1(67100) <= 11071266;
srom_1(67101) <= 10521020;
srom_1(67102) <= 9960775;
srom_1(67103) <= 9393156;
srom_1(67104) <= 8820828;
srom_1(67105) <= 8246472;
srom_1(67106) <= 7672783;
srom_1(67107) <= 7102451;
srom_1(67108) <= 6538149;
srom_1(67109) <= 5982526;
srom_1(67110) <= 5438185;
srom_1(67111) <= 4907680;
srom_1(67112) <= 4393498;
srom_1(67113) <= 3898050;
srom_1(67114) <= 3423661;
srom_1(67115) <= 2972553;
srom_1(67116) <= 2546843;
srom_1(67117) <= 2148528;
srom_1(67118) <= 1779474;
srom_1(67119) <= 1441413;
srom_1(67120) <= 1135929;
srom_1(67121) <= 864456;
srom_1(67122) <= 628266;
srom_1(67123) <= 428467;
srom_1(67124) <= 265996;
srom_1(67125) <= 141615;
srom_1(67126) <= 55906;
srom_1(67127) <= 9272;
srom_1(67128) <= 1932;
srom_1(67129) <= 33921;
srom_1(67130) <= 105086;
srom_1(67131) <= 215097;
srom_1(67132) <= 363435;
srom_1(67133) <= 549407;
srom_1(67134) <= 772139;
srom_1(67135) <= 1030587;
srom_1(67136) <= 1323540;
srom_1(67137) <= 1649623;
srom_1(67138) <= 2007308;
srom_1(67139) <= 2394917;
srom_1(67140) <= 2810632;
srom_1(67141) <= 3252504;
srom_1(67142) <= 3718461;
srom_1(67143) <= 4206318;
srom_1(67144) <= 4713787;
srom_1(67145) <= 5238489;
srom_1(67146) <= 5777963;
srom_1(67147) <= 6329679;
srom_1(67148) <= 6891050;
srom_1(67149) <= 7459443;
srom_1(67150) <= 8032194;
srom_1(67151) <= 8606616;
srom_1(67152) <= 9180016;
srom_1(67153) <= 9749704;
srom_1(67154) <= 10313010;
srom_1(67155) <= 10867292;
srom_1(67156) <= 11409950;
srom_1(67157) <= 11938440;
srom_1(67158) <= 12450284;
srom_1(67159) <= 12943081;
srom_1(67160) <= 13414521;
srom_1(67161) <= 13862392;
srom_1(67162) <= 14284595;
srom_1(67163) <= 14679150;
srom_1(67164) <= 15044206;
srom_1(67165) <= 15378052;
srom_1(67166) <= 15679121;
srom_1(67167) <= 15946003;
srom_1(67168) <= 16177446;
srom_1(67169) <= 16372365;
srom_1(67170) <= 16529844;
srom_1(67171) <= 16649147;
srom_1(67172) <= 16729713;
srom_1(67173) <= 16771165;
srom_1(67174) <= 16773308;
srom_1(67175) <= 16736133;
srom_1(67176) <= 16659813;
srom_1(67177) <= 16544706;
srom_1(67178) <= 16391353;
srom_1(67179) <= 16200472;
srom_1(67180) <= 15972958;
srom_1(67181) <= 15709879;
srom_1(67182) <= 15412468;
srom_1(67183) <= 15082120;
srom_1(67184) <= 14720383;
srom_1(67185) <= 14328955;
srom_1(67186) <= 13909670;
srom_1(67187) <= 13464495;
srom_1(67188) <= 12995518;
srom_1(67189) <= 12504937;
srom_1(67190) <= 11995053;
srom_1(67191) <= 11468258;
srom_1(67192) <= 10927020;
srom_1(67193) <= 10373880;
srom_1(67194) <= 9811429;
srom_1(67195) <= 9242307;
srom_1(67196) <= 8669181;
srom_1(67197) <= 8094740;
srom_1(67198) <= 7521677;
srom_1(67199) <= 6952679;
srom_1(67200) <= 6390414;
srom_1(67201) <= 5837520;
srom_1(67202) <= 5296588;
srom_1(67203) <= 4770157;
srom_1(67204) <= 4260693;
srom_1(67205) <= 3770587;
srom_1(67206) <= 3302136;
srom_1(67207) <= 2857537;
srom_1(67208) <= 2438875;
srom_1(67209) <= 2048114;
srom_1(67210) <= 1687085;
srom_1(67211) <= 1357482;
srom_1(67212) <= 1060851;
srom_1(67213) <= 798582;
srom_1(67214) <= 571905;
srom_1(67215) <= 381883;
srom_1(67216) <= 229408;
srom_1(67217) <= 115194;
srom_1(67218) <= 39776;
srom_1(67219) <= 3510;
srom_1(67220) <= 6563;
srom_1(67221) <= 48924;
srom_1(67222) <= 130391;
srom_1(67223) <= 250585;
srom_1(67224) <= 408940;
srom_1(67225) <= 604715;
srom_1(67226) <= 836991;
srom_1(67227) <= 1104679;
srom_1(67228) <= 1406524;
srom_1(67229) <= 1741111;
srom_1(67230) <= 2106870;
srom_1(67231) <= 2502086;
srom_1(67232) <= 2924906;
srom_1(67233) <= 3373347;
srom_1(67234) <= 3845306;
srom_1(67235) <= 4338571;
srom_1(67236) <= 4850827;
srom_1(67237) <= 5379674;
srom_1(67238) <= 5922630;
srom_1(67239) <= 6477150;
srom_1(67240) <= 7040634;
srom_1(67241) <= 7610439;
srom_1(67242) <= 8183892;
srom_1(67243) <= 8758306;
srom_1(67244) <= 9330986;
srom_1(67245) <= 9899247;
srom_1(67246) <= 10460424;
srom_1(67247) <= 11011886;
srom_1(67248) <= 11551046;
srom_1(67249) <= 12075376;
srom_1(67250) <= 12582418;
srom_1(67251) <= 13069794;
srom_1(67252) <= 13535218;
srom_1(67253) <= 13976508;
srom_1(67254) <= 14391594;
srom_1(67255) <= 14778530;
srom_1(67256) <= 15135501;
srom_1(67257) <= 15460834;
srom_1(67258) <= 15753003;
srom_1(67259) <= 16010638;
srom_1(67260) <= 16232530;
srom_1(67261) <= 16417640;
srom_1(67262) <= 16565098;
srom_1(67263) <= 16674215;
srom_1(67264) <= 16744477;
srom_1(67265) <= 16775555;
srom_1(67266) <= 16767305;
srom_1(67267) <= 16719764;
srom_1(67268) <= 16633155;
srom_1(67269) <= 16507884;
srom_1(67270) <= 16344540;
srom_1(67271) <= 16143887;
srom_1(67272) <= 15906867;
srom_1(67273) <= 15634592;
srom_1(67274) <= 15328337;
srom_1(67275) <= 14989540;
srom_1(67276) <= 14619789;
srom_1(67277) <= 14220818;
srom_1(67278) <= 13794497;
srom_1(67279) <= 13342826;
srom_1(67280) <= 12867924;
srom_1(67281) <= 12372016;
srom_1(67282) <= 11857428;
srom_1(67283) <= 11326575;
srom_1(67284) <= 10781944;
srom_1(67285) <= 10226089;
srom_1(67286) <= 9661619;
srom_1(67287) <= 9091178;
srom_1(67288) <= 8517443;
srom_1(67289) <= 7943104;
srom_1(67290) <= 7370854;
srom_1(67291) <= 6803377;
srom_1(67292) <= 6243333;
srom_1(67293) <= 5693349;
srom_1(67294) <= 5156004;
srom_1(67295) <= 4633818;
srom_1(67296) <= 4129240;
srom_1(67297) <= 3644635;
srom_1(67298) <= 3182276;
srom_1(67299) <= 2744331;
srom_1(67300) <= 2332855;
srom_1(67301) <= 1949776;
srom_1(67302) <= 1596890;
srom_1(67303) <= 1275854;
srom_1(67304) <= 988172;
srom_1(67305) <= 735192;
srom_1(67306) <= 518103;
srom_1(67307) <= 337921;
srom_1(67308) <= 195491;
srom_1(67309) <= 91481;
srom_1(67310) <= 26380;
srom_1(67311) <= 492;
srom_1(67312) <= 13939;
srom_1(67313) <= 66657;
srom_1(67314) <= 158400;
srom_1(67315) <= 288737;
srom_1(67316) <= 457057;
srom_1(67317) <= 662571;
srom_1(67318) <= 904316;
srom_1(67319) <= 1181156;
srom_1(67320) <= 1491795;
srom_1(67321) <= 1834775;
srom_1(67322) <= 2208488;
srom_1(67323) <= 2611182;
srom_1(67324) <= 3040969;
srom_1(67325) <= 3495832;
srom_1(67326) <= 3973639;
srom_1(67327) <= 4472150;
srom_1(67328) <= 4989026;
srom_1(67329) <= 5521844;
srom_1(67330) <= 6068105;
srom_1(67331) <= 6625248;
srom_1(67332) <= 7190659;
srom_1(67333) <= 7761689;
srom_1(67334) <= 8335658;
srom_1(67335) <= 8909875;
srom_1(67336) <= 9481648;
srom_1(67337) <= 10048296;
srom_1(67338) <= 10607160;
srom_1(67339) <= 11155621;
srom_1(67340) <= 11691107;
srom_1(67341) <= 12211106;
srom_1(67342) <= 12713180;
srom_1(67343) <= 13194974;
srom_1(67344) <= 13654230;
srom_1(67345) <= 14088794;
srom_1(67346) <= 14496627;
srom_1(67347) <= 14875818;
srom_1(67348) <= 15224588;
srom_1(67349) <= 15541302;
srom_1(67350) <= 15824474;
srom_1(67351) <= 16072777;
srom_1(67352) <= 16285046;
srom_1(67353) <= 16460286;
srom_1(67354) <= 16597676;
srom_1(67355) <= 16696570;
srom_1(67356) <= 16756505;
srom_1(67357) <= 16777200;
srom_1(67358) <= 16758558;
srom_1(67359) <= 16700667;
srom_1(67360) <= 16603798;
srom_1(67361) <= 16468404;
srom_1(67362) <= 16295122;
srom_1(67363) <= 16084764;
srom_1(67364) <= 15838315;
srom_1(67365) <= 15556932;
srom_1(67366) <= 15241935;
srom_1(67367) <= 14894800;
srom_1(67368) <= 14517155;
srom_1(67369) <= 14110771;
srom_1(67370) <= 13677554;
srom_1(67371) <= 13219535;
srom_1(67372) <= 12738863;
srom_1(67373) <= 12237790;
srom_1(67374) <= 11718668;
srom_1(67375) <= 11183930;
srom_1(67376) <= 10636083;
srom_1(67377) <= 10077697;
srom_1(67378) <= 9511391;
srom_1(67379) <= 8939819;
srom_1(67380) <= 8365663;
srom_1(67381) <= 7791614;
srom_1(67382) <= 7220365;
srom_1(67383) <= 6654594;
srom_1(67384) <= 6096954;
srom_1(67385) <= 5550061;
srom_1(67386) <= 5016478;
srom_1(67387) <= 4498709;
srom_1(67388) <= 3999181;
srom_1(67389) <= 3520236;
srom_1(67390) <= 3064121;
srom_1(67391) <= 2632974;
srom_1(67392) <= 2228817;
srom_1(67393) <= 1853546;
srom_1(67394) <= 1508919;
srom_1(67395) <= 1196554;
srom_1(67396) <= 917915;
srom_1(67397) <= 674309;
srom_1(67398) <= 466877;
srom_1(67399) <= 296594;
srom_1(67400) <= 164256;
srom_1(67401) <= 70485;
srom_1(67402) <= 15721;
srom_1(67403) <= 220;
srom_1(67404) <= 24056;
srom_1(67405) <= 87115;
srom_1(67406) <= 189103;
srom_1(67407) <= 329541;
srom_1(67408) <= 507771;
srom_1(67409) <= 722957;
srom_1(67410) <= 974090;
srom_1(67411) <= 1259992;
srom_1(67412) <= 1579323;
srom_1(67413) <= 1930584;
srom_1(67414) <= 2312130;
srom_1(67415) <= 2722170;
srom_1(67416) <= 3158782;
srom_1(67417) <= 3619919;
srom_1(67418) <= 4103417;
srom_1(67419) <= 4607011;
srom_1(67420) <= 5128337;
srom_1(67421) <= 5664952;
srom_1(67422) <= 6214339;
srom_1(67423) <= 6773922;
srom_1(67424) <= 7341077;
srom_1(67425) <= 7913144;
srom_1(67426) <= 8487441;
srom_1(67427) <= 9061274;
srom_1(67428) <= 9631953;
srom_1(67429) <= 10196801;
srom_1(67430) <= 10753170;
srom_1(67431) <= 11298451;
srom_1(67432) <= 11830087;
srom_1(67433) <= 12345584;
srom_1(67434) <= 12842525;
srom_1(67435) <= 13318581;
srom_1(67436) <= 13771519;
srom_1(67437) <= 14199214;
srom_1(67438) <= 14599661;
srom_1(67439) <= 14970982;
srom_1(67440) <= 15311436;
srom_1(67441) <= 15619427;
srom_1(67442) <= 15893510;
srom_1(67443) <= 16132400;
srom_1(67444) <= 16334977;
srom_1(67445) <= 16500290;
srom_1(67446) <= 16627565;
srom_1(67447) <= 16716205;
srom_1(67448) <= 16765793;
srom_1(67449) <= 16776098;
srom_1(67450) <= 16747072;
srom_1(67451) <= 16678849;
srom_1(67452) <= 16571751;
srom_1(67453) <= 16426279;
srom_1(67454) <= 16243116;
srom_1(67455) <= 16023120;
srom_1(67456) <= 15767324;
srom_1(67457) <= 15476926;
srom_1(67458) <= 15153288;
srom_1(67459) <= 14797929;
srom_1(67460) <= 14412514;
srom_1(67461) <= 13998851;
srom_1(67462) <= 13558879;
srom_1(67463) <= 13094663;
srom_1(67464) <= 12608378;
srom_1(67465) <= 12102305;
srom_1(67466) <= 11578817;
srom_1(67467) <= 11040370;
srom_1(67468) <= 10489487;
srom_1(67469) <= 9928752;
srom_1(67470) <= 9360796;
srom_1(67471) <= 8788280;
srom_1(67472) <= 8213890;
srom_1(67473) <= 7640319;
srom_1(67474) <= 7070258;
srom_1(67475) <= 6506378;
srom_1(67476) <= 5951325;
srom_1(67477) <= 5407702;
srom_1(67478) <= 4878056;
srom_1(67479) <= 4364873;
srom_1(67480) <= 3870559;
srom_1(67481) <= 3397431;
srom_1(67482) <= 2947709;
srom_1(67483) <= 2523501;
srom_1(67484) <= 2126796;
srom_1(67485) <= 1759455;
srom_1(67486) <= 1423200;
srom_1(67487) <= 1119609;
srom_1(67488) <= 850105;
srom_1(67489) <= 615951;
srom_1(67490) <= 418245;
srom_1(67491) <= 257916;
srom_1(67492) <= 135714;
srom_1(67493) <= 52213;
srom_1(67494) <= 7804;
srom_1(67495) <= 2695;
srom_1(67496) <= 36911;
srom_1(67497) <= 110291;
srom_1(67498) <= 222491;
srom_1(67499) <= 372984;
srom_1(67500) <= 561066;
srom_1(67501) <= 785853;
srom_1(67502) <= 1046292;
srom_1(67503) <= 1341162;
srom_1(67504) <= 1669080;
srom_1(67505) <= 2028508;
srom_1(67506) <= 2417761;
srom_1(67507) <= 2835013;
srom_1(67508) <= 3278308;
srom_1(67509) <= 3745567;
srom_1(67510) <= 4234598;
srom_1(67511) <= 4743110;
srom_1(67512) <= 5268716;
srom_1(67513) <= 5808952;
srom_1(67514) <= 6361285;
srom_1(67515) <= 6923125;
srom_1(67516) <= 7491837;
srom_1(67517) <= 8064755;
srom_1(67518) <= 8639191;
srom_1(67519) <= 9212452;
srom_1(67520) <= 9781850;
srom_1(67521) <= 10344714;
srom_1(67522) <= 10898406;
srom_1(67523) <= 11440328;
srom_1(67524) <= 11967939;
srom_1(67525) <= 12478766;
srom_1(67526) <= 12970413;
srom_1(67527) <= 13440574;
srom_1(67528) <= 13887045;
srom_1(67529) <= 14307731;
srom_1(67530) <= 14700661;
srom_1(67531) <= 15063991;
srom_1(67532) <= 15396019;
srom_1(67533) <= 15695186;
srom_1(67534) <= 15960090;
srom_1(67535) <= 16189488;
srom_1(67536) <= 16382306;
srom_1(67537) <= 16537638;
srom_1(67538) <= 16654757;
srom_1(67539) <= 16733113;
srom_1(67540) <= 16772339;
srom_1(67541) <= 16772251;
srom_1(67542) <= 16732848;
srom_1(67543) <= 16654317;
srom_1(67544) <= 16537025;
srom_1(67545) <= 16381522;
srom_1(67546) <= 16188538;
srom_1(67547) <= 15958977;
srom_1(67548) <= 15693917;
srom_1(67549) <= 15394599;
srom_1(67550) <= 15062427;
srom_1(67551) <= 14698960;
srom_1(67552) <= 14305901;
srom_1(67553) <= 13885094;
srom_1(67554) <= 13438512;
srom_1(67555) <= 12968249;
srom_1(67556) <= 12476511;
srom_1(67557) <= 11965604;
srom_1(67558) <= 11437922;
srom_1(67559) <= 10895941;
srom_1(67560) <= 10342203;
srom_1(67561) <= 9779303;
srom_1(67562) <= 9209882;
srom_1(67563) <= 8636610;
srom_1(67564) <= 8062174;
srom_1(67565) <= 7489270;
srom_1(67566) <= 6920583;
srom_1(67567) <= 6358779;
srom_1(67568) <= 5806495;
srom_1(67569) <= 5266319;
srom_1(67570) <= 4740784;
srom_1(67571) <= 4232355;
srom_1(67572) <= 3743416;
srom_1(67573) <= 3276260;
srom_1(67574) <= 2833078;
srom_1(67575) <= 2415948;
srom_1(67576) <= 2026825;
srom_1(67577) <= 1667535;
srom_1(67578) <= 1339762;
srom_1(67579) <= 1045044;
srom_1(67580) <= 784762;
srom_1(67581) <= 560137;
srom_1(67582) <= 372223;
srom_1(67583) <= 221900;
srom_1(67584) <= 109874;
srom_1(67585) <= 36670;
srom_1(67586) <= 2630;
srom_1(67587) <= 7916;
srom_1(67588) <= 52501;
srom_1(67589) <= 136177;
srom_1(67590) <= 258552;
srom_1(67591) <= 419051;
srom_1(67592) <= 616922;
srom_1(67593) <= 851238;
srom_1(67594) <= 1120898;
srom_1(67595) <= 1424640;
srom_1(67596) <= 1761038;
srom_1(67597) <= 2128515;
srom_1(67598) <= 2525347;
srom_1(67599) <= 2949675;
srom_1(67600) <= 3399507;
srom_1(67601) <= 3872735;
srom_1(67602) <= 4367140;
srom_1(67603) <= 4880402;
srom_1(67604) <= 5410116;
srom_1(67605) <= 5953797;
srom_1(67606) <= 6508895;
srom_1(67607) <= 7072808;
srom_1(67608) <= 7642892;
srom_1(67609) <= 8216472;
srom_1(67610) <= 8790859;
srom_1(67611) <= 9363361;
srom_1(67612) <= 9931291;
srom_1(67613) <= 10491987;
srom_1(67614) <= 11042819;
srom_1(67615) <= 11581206;
srom_1(67616) <= 12104620;
srom_1(67617) <= 12610610;
srom_1(67618) <= 13096800;
srom_1(67619) <= 13560913;
srom_1(67620) <= 14000771;
srom_1(67621) <= 14414311;
srom_1(67622) <= 14799595;
srom_1(67623) <= 15154815;
srom_1(67624) <= 15478306;
srom_1(67625) <= 15768552;
srom_1(67626) <= 16024190;
srom_1(67627) <= 16244022;
srom_1(67628) <= 16427018;
srom_1(67629) <= 16572319;
srom_1(67630) <= 16679243;
srom_1(67631) <= 16747290;
srom_1(67632) <= 16776140;
srom_1(67633) <= 16765658;
srom_1(67634) <= 16715893;
srom_1(67635) <= 16627079;
srom_1(67636) <= 16499632;
srom_1(67637) <= 16334149;
srom_1(67638) <= 16131407;
srom_1(67639) <= 15892356;
srom_1(67640) <= 15618118;
srom_1(67641) <= 15309978;
srom_1(67642) <= 14969381;
srom_1(67643) <= 14597925;
srom_1(67644) <= 14197351;
srom_1(67645) <= 13769538;
srom_1(67646) <= 13316492;
srom_1(67647) <= 12840337;
srom_1(67648) <= 12343306;
srom_1(67649) <= 11827731;
srom_1(67650) <= 11296029;
srom_1(67651) <= 10750692;
srom_1(67652) <= 10194279;
srom_1(67653) <= 9629399;
srom_1(67654) <= 9058700;
srom_1(67655) <= 8484858;
srom_1(67656) <= 7910566;
srom_1(67657) <= 7338515;
srom_1(67658) <= 6771388;
srom_1(67659) <= 6211845;
srom_1(67660) <= 5662509;
srom_1(67661) <= 5125958;
srom_1(67662) <= 4604706;
srom_1(67663) <= 4101197;
srom_1(67664) <= 3617794;
srom_1(67665) <= 3156763;
srom_1(67666) <= 2720266;
srom_1(67667) <= 2310350;
srom_1(67668) <= 1928937;
srom_1(67669) <= 1577815;
srom_1(67670) <= 1258631;
srom_1(67671) <= 972883;
srom_1(67672) <= 721909;
srom_1(67673) <= 506887;
srom_1(67674) <= 328825;
srom_1(67675) <= 188558;
srom_1(67676) <= 86744;
srom_1(67677) <= 23861;
srom_1(67678) <= 202;
srom_1(67679) <= 15880;
srom_1(67680) <= 70820;
srom_1(67681) <= 164765;
srom_1(67682) <= 297275;
srom_1(67683) <= 467727;
srom_1(67684) <= 675324;
srom_1(67685) <= 919090;
srom_1(67686) <= 1197884;
srom_1(67687) <= 1510397;
srom_1(67688) <= 1855165;
srom_1(67689) <= 2230570;
srom_1(67690) <= 2634853;
srom_1(67691) <= 3066117;
srom_1(67692) <= 3522339;
srom_1(67693) <= 4001382;
srom_1(67694) <= 4500997;
srom_1(67695) <= 5018843;
srom_1(67696) <= 5552491;
srom_1(67697) <= 6099438;
srom_1(67698) <= 6657120;
srom_1(67699) <= 7222922;
srom_1(67700) <= 7794190;
srom_1(67701) <= 8368245;
srom_1(67702) <= 8942396;
srom_1(67703) <= 9513950;
srom_1(67704) <= 10080227;
srom_1(67705) <= 10638571;
srom_1(67706) <= 11186364;
srom_1(67707) <= 11721038;
srom_1(67708) <= 12240085;
srom_1(67709) <= 12741071;
srom_1(67710) <= 13221646;
srom_1(67711) <= 13679558;
srom_1(67712) <= 14112659;
srom_1(67713) <= 14518918;
srom_1(67714) <= 14896429;
srom_1(67715) <= 15243424;
srom_1(67716) <= 15558273;
srom_1(67717) <= 15839502;
srom_1(67718) <= 16085791;
srom_1(67719) <= 16295985;
srom_1(67720) <= 16469098;
srom_1(67721) <= 16604320;
srom_1(67722) <= 16701015;
srom_1(67723) <= 16758730;
srom_1(67724) <= 16777195;
srom_1(67725) <= 16756323;
srom_1(67726) <= 16696212;
srom_1(67727) <= 16597144;
srom_1(67728) <= 16459583;
srom_1(67729) <= 16284174;
srom_1(67730) <= 16071741;
srom_1(67731) <= 15823278;
srom_1(67732) <= 15539952;
srom_1(67733) <= 15223091;
srom_1(67734) <= 14874180;
srom_1(67735) <= 14494857;
srom_1(67736) <= 14086899;
srom_1(67737) <= 13652220;
srom_1(67738) <= 13192858;
srom_1(67739) <= 12710967;
srom_1(67740) <= 12208807;
srom_1(67741) <= 11688733;
srom_1(67742) <= 11153183;
srom_1(67743) <= 10604670;
srom_1(67744) <= 10045764;
srom_1(67745) <= 9479088;
srom_1(67746) <= 8907298;
srom_1(67747) <= 8333075;
srom_1(67748) <= 7759113;
srom_1(67749) <= 7188103;
srom_1(67750) <= 6622723;
srom_1(67751) <= 6065623;
srom_1(67752) <= 5519417;
srom_1(67753) <= 4986665;
srom_1(67754) <= 4469866;
srom_1(67755) <= 3971443;
srom_1(67756) <= 3493734;
srom_1(67757) <= 3038979;
srom_1(67758) <= 2609310;
srom_1(67759) <= 2206742;
srom_1(67760) <= 1833163;
srom_1(67761) <= 1490325;
srom_1(67762) <= 1179835;
srom_1(67763) <= 903150;
srom_1(67764) <= 661566;
srom_1(67765) <= 456217;
srom_1(67766) <= 288066;
srom_1(67767) <= 157901;
srom_1(67768) <= 66333;
srom_1(67769) <= 13790;
srom_1(67770) <= 520;
srom_1(67771) <= 26585;
srom_1(67772) <= 91862;
srom_1(67773) <= 196045;
srom_1(67774) <= 338647;
srom_1(67775) <= 518997;
srom_1(67776) <= 736250;
srom_1(67777) <= 989388;
srom_1(67778) <= 1277223;
srom_1(67779) <= 1598407;
srom_1(67780) <= 1951431;
srom_1(67781) <= 2334642;
srom_1(67782) <= 2746242;
srom_1(67783) <= 3184301;
srom_1(67784) <= 3646765;
srom_1(67785) <= 4131465;
srom_1(67786) <= 4636128;
srom_1(67787) <= 5158387;
srom_1(67788) <= 5695795;
srom_1(67789) <= 6245830;
srom_1(67790) <= 6805913;
srom_1(67791) <= 7373417;
srom_1(67792) <= 7945683;
srom_1(67793) <= 8520025;
srom_1(67794) <= 9093752;
srom_1(67795) <= 9664171;
srom_1(67796) <= 10228609;
srom_1(67797) <= 10784419;
srom_1(67798) <= 11328993;
srom_1(67799) <= 11859780;
srom_1(67800) <= 12374288;
srom_1(67801) <= 12870107;
srom_1(67802) <= 13344910;
srom_1(67803) <= 13796472;
srom_1(67804) <= 14222674;
srom_1(67805) <= 14621518;
srom_1(67806) <= 14991134;
srom_1(67807) <= 15329788;
srom_1(67808) <= 15635893;
srom_1(67809) <= 15908012;
srom_1(67810) <= 16144871;
srom_1(67811) <= 16345358;
srom_1(67812) <= 16508533;
srom_1(67813) <= 16633631;
srom_1(67814) <= 16720065;
srom_1(67815) <= 16767430;
srom_1(67816) <= 16775504;
srom_1(67817) <= 16744248;
srom_1(67818) <= 16673811;
srom_1(67819) <= 16564521;
srom_1(67820) <= 16416891;
srom_1(67821) <= 16231614;
srom_1(67822) <= 16009559;
srom_1(67823) <= 15751766;
srom_1(67824) <= 15459445;
srom_1(67825) <= 15133966;
srom_1(67826) <= 14776856;
srom_1(67827) <= 14389790;
srom_1(67828) <= 13974581;
srom_1(67829) <= 13533178;
srom_1(67830) <= 13067651;
srom_1(67831) <= 12580182;
srom_1(67832) <= 12073057;
srom_1(67833) <= 11548654;
srom_1(67834) <= 11009433;
srom_1(67835) <= 10457922;
srom_1(67836) <= 9896707;
srom_1(67837) <= 9328420;
srom_1(67838) <= 8755726;
srom_1(67839) <= 8181311;
srom_1(67840) <= 7607867;
srom_1(67841) <= 7038085;
srom_1(67842) <= 6474636;
srom_1(67843) <= 5920162;
srom_1(67844) <= 5377263;
srom_1(67845) <= 4848486;
srom_1(67846) <= 4336310;
srom_1(67847) <= 3843136;
srom_1(67848) <= 3371277;
srom_1(67849) <= 2922946;
srom_1(67850) <= 2500246;
srom_1(67851) <= 2105158;
srom_1(67852) <= 1739536;
srom_1(67853) <= 1405093;
srom_1(67854) <= 1103399;
srom_1(67855) <= 835867;
srom_1(67856) <= 603753;
srom_1(67857) <= 408144;
srom_1(67858) <= 249959;
srom_1(67859) <= 129938;
srom_1(67860) <= 48646;
srom_1(67861) <= 6462;
srom_1(67862) <= 3585;
srom_1(67863) <= 40028;
srom_1(67864) <= 115620;
srom_1(67865) <= 230008;
srom_1(67866) <= 382654;
srom_1(67867) <= 572842;
srom_1(67868) <= 799682;
srom_1(67869) <= 1062108;
srom_1(67870) <= 1358891;
srom_1(67871) <= 1688639;
srom_1(67872) <= 2049805;
srom_1(67873) <= 2440696;
srom_1(67874) <= 2859479;
srom_1(67875) <= 3304189;
srom_1(67876) <= 3772743;
srom_1(67877) <= 4262941;
srom_1(67878) <= 4772487;
srom_1(67879) <= 5298989;
srom_1(67880) <= 5839980;
srom_1(67881) <= 6392922;
srom_1(67882) <= 6955223;
srom_1(67883) <= 7524245;
srom_1(67884) <= 8097321;
srom_1(67885) <= 8671762;
srom_1(67886) <= 9244876;
srom_1(67887) <= 9813974;
srom_1(67888) <= 10376389;
srom_1(67889) <= 10929482;
srom_1(67890) <= 11470660;
srom_1(67891) <= 11997385;
srom_1(67892) <= 12507187;
srom_1(67893) <= 12997676;
srom_1(67894) <= 13466551;
srom_1(67895) <= 13911614;
srom_1(67896) <= 14330778;
srom_1(67897) <= 14722077;
srom_1(67898) <= 15083676;
srom_1(67899) <= 15413880;
srom_1(67900) <= 15711140;
srom_1(67901) <= 15974061;
srom_1(67902) <= 16201412;
srom_1(67903) <= 16392127;
srom_1(67904) <= 16545309;
srom_1(67905) <= 16660243;
srom_1(67906) <= 16736387;
srom_1(67907) <= 16773387;
srom_1(67908) <= 16771067;
srom_1(67909) <= 16729438;
srom_1(67910) <= 16648697;
srom_1(67911) <= 16529221;
srom_1(67912) <= 16371572;
srom_1(67913) <= 16176487;
srom_1(67914) <= 15944882;
srom_1(67915) <= 15677844;
srom_1(67916) <= 15376623;
srom_1(67917) <= 15042634;
srom_1(67918) <= 14677441;
srom_1(67919) <= 14282758;
srom_1(67920) <= 13860435;
srom_1(67921) <= 13412453;
srom_1(67922) <= 12940912;
srom_1(67923) <= 12448024;
srom_1(67924) <= 11936100;
srom_1(67925) <= 11407541;
srom_1(67926) <= 10864824;
srom_1(67927) <= 10310496;
srom_1(67928) <= 9747156;
srom_1(67929) <= 9177445;
srom_1(67930) <= 8604034;
srom_1(67931) <= 8029614;
srom_1(67932) <= 7456877;
srom_1(67933) <= 6888509;
srom_1(67934) <= 6327175;
srom_1(67935) <= 5775509;
srom_1(67936) <= 5236096;
srom_1(67937) <= 4711466;
srom_1(67938) <= 4204080;
srom_1(67939) <= 3716316;
srom_1(67940) <= 3250462;
srom_1(67941) <= 2808703;
srom_1(67942) <= 2393110;
srom_1(67943) <= 2005632;
srom_1(67944) <= 1648086;
srom_1(67945) <= 1322148;
srom_1(67946) <= 1029348;
srom_1(67947) <= 771057;
srom_1(67948) <= 548488;
srom_1(67949) <= 362684;
srom_1(67950) <= 214516;
srom_1(67951) <= 104679;
srom_1(67952) <= 33689;
srom_1(67953) <= 1877;
srom_1(67954) <= 9394;
srom_1(67955) <= 56204;
srom_1(67956) <= 142087;
srom_1(67957) <= 266642;
srom_1(67958) <= 429282;
srom_1(67959) <= 629247;
srom_1(67960) <= 865598;
srom_1(67961) <= 1137227;
srom_1(67962) <= 1442860;
srom_1(67963) <= 1781065;
srom_1(67964) <= 2150254;
srom_1(67965) <= 2548697;
srom_1(67966) <= 2974525;
srom_1(67967) <= 3425742;
srom_1(67968) <= 3900232;
srom_1(67969) <= 4395769;
srom_1(67970) <= 4910030;
srom_1(67971) <= 5440603;
srom_1(67972) <= 5985000;
srom_1(67973) <= 6540668;
srom_1(67974) <= 7105003;
srom_1(67975) <= 7675356;
srom_1(67976) <= 8249054;
srom_1(67977) <= 8823407;
srom_1(67978) <= 9395720;
srom_1(67979) <= 9963311;
srom_1(67980) <= 10523518;
srom_1(67981) <= 11073713;
srom_1(67982) <= 11611317;
srom_1(67983) <= 12133808;
srom_1(67984) <= 12638737;
srom_1(67985) <= 13123736;
srom_1(67986) <= 13586530;
srom_1(67987) <= 14024949;
srom_1(67988) <= 14436937;
srom_1(67989) <= 14820563;
srom_1(67990) <= 15174027;
srom_1(67991) <= 15495672;
srom_1(67992) <= 15783989;
srom_1(67993) <= 16037627;
srom_1(67994) <= 16255396;
srom_1(67995) <= 16436275;
srom_1(67996) <= 16579415;
srom_1(67997) <= 16684146;
srom_1(67998) <= 16749977;
srom_1(67999) <= 16776598;
srom_1(68000) <= 16763885;
srom_1(68001) <= 16711897;
srom_1(68002) <= 16620879;
srom_1(68003) <= 16491257;
srom_1(68004) <= 16323638;
srom_1(68005) <= 16118810;
srom_1(68006) <= 15877732;
srom_1(68007) <= 15601534;
srom_1(68008) <= 15291513;
srom_1(68009) <= 14949122;
srom_1(68010) <= 14575967;
srom_1(68011) <= 14173796;
srom_1(68012) <= 13744497;
srom_1(68013) <= 13290082;
srom_1(68014) <= 12812683;
srom_1(68015) <= 12314538;
srom_1(68016) <= 11797982;
srom_1(68017) <= 11265439;
srom_1(68018) <= 10719405;
srom_1(68019) <= 10162442;
srom_1(68020) <= 9597160;
srom_1(68021) <= 9026211;
srom_1(68022) <= 8452272;
srom_1(68023) <= 7878034;
srom_1(68024) <= 7306191;
srom_1(68025) <= 6739424;
srom_1(68026) <= 6180390;
srom_1(68027) <= 5631711;
srom_1(68028) <= 5095960;
srom_1(68029) <= 4575650;
srom_1(68030) <= 4073220;
srom_1(68031) <= 3591026;
srom_1(68032) <= 3131330;
srom_1(68033) <= 2696287;
srom_1(68034) <= 2287937;
srom_1(68035) <= 1908195;
srom_1(68036) <= 1558842;
srom_1(68037) <= 1241516;
srom_1(68038) <= 957706;
srom_1(68039) <= 708741;
srom_1(68040) <= 495790;
srom_1(68041) <= 319851;
srom_1(68042) <= 181750;
srom_1(68043) <= 82133;
srom_1(68044) <= 21468;
srom_1(68045) <= 39;
srom_1(68046) <= 17947;
srom_1(68047) <= 75108;
srom_1(68048) <= 171254;
srom_1(68049) <= 305934;
srom_1(68050) <= 478517;
srom_1(68051) <= 688192;
srom_1(68052) <= 933977;
srom_1(68053) <= 1214720;
srom_1(68054) <= 1529104;
srom_1(68055) <= 1875654;
srom_1(68056) <= 2252745;
srom_1(68057) <= 2658610;
srom_1(68058) <= 3091345;
srom_1(68059) <= 3548920;
srom_1(68060) <= 4029190;
srom_1(68061) <= 4529903;
srom_1(68062) <= 5048711;
srom_1(68063) <= 5583181;
srom_1(68064) <= 6130807;
srom_1(68065) <= 6689020;
srom_1(68066) <= 7255202;
srom_1(68067) <= 7826700;
srom_1(68068) <= 8400833;
srom_1(68069) <= 8974909;
srom_1(68070) <= 9546235;
srom_1(68071) <= 10112132;
srom_1(68072) <= 10669948;
srom_1(68073) <= 11217065;
srom_1(68074) <= 11750919;
srom_1(68075) <= 12269006;
srom_1(68076) <= 12768896;
srom_1(68077) <= 13248245;
srom_1(68078) <= 13704807;
srom_1(68079) <= 14136438;
srom_1(68080) <= 14541116;
srom_1(68081) <= 14916943;
srom_1(68082) <= 15262156;
srom_1(68083) <= 15575137;
srom_1(68084) <= 15854417;
srom_1(68085) <= 16098688;
srom_1(68086) <= 16306804;
srom_1(68087) <= 16477788;
srom_1(68088) <= 16610840;
srom_1(68089) <= 16705334;
srom_1(68090) <= 16760829;
srom_1(68091) <= 16777063;
srom_1(68092) <= 16753962;
srom_1(68093) <= 16691632;
srom_1(68094) <= 16590366;
srom_1(68095) <= 16450639;
srom_1(68096) <= 16273107;
srom_1(68097) <= 16058602;
srom_1(68098) <= 15808129;
srom_1(68099) <= 15522864;
srom_1(68100) <= 15204144;
srom_1(68101) <= 14853463;
srom_1(68102) <= 14472466;
srom_1(68103) <= 14062941;
srom_1(68104) <= 13626806;
srom_1(68105) <= 13166107;
srom_1(68106) <= 12683005;
srom_1(68107) <= 12179766;
srom_1(68108) <= 11658748;
srom_1(68109) <= 11122395;
srom_1(68110) <= 10573223;
srom_1(68111) <= 10013806;
srom_1(68112) <= 9446768;
srom_1(68113) <= 8874768;
srom_1(68114) <= 8300489;
srom_1(68115) <= 7726622;
srom_1(68116) <= 7155860;
srom_1(68117) <= 6590879;
srom_1(68118) <= 6034327;
srom_1(68119) <= 5488816;
srom_1(68120) <= 4956903;
srom_1(68121) <= 4441082;
srom_1(68122) <= 3943773;
srom_1(68123) <= 3467307;
srom_1(68124) <= 3013918;
srom_1(68125) <= 2585734;
srom_1(68126) <= 2184761;
srom_1(68127) <= 1812880;
srom_1(68128) <= 1471835;
srom_1(68129) <= 1163225;
srom_1(68130) <= 888497;
srom_1(68131) <= 648940;
srom_1(68132) <= 445676;
srom_1(68133) <= 279660;
srom_1(68134) <= 151670;
srom_1(68135) <= 62305;
srom_1(68136) <= 11986;
srom_1(68137) <= 947;
srom_1(68138) <= 29241;
srom_1(68139) <= 96734;
srom_1(68140) <= 203111;
srom_1(68141) <= 347873;
srom_1(68142) <= 530341;
srom_1(68143) <= 749658;
srom_1(68144) <= 1004797;
srom_1(68145) <= 1294562;
srom_1(68146) <= 1617593;
srom_1(68147) <= 1972375;
srom_1(68148) <= 2357246;
srom_1(68149) <= 2770399;
srom_1(68150) <= 3209898;
srom_1(68151) <= 3673682;
srom_1(68152) <= 4159576;
srom_1(68153) <= 4665301;
srom_1(68154) <= 5188487;
srom_1(68155) <= 5726678;
srom_1(68156) <= 6277352;
srom_1(68157) <= 6837927;
srom_1(68158) <= 7405773;
srom_1(68159) <= 7978229;
srom_1(68160) <= 8552608;
srom_1(68161) <= 9126219;
srom_1(68162) <= 9696370;
srom_1(68163) <= 10260389;
srom_1(68164) <= 10815631;
srom_1(68165) <= 11359491;
srom_1(68166) <= 11889420;
srom_1(68167) <= 12402933;
srom_1(68168) <= 12897621;
srom_1(68169) <= 13371164;
srom_1(68170) <= 13821343;
srom_1(68171) <= 14246046;
srom_1(68172) <= 14643281;
srom_1(68173) <= 15011185;
srom_1(68174) <= 15348035;
srom_1(68175) <= 15652249;
srom_1(68176) <= 15922401;
srom_1(68177) <= 16157225;
srom_1(68178) <= 16355619;
srom_1(68179) <= 16516653;
srom_1(68180) <= 16639572;
srom_1(68181) <= 16723799;
srom_1(68182) <= 16768940;
srom_1(68183) <= 16774783;
srom_1(68184) <= 16741299;
srom_1(68185) <= 16668647;
srom_1(68186) <= 16557168;
srom_1(68187) <= 16407382;
srom_1(68188) <= 16219995;
srom_1(68189) <= 15995883;
srom_1(68190) <= 15736098;
srom_1(68191) <= 15441858;
srom_1(68192) <= 15114543;
srom_1(68193) <= 14755687;
srom_1(68194) <= 14366975;
srom_1(68195) <= 13950227;
srom_1(68196) <= 13507400;
srom_1(68197) <= 13040568;
srom_1(68198) <= 12551922;
srom_1(68199) <= 12043753;
srom_1(68200) <= 11518443;
srom_1(68201) <= 10978457;
srom_1(68202) <= 10426325;
srom_1(68203) <= 9864639;
srom_1(68204) <= 9296030;
srom_1(68205) <= 8723167;
srom_1(68206) <= 8148734;
srom_1(68207) <= 7575427;
srom_1(68208) <= 7005933;
srom_1(68209) <= 6442922;
srom_1(68210) <= 5889036;
srom_1(68211) <= 5346870;
srom_1(68212) <= 4818969;
srom_1(68213) <= 4307807;
srom_1(68214) <= 3815781;
srom_1(68215) <= 3345199;
srom_1(68216) <= 2898267;
srom_1(68217) <= 2477081;
srom_1(68218) <= 2083616;
srom_1(68219) <= 1719717;
srom_1(68220) <= 1387092;
srom_1(68221) <= 1087298;
srom_1(68222) <= 821743;
srom_1(68223) <= 591672;
srom_1(68224) <= 398163;
srom_1(68225) <= 242124;
srom_1(68226) <= 124287;
srom_1(68227) <= 45204;
srom_1(68228) <= 5246;
srom_1(68229) <= 4601;
srom_1(68230) <= 43271;
srom_1(68231) <= 121075;
srom_1(68232) <= 237648;
srom_1(68233) <= 392444;
srom_1(68234) <= 584737;
srom_1(68235) <= 813625;
srom_1(68236) <= 1078035;
srom_1(68237) <= 1376726;
srom_1(68238) <= 1708299;
srom_1(68239) <= 2071197;
srom_1(68240) <= 2463720;
srom_1(68241) <= 2884028;
srom_1(68242) <= 3330147;
srom_1(68243) <= 3799988;
srom_1(68244) <= 4291347;
srom_1(68245) <= 4801918;
srom_1(68246) <= 5329309;
srom_1(68247) <= 5871047;
srom_1(68248) <= 6424589;
srom_1(68249) <= 6987342;
srom_1(68250) <= 7556666;
srom_1(68251) <= 8129891;
srom_1(68252) <= 8704329;
srom_1(68253) <= 9277287;
srom_1(68254) <= 9846078;
srom_1(68255) <= 10408033;
srom_1(68256) <= 10960519;
srom_1(68257) <= 11500945;
srom_1(68258) <= 12026776;
srom_1(68259) <= 12535546;
srom_1(68260) <= 13024869;
srom_1(68261) <= 13492452;
srom_1(68262) <= 13936101;
srom_1(68263) <= 14353735;
srom_1(68264) <= 14743398;
srom_1(68265) <= 15103260;
srom_1(68266) <= 15431635;
srom_1(68267) <= 15726983;
srom_1(68268) <= 15987919;
srom_1(68269) <= 16213219;
srom_1(68270) <= 16401826;
srom_1(68271) <= 16552857;
srom_1(68272) <= 16665603;
srom_1(68273) <= 16739536;
srom_1(68274) <= 16774308;
srom_1(68275) <= 16769756;
srom_1(68276) <= 16725902;
srom_1(68277) <= 16642952;
srom_1(68278) <= 16521295;
srom_1(68279) <= 16361500;
srom_1(68280) <= 16164318;
srom_1(68281) <= 15930673;
srom_1(68282) <= 15661661;
srom_1(68283) <= 15358542;
srom_1(68284) <= 15022740;
srom_1(68285) <= 14655827;
srom_1(68286) <= 14259526;
srom_1(68287) <= 13835693;
srom_1(68288) <= 13386318;
srom_1(68289) <= 12913506;
srom_1(68290) <= 12419475;
srom_1(68291) <= 11906543;
srom_1(68292) <= 11377114;
srom_1(68293) <= 10833670;
srom_1(68294) <= 10278761;
srom_1(68295) <= 9714988;
srom_1(68296) <= 9144995;
srom_1(68297) <= 8571456;
srom_1(68298) <= 7997059;
srom_1(68299) <= 7424498;
srom_1(68300) <= 6856458;
srom_1(68301) <= 6295602;
srom_1(68302) <= 5744562;
srom_1(68303) <= 5205921;
srom_1(68304) <= 4682204;
srom_1(68305) <= 4175868;
srom_1(68306) <= 3689286;
srom_1(68307) <= 3224742;
srom_1(68308) <= 2784412;
srom_1(68309) <= 2370363;
srom_1(68310) <= 1984535;
srom_1(68311) <= 1628738;
srom_1(68312) <= 1304641;
srom_1(68313) <= 1013762;
srom_1(68314) <= 757467;
srom_1(68315) <= 536957;
srom_1(68316) <= 353266;
srom_1(68317) <= 207255;
srom_1(68318) <= 99610;
srom_1(68319) <= 30834;
srom_1(68320) <= 1251;
srom_1(68321) <= 10999;
srom_1(68322) <= 60033;
srom_1(68323) <= 148122;
srom_1(68324) <= 274854;
srom_1(68325) <= 439634;
srom_1(68326) <= 641689;
srom_1(68327) <= 880072;
srom_1(68328) <= 1153665;
srom_1(68329) <= 1461186;
srom_1(68330) <= 1801191;
srom_1(68331) <= 2172088;
srom_1(68332) <= 2572135;
srom_1(68333) <= 2999458;
srom_1(68334) <= 3452053;
srom_1(68335) <= 3927796;
srom_1(68336) <= 4424458;
srom_1(68337) <= 4939710;
srom_1(68338) <= 5471134;
srom_1(68339) <= 6016239;
srom_1(68340) <= 6572470;
srom_1(68341) <= 7137216;
srom_1(68342) <= 7707831;
srom_1(68343) <= 8281638;
srom_1(68344) <= 8855947;
srom_1(68345) <= 9428065;
srom_1(68346) <= 9995308;
srom_1(68347) <= 10555016;
srom_1(68348) <= 11104566;
srom_1(68349) <= 11641379;
srom_1(68350) <= 12162940;
srom_1(68351) <= 12666801;
srom_1(68352) <= 13150600;
srom_1(68353) <= 13612068;
srom_1(68354) <= 14049042;
srom_1(68355) <= 14459472;
srom_1(68356) <= 14841434;
srom_1(68357) <= 15193136;
srom_1(68358) <= 15512930;
srom_1(68359) <= 15799315;
srom_1(68360) <= 16050948;
srom_1(68361) <= 16266651;
srom_1(68362) <= 16445410;
srom_1(68363) <= 16586389;
srom_1(68364) <= 16688925;
srom_1(68365) <= 16752538;
srom_1(68366) <= 16776930;
srom_1(68367) <= 16761986;
srom_1(68368) <= 16707776;
srom_1(68369) <= 16614555;
srom_1(68370) <= 16482760;
srom_1(68371) <= 16313008;
srom_1(68372) <= 16106096;
srom_1(68373) <= 15862994;
srom_1(68374) <= 15584842;
srom_1(68375) <= 15272945;
srom_1(68376) <= 14928765;
srom_1(68377) <= 14553915;
srom_1(68378) <= 14150154;
srom_1(68379) <= 13719376;
srom_1(68380) <= 13263599;
srom_1(68381) <= 12784962;
srom_1(68382) <= 12285709;
srom_1(68383) <= 11768181;
srom_1(68384) <= 11234806;
srom_1(68385) <= 10688083;
srom_1(68386) <= 10130577;
srom_1(68387) <= 9564903;
srom_1(68388) <= 8993713;
srom_1(68389) <= 8419685;
srom_1(68390) <= 7845511;
srom_1(68391) <= 7273884;
srom_1(68392) <= 6707484;
srom_1(68393) <= 6148968;
srom_1(68394) <= 5600954;
srom_1(68395) <= 5066013;
srom_1(68396) <= 4546652;
srom_1(68397) <= 4045307;
srom_1(68398) <= 3564330;
srom_1(68399) <= 3105975;
srom_1(68400) <= 2672393;
srom_1(68401) <= 2265616;
srom_1(68402) <= 1887551;
srom_1(68403) <= 1539972;
srom_1(68404) <= 1224509;
srom_1(68405) <= 942641;
srom_1(68406) <= 695689;
srom_1(68407) <= 484813;
srom_1(68408) <= 310999;
srom_1(68409) <= 175065;
srom_1(68410) <= 77646;
srom_1(68411) <= 19201;
srom_1(68412) <= 2;
srom_1(68413) <= 20141;
srom_1(68414) <= 79522;
srom_1(68415) <= 177867;
srom_1(68416) <= 314716;
srom_1(68417) <= 489425;
srom_1(68418) <= 701177;
srom_1(68419) <= 948977;
srom_1(68420) <= 1231665;
srom_1(68421) <= 1547914;
srom_1(68422) <= 1896241;
srom_1(68423) <= 2275013;
srom_1(68424) <= 2682454;
srom_1(68425) <= 3116653;
srom_1(68426) <= 3575574;
srom_1(68427) <= 4057065;
srom_1(68428) <= 4558868;
srom_1(68429) <= 5078630;
srom_1(68430) <= 5613914;
srom_1(68431) <= 6162209;
srom_1(68432) <= 6720944;
srom_1(68433) <= 7287500;
srom_1(68434) <= 7859219;
srom_1(68435) <= 8433421;
srom_1(68436) <= 9007412;
srom_1(68437) <= 9578502;
srom_1(68438) <= 10144012;
srom_1(68439) <= 10701290;
srom_1(68440) <= 11247723;
srom_1(68441) <= 11780749;
srom_1(68442) <= 12297868;
srom_1(68443) <= 12796655;
srom_1(68444) <= 13274771;
srom_1(68445) <= 13729975;
srom_1(68446) <= 14160130;
srom_1(68447) <= 14563221;
srom_1(68448) <= 14937358;
srom_1(68449) <= 15280785;
srom_1(68450) <= 15591892;
srom_1(68451) <= 15869220;
srom_1(68452) <= 16111469;
srom_1(68453) <= 16317503;
srom_1(68454) <= 16486356;
srom_1(68455) <= 16617236;
srom_1(68456) <= 16709529;
srom_1(68457) <= 16762802;
srom_1(68458) <= 16776805;
srom_1(68459) <= 16751474;
srom_1(68460) <= 16686926;
srom_1(68461) <= 16583464;
srom_1(68462) <= 16441574;
srom_1(68463) <= 16261921;
srom_1(68464) <= 16045347;
srom_1(68465) <= 15792868;
srom_1(68466) <= 15505668;
srom_1(68467) <= 15185094;
srom_1(68468) <= 14832648;
srom_1(68469) <= 14449984;
srom_1(68470) <= 14038897;
srom_1(68471) <= 13601313;
srom_1(68472) <= 13139285;
srom_1(68473) <= 12654979;
srom_1(68474) <= 12150667;
srom_1(68475) <= 11628714;
srom_1(68476) <= 11091566;
srom_1(68477) <= 10541743;
srom_1(68478) <= 9981824;
srom_1(68479) <= 9414433;
srom_1(68480) <= 8842232;
srom_1(68481) <= 8267903;
srom_1(68482) <= 7694141;
srom_1(68483) <= 7123635;
srom_1(68484) <= 6559062;
srom_1(68485) <= 6003067;
srom_1(68486) <= 5458259;
srom_1(68487) <= 4927193;
srom_1(68488) <= 4412358;
srom_1(68489) <= 3916169;
srom_1(68490) <= 3440953;
srom_1(68491) <= 2988939;
srom_1(68492) <= 2562245;
srom_1(68493) <= 2162873;
srom_1(68494) <= 1792696;
srom_1(68495) <= 1453449;
srom_1(68496) <= 1146723;
srom_1(68497) <= 873957;
srom_1(68498) <= 636430;
srom_1(68499) <= 435256;
srom_1(68500) <= 271377;
srom_1(68501) <= 145563;
srom_1(68502) <= 58404;
srom_1(68503) <= 10307;
srom_1(68504) <= 1500;
srom_1(68505) <= 32022;
srom_1(68506) <= 101731;
srom_1(68507) <= 210301;
srom_1(68508) <= 357221;
srom_1(68509) <= 541803;
srom_1(68510) <= 763181;
srom_1(68511) <= 1020318;
srom_1(68512) <= 1312007;
srom_1(68513) <= 1636881;
srom_1(68514) <= 1993416;
srom_1(68515) <= 2379940;
srom_1(68516) <= 2794641;
srom_1(68517) <= 3235574;
srom_1(68518) <= 3700671;
srom_1(68519) <= 4187752;
srom_1(68520) <= 4694531;
srom_1(68521) <= 5218634;
srom_1(68522) <= 5757602;
srom_1(68523) <= 6308907;
srom_1(68524) <= 6869965;
srom_1(68525) <= 7438144;
srom_1(68526) <= 8010780;
srom_1(68527) <= 8585188;
srom_1(68528) <= 9158675;
srom_1(68529) <= 9728550;
srom_1(68530) <= 10292141;
srom_1(68531) <= 10846807;
srom_1(68532) <= 11389945;
srom_1(68533) <= 11919008;
srom_1(68534) <= 12431517;
srom_1(68535) <= 12925066;
srom_1(68536) <= 13397343;
srom_1(68537) <= 13846132;
srom_1(68538) <= 14269329;
srom_1(68539) <= 14664949;
srom_1(68540) <= 15031137;
srom_1(68541) <= 15366176;
srom_1(68542) <= 15668495;
srom_1(68543) <= 15936676;
srom_1(68544) <= 16169462;
srom_1(68545) <= 16365760;
srom_1(68546) <= 16524651;
srom_1(68547) <= 16645389;
srom_1(68548) <= 16727408;
srom_1(68549) <= 16770324;
srom_1(68550) <= 16773935;
srom_1(68551) <= 16738224;
srom_1(68552) <= 16663359;
srom_1(68553) <= 16549691;
srom_1(68554) <= 16397753;
srom_1(68555) <= 16208257;
srom_1(68556) <= 15982092;
srom_1(68557) <= 15720318;
srom_1(68558) <= 15424164;
srom_1(68559) <= 15095017;
srom_1(68560) <= 14734422;
srom_1(68561) <= 14344069;
srom_1(68562) <= 13925789;
srom_1(68563) <= 13481544;
srom_1(68564) <= 13013415;
srom_1(68565) <= 12523600;
srom_1(68566) <= 12014394;
srom_1(68567) <= 11488185;
srom_1(68568) <= 10947441;
srom_1(68569) <= 10394698;
srom_1(68570) <= 9832548;
srom_1(68571) <= 9263627;
srom_1(68572) <= 8690603;
srom_1(68573) <= 8116162;
srom_1(68574) <= 7542999;
srom_1(68575) <= 6973801;
srom_1(68576) <= 6411238;
srom_1(68577) <= 5857947;
srom_1(68578) <= 5316523;
srom_1(68579) <= 4789506;
srom_1(68580) <= 4279366;
srom_1(68581) <= 3788495;
srom_1(68582) <= 3319196;
srom_1(68583) <= 2873670;
srom_1(68584) <= 2454004;
srom_1(68585) <= 2062168;
srom_1(68586) <= 1699999;
srom_1(68587) <= 1369195;
srom_1(68588) <= 1071308;
srom_1(68589) <= 807734;
srom_1(68590) <= 579709;
srom_1(68591) <= 388303;
srom_1(68592) <= 234413;
srom_1(68593) <= 118761;
srom_1(68594) <= 41888;
srom_1(68595) <= 4157;
srom_1(68596) <= 5743;
srom_1(68597) <= 46639;
srom_1(68598) <= 126654;
srom_1(68599) <= 245412;
srom_1(68600) <= 402356;
srom_1(68601) <= 596750;
srom_1(68602) <= 827683;
srom_1(68603) <= 1094071;
srom_1(68604) <= 1394667;
srom_1(68605) <= 1728059;
srom_1(68606) <= 2092685;
srom_1(68607) <= 2486834;
srom_1(68608) <= 2908659;
srom_1(68609) <= 3356182;
srom_1(68610) <= 3827303;
srom_1(68611) <= 4319814;
srom_1(68612) <= 4831404;
srom_1(68613) <= 5359676;
srom_1(68614) <= 5902151;
srom_1(68615) <= 6456286;
srom_1(68616) <= 7019483;
srom_1(68617) <= 7589099;
srom_1(68618) <= 8162465;
srom_1(68619) <= 8736892;
srom_1(68620) <= 9309685;
srom_1(68621) <= 9878159;
srom_1(68622) <= 10439648;
srom_1(68623) <= 10991518;
srom_1(68624) <= 11531183;
srom_1(68625) <= 12056111;
srom_1(68626) <= 12563841;
srom_1(68627) <= 13051992;
srom_1(68628) <= 13518275;
srom_1(68629) <= 13960503;
srom_1(68630) <= 14376602;
srom_1(68631) <= 14764622;
srom_1(68632) <= 15122742;
srom_1(68633) <= 15449284;
srom_1(68634) <= 15742716;
srom_1(68635) <= 16001661;
srom_1(68636) <= 16224907;
srom_1(68637) <= 16411405;
srom_1(68638) <= 16560282;
srom_1(68639) <= 16670839;
srom_1(68640) <= 16742558;
srom_1(68641) <= 16775102;
srom_1(68642) <= 16768319;
srom_1(68643) <= 16722241;
srom_1(68644) <= 16637083;
srom_1(68645) <= 16513245;
srom_1(68646) <= 16351309;
srom_1(68647) <= 16152032;
srom_1(68648) <= 15916350;
srom_1(68649) <= 15645368;
srom_1(68650) <= 15340356;
srom_1(68651) <= 15002745;
srom_1(68652) <= 14634119;
srom_1(68653) <= 14236205;
srom_1(68654) <= 13810869;
srom_1(68655) <= 13360107;
srom_1(68656) <= 12886031;
srom_1(68657) <= 12390866;
srom_1(68658) <= 11876933;
srom_1(68659) <= 11346641;
srom_1(68660) <= 10802479;
srom_1(68661) <= 10246997;
srom_1(68662) <= 9682800;
srom_1(68663) <= 9112535;
srom_1(68664) <= 8538874;
srom_1(68665) <= 7964509;
srom_1(68666) <= 7392133;
srom_1(68667) <= 6824430;
srom_1(68668) <= 6264061;
srom_1(68669) <= 5713655;
srom_1(68670) <= 5175793;
srom_1(68671) <= 4652997;
srom_1(68672) <= 4147719;
srom_1(68673) <= 3662328;
srom_1(68674) <= 3199099;
srom_1(68675) <= 2760206;
srom_1(68676) <= 2347707;
srom_1(68677) <= 1963535;
srom_1(68678) <= 1609493;
srom_1(68679) <= 1287240;
srom_1(68680) <= 998289;
srom_1(68681) <= 743992;
srom_1(68682) <= 525544;
srom_1(68683) <= 343969;
srom_1(68684) <= 200118;
srom_1(68685) <= 94665;
srom_1(68686) <= 28106;
srom_1(68687) <= 752;
srom_1(68688) <= 12731;
srom_1(68689) <= 63988;
srom_1(68690) <= 154281;
srom_1(68691) <= 283189;
srom_1(68692) <= 450105;
srom_1(68693) <= 654248;
srom_1(68694) <= 894659;
srom_1(68695) <= 1170213;
srom_1(68696) <= 1479616;
srom_1(68697) <= 1821417;
srom_1(68698) <= 2194015;
srom_1(68699) <= 2595661;
srom_1(68700) <= 3024472;
srom_1(68701) <= 3478437;
srom_1(68702) <= 3955428;
srom_1(68703) <= 4453208;
srom_1(68704) <= 4969442;
srom_1(68705) <= 5501709;
srom_1(68706) <= 6047515;
srom_1(68707) <= 6604298;
srom_1(68708) <= 7169449;
srom_1(68709) <= 7740317;
srom_1(68710) <= 8314224;
srom_1(68711) <= 8888481;
srom_1(68712) <= 9460393;
srom_1(68713) <= 10027280;
srom_1(68714) <= 10586482;
srom_1(68715) <= 11135378;
srom_1(68716) <= 11671393;
srom_1(68717) <= 12192014;
srom_1(68718) <= 12694799;
srom_1(68719) <= 13177392;
srom_1(68720) <= 13637528;
srom_1(68721) <= 14073050;
srom_1(68722) <= 14481915;
srom_1(68723) <= 14862208;
srom_1(68724) <= 15212143;
srom_1(68725) <= 15530080;
srom_1(68726) <= 15814528;
srom_1(68727) <= 16064154;
srom_1(68728) <= 16277787;
srom_1(68729) <= 16454424;
srom_1(68730) <= 16593238;
srom_1(68731) <= 16693578;
srom_1(68732) <= 16754972;
srom_1(68733) <= 16777134;
srom_1(68734) <= 16759960;
srom_1(68735) <= 16703529;
srom_1(68736) <= 16608107;
srom_1(68737) <= 16474140;
srom_1(68738) <= 16302258;
srom_1(68739) <= 16093266;
srom_1(68740) <= 15848144;
srom_1(68741) <= 15568042;
srom_1(68742) <= 15254273;
srom_1(68743) <= 14908308;
srom_1(68744) <= 14531770;
srom_1(68745) <= 14126425;
srom_1(68746) <= 13694174;
srom_1(68747) <= 13237043;
srom_1(68748) <= 12757175;
srom_1(68749) <= 12256822;
srom_1(68750) <= 11738330;
srom_1(68751) <= 11204130;
srom_1(68752) <= 10656726;
srom_1(68753) <= 10098687;
srom_1(68754) <= 9532628;
srom_1(68755) <= 8961205;
srom_1(68756) <= 8387097;
srom_1(68757) <= 7812996;
srom_1(68758) <= 7241594;
srom_1(68759) <= 6675570;
srom_1(68760) <= 6117580;
srom_1(68761) <= 5570240;
srom_1(68762) <= 5036115;
srom_1(68763) <= 4517712;
srom_1(68764) <= 4017461;
srom_1(68765) <= 3537707;
srom_1(68766) <= 3080701;
srom_1(68767) <= 2648585;
srom_1(68768) <= 2243387;
srom_1(68769) <= 1867006;
srom_1(68770) <= 1521206;
srom_1(68771) <= 1207610;
srom_1(68772) <= 927689;
srom_1(68773) <= 682754;
srom_1(68774) <= 473954;
srom_1(68775) <= 302269;
srom_1(68776) <= 168504;
srom_1(68777) <= 73285;
srom_1(68778) <= 17060;
srom_1(68779) <= 92;
srom_1(68780) <= 22461;
srom_1(68781) <= 84061;
srom_1(68782) <= 184604;
srom_1(68783) <= 323619;
srom_1(68784) <= 500453;
srom_1(68785) <= 714277;
srom_1(68786) <= 964089;
srom_1(68787) <= 1248717;
srom_1(68788) <= 1566827;
srom_1(68789) <= 1916926;
srom_1(68790) <= 2297373;
srom_1(68791) <= 2706384;
srom_1(68792) <= 3142041;
srom_1(68793) <= 3602300;
srom_1(68794) <= 4085005;
srom_1(68795) <= 4587890;
srom_1(68796) <= 5108599;
srom_1(68797) <= 5644688;
srom_1(68798) <= 6193645;
srom_1(68799) <= 6752894;
srom_1(68800) <= 7319814;
srom_1(68801) <= 7891746;
srom_1(68802) <= 8466008;
srom_1(68803) <= 9039907;
srom_1(68804) <= 9610751;
srom_1(68805) <= 10175865;
srom_1(68806) <= 10732597;
srom_1(68807) <= 11278338;
srom_1(68808) <= 11810528;
srom_1(68809) <= 12326671;
srom_1(68810) <= 12824348;
srom_1(68811) <= 13301223;
srom_1(68812) <= 13755062;
srom_1(68813) <= 14183735;
srom_1(68814) <= 14585234;
srom_1(68815) <= 14957674;
srom_1(68816) <= 15299309;
srom_1(68817) <= 15608538;
srom_1(68818) <= 15883910;
srom_1(68819) <= 16124134;
srom_1(68820) <= 16328083;
srom_1(68821) <= 16494802;
srom_1(68822) <= 16623508;
srom_1(68823) <= 16713597;
srom_1(68824) <= 16764648;
srom_1(68825) <= 16776420;
srom_1(68826) <= 16748860;
srom_1(68827) <= 16682095;
srom_1(68828) <= 16576439;
srom_1(68829) <= 16432388;
srom_1(68830) <= 16250616;
srom_1(68831) <= 16031977;
srom_1(68832) <= 15777496;
srom_1(68833) <= 15488365;
srom_1(68834) <= 15165941;
srom_1(68835) <= 14811736;
srom_1(68836) <= 14427411;
srom_1(68837) <= 14014768;
srom_1(68838) <= 13575741;
srom_1(68839) <= 13112391;
srom_1(68840) <= 12626889;
srom_1(68841) <= 12121512;
srom_1(68842) <= 11598630;
srom_1(68843) <= 11060696;
srom_1(68844) <= 10510231;
srom_1(68845) <= 9949817;
srom_1(68846) <= 9382082;
srom_1(68847) <= 8809688;
srom_1(68848) <= 8235320;
srom_1(68849) <= 7661671;
srom_1(68850) <= 7091430;
srom_1(68851) <= 6527272;
srom_1(68852) <= 5971843;
srom_1(68853) <= 5427747;
srom_1(68854) <= 4897535;
srom_1(68855) <= 4383694;
srom_1(68856) <= 3888633;
srom_1(68857) <= 3414675;
srom_1(68858) <= 2964040;
srom_1(68859) <= 2538844;
srom_1(68860) <= 2141079;
srom_1(68861) <= 1772611;
srom_1(68862) <= 1435167;
srom_1(68863) <= 1130331;
srom_1(68864) <= 859531;
srom_1(68865) <= 624038;
srom_1(68866) <= 424955;
srom_1(68867) <= 263217;
srom_1(68868) <= 139581;
srom_1(68869) <= 54628;
srom_1(68870) <= 8756;
srom_1(68871) <= 2179;
srom_1(68872) <= 34930;
srom_1(68873) <= 106854;
srom_1(68874) <= 217614;
srom_1(68875) <= 366690;
srom_1(68876) <= 553384;
srom_1(68877) <= 776820;
srom_1(68878) <= 1035950;
srom_1(68879) <= 1329560;
srom_1(68880) <= 1656271;
srom_1(68881) <= 2014553;
srom_1(68882) <= 2402725;
srom_1(68883) <= 2818967;
srom_1(68884) <= 3261327;
srom_1(68885) <= 3727731;
srom_1(68886) <= 4215990;
srom_1(68887) <= 4723817;
srom_1(68888) <= 5248829;
srom_1(68889) <= 5788565;
srom_1(68890) <= 6340493;
srom_1(68891) <= 6902026;
srom_1(68892) <= 7470529;
srom_1(68893) <= 8043338;
srom_1(68894) <= 8617766;
srom_1(68895) <= 9191119;
srom_1(68896) <= 9760709;
srom_1(68897) <= 10323865;
srom_1(68898) <= 10877945;
srom_1(68899) <= 11420352;
srom_1(68900) <= 11948543;
srom_1(68901) <= 12460039;
srom_1(68902) <= 12952444;
srom_1(68903) <= 13423446;
srom_1(68904) <= 13870839;
srom_1(68905) <= 14292524;
srom_1(68906) <= 14686523;
srom_1(68907) <= 15050989;
srom_1(68908) <= 15384213;
srom_1(68909) <= 15684632;
srom_1(68910) <= 15950837;
srom_1(68911) <= 16181581;
srom_1(68912) <= 16375781;
srom_1(68913) <= 16532526;
srom_1(68914) <= 16651081;
srom_1(68915) <= 16730891;
srom_1(68916) <= 16771581;
srom_1(68917) <= 16772960;
srom_1(68918) <= 16735023;
srom_1(68919) <= 16657946;
srom_1(68920) <= 16542091;
srom_1(68921) <= 16388002;
srom_1(68922) <= 16196401;
srom_1(68923) <= 15968186;
srom_1(68924) <= 15704428;
srom_1(68925) <= 15406364;
srom_1(68926) <= 15075391;
srom_1(68927) <= 14713062;
srom_1(68928) <= 14321074;
srom_1(68929) <= 13901268;
srom_1(68930) <= 13455611;
srom_1(68931) <= 12986193;
srom_1(68932) <= 12495215;
srom_1(68933) <= 11984980;
srom_1(68934) <= 11457880;
srom_1(68935) <= 10916387;
srom_1(68936) <= 10363041;
srom_1(68937) <= 9800436;
srom_1(68938) <= 9231210;
srom_1(68939) <= 8658034;
srom_1(68940) <= 8083593;
srom_1(68941) <= 7510583;
srom_1(68942) <= 6941691;
srom_1(68943) <= 6379583;
srom_1(68944) <= 5826897;
srom_1(68945) <= 5286223;
srom_1(68946) <= 4760097;
srom_1(68947) <= 4250987;
srom_1(68948) <= 3761279;
srom_1(68949) <= 3293271;
srom_1(68950) <= 2849156;
srom_1(68951) <= 2431018;
srom_1(68952) <= 2040817;
srom_1(68953) <= 1680382;
srom_1(68954) <= 1351405;
srom_1(68955) <= 1055428;
srom_1(68956) <= 793839;
srom_1(68957) <= 567864;
srom_1(68958) <= 378563;
srom_1(68959) <= 226824;
srom_1(68960) <= 113359;
srom_1(68961) <= 38699;
srom_1(68962) <= 3194;
srom_1(68963) <= 7012;
srom_1(68964) <= 50134;
srom_1(68965) <= 132358;
srom_1(68966) <= 253298;
srom_1(68967) <= 412387;
srom_1(68968) <= 608880;
srom_1(68969) <= 841854;
srom_1(68970) <= 1110218;
srom_1(68971) <= 1412713;
srom_1(68972) <= 1747920;
srom_1(68973) <= 2114267;
srom_1(68974) <= 2510037;
srom_1(68975) <= 2933374;
srom_1(68976) <= 3382292;
srom_1(68977) <= 3854687;
srom_1(68978) <= 4348342;
srom_1(68979) <= 4860944;
srom_1(68980) <= 5390088;
srom_1(68981) <= 5933293;
srom_1(68982) <= 6488012;
srom_1(68983) <= 7051644;
srom_1(68984) <= 7621545;
srom_1(68985) <= 8195043;
srom_1(68986) <= 8769449;
srom_1(68987) <= 9342069;
srom_1(68988) <= 9910217;
srom_1(68989) <= 10471231;
srom_1(68990) <= 11022478;
srom_1(68991) <= 11561374;
srom_1(68992) <= 12085392;
srom_1(68993) <= 12592074;
srom_1(68994) <= 13079045;
srom_1(68995) <= 13544021;
srom_1(68996) <= 13984822;
srom_1(68997) <= 14399379;
srom_1(68998) <= 14785750;
srom_1(68999) <= 15142123;
srom_1(69000) <= 15466826;
srom_1(69001) <= 15758337;
srom_1(69002) <= 16015289;
srom_1(69003) <= 16236477;
srom_1(69004) <= 16420863;
srom_1(69005) <= 16567584;
srom_1(69006) <= 16675950;
srom_1(69007) <= 16745454;
srom_1(69008) <= 16775770;
srom_1(69009) <= 16766755;
srom_1(69010) <= 16718453;
srom_1(69011) <= 16631089;
srom_1(69012) <= 16505073;
srom_1(69013) <= 16340997;
srom_1(69014) <= 16139629;
srom_1(69015) <= 15901913;
srom_1(69016) <= 15628966;
srom_1(69017) <= 15322065;
srom_1(69018) <= 14982652;
srom_1(69019) <= 14612316;
srom_1(69020) <= 14212796;
srom_1(69021) <= 13785963;
srom_1(69022) <= 13333821;
srom_1(69023) <= 12858489;
srom_1(69024) <= 12362196;
srom_1(69025) <= 11847270;
srom_1(69026) <= 11316125;
srom_1(69027) <= 10771251;
srom_1(69028) <= 10215205;
srom_1(69029) <= 9650593;
srom_1(69030) <= 9080063;
srom_1(69031) <= 8506291;
srom_1(69032) <= 7931966;
srom_1(69033) <= 7359784;
srom_1(69034) <= 6792425;
srom_1(69035) <= 6232552;
srom_1(69036) <= 5682789;
srom_1(69037) <= 5145715;
srom_1(69038) <= 4623847;
srom_1(69039) <= 4119634;
srom_1(69040) <= 3635440;
srom_1(69041) <= 3173535;
srom_1(69042) <= 2736085;
srom_1(69043) <= 2325142;
srom_1(69044) <= 1942632;
srom_1(69045) <= 1590350;
srom_1(69046) <= 1269947;
srom_1(69047) <= 982926;
srom_1(69048) <= 730633;
srom_1(69049) <= 514251;
srom_1(69050) <= 334794;
srom_1(69051) <= 193104;
srom_1(69052) <= 89846;
srom_1(69053) <= 25503;
srom_1(69054) <= 379;
srom_1(69055) <= 14589;
srom_1(69056) <= 68068;
srom_1(69057) <= 160565;
srom_1(69058) <= 291646;
srom_1(69059) <= 460696;
srom_1(69060) <= 666923;
srom_1(69061) <= 909360;
srom_1(69062) <= 1186869;
srom_1(69063) <= 1498150;
srom_1(69064) <= 1841743;
srom_1(69065) <= 2216036;
srom_1(69066) <= 2619274;
srom_1(69067) <= 3049567;
srom_1(69068) <= 3504896;
srom_1(69069) <= 3983127;
srom_1(69070) <= 4482017;
srom_1(69071) <= 4999225;
srom_1(69072) <= 5532328;
srom_1(69073) <= 6078825;
srom_1(69074) <= 6636154;
srom_1(69075) <= 7201700;
srom_1(69076) <= 7772812;
srom_1(69077) <= 8346811;
srom_1(69078) <= 8921007;
srom_1(69079) <= 9492706;
srom_1(69080) <= 10059228;
srom_1(69081) <= 10617915;
srom_1(69082) <= 11166148;
srom_1(69083) <= 11701357;
srom_1(69084) <= 12221031;
srom_1(69085) <= 12722733;
srom_1(69086) <= 13204112;
srom_1(69087) <= 13662908;
srom_1(69088) <= 14096972;
srom_1(69089) <= 14504267;
srom_1(69090) <= 14882884;
srom_1(69091) <= 15231046;
srom_1(69092) <= 15547123;
srom_1(69093) <= 15829630;
srom_1(69094) <= 16077244;
srom_1(69095) <= 16288803;
srom_1(69096) <= 16463316;
srom_1(69097) <= 16599964;
srom_1(69098) <= 16698105;
srom_1(69099) <= 16757281;
srom_1(69100) <= 16777213;
srom_1(69101) <= 16757808;
srom_1(69102) <= 16699156;
srom_1(69103) <= 16601534;
srom_1(69104) <= 16465399;
srom_1(69105) <= 16291388;
srom_1(69106) <= 16080319;
srom_1(69107) <= 15833181;
srom_1(69108) <= 15551133;
srom_1(69109) <= 15235497;
srom_1(69110) <= 14887753;
srom_1(69111) <= 14509533;
srom_1(69112) <= 14102610;
srom_1(69113) <= 13668892;
srom_1(69114) <= 13210413;
srom_1(69115) <= 12729322;
srom_1(69116) <= 12227877;
srom_1(69117) <= 11708428;
srom_1(69118) <= 11173411;
srom_1(69119) <= 10625335;
srom_1(69120) <= 10066771;
srom_1(69121) <= 9500336;
srom_1(69122) <= 8928689;
srom_1(69123) <= 8354509;
srom_1(69124) <= 7780489;
srom_1(69125) <= 7209321;
srom_1(69126) <= 6643682;
srom_1(69127) <= 6086227;
srom_1(69128) <= 5539567;
srom_1(69129) <= 5006268;
srom_1(69130) <= 4488830;
srom_1(69131) <= 3989680;
srom_1(69132) <= 3511157;
srom_1(69133) <= 3055507;
srom_1(69134) <= 2624865;
srom_1(69135) <= 2221251;
srom_1(69136) <= 1846558;
srom_1(69137) <= 1502543;
srom_1(69138) <= 1190820;
srom_1(69139) <= 912849;
srom_1(69140) <= 669934;
srom_1(69141) <= 463215;
srom_1(69142) <= 293661;
srom_1(69143) <= 162067;
srom_1(69144) <= 69050;
srom_1(69145) <= 15046;
srom_1(69146) <= 309;
srom_1(69147) <= 24907;
srom_1(69148) <= 88726;
srom_1(69149) <= 191465;
srom_1(69150) <= 332644;
srom_1(69151) <= 511600;
srom_1(69152) <= 727494;
srom_1(69153) <= 979314;
srom_1(69154) <= 1265878;
srom_1(69155) <= 1585843;
srom_1(69156) <= 1937709;
srom_1(69157) <= 2319825;
srom_1(69158) <= 2730400;
srom_1(69159) <= 3167508;
srom_1(69160) <= 3629099;
srom_1(69161) <= 4113010;
srom_1(69162) <= 4616970;
srom_1(69163) <= 5138617;
srom_1(69164) <= 5675504;
srom_1(69165) <= 6225114;
srom_1(69166) <= 6784869;
srom_1(69167) <= 7352144;
srom_1(69168) <= 7924280;
srom_1(69169) <= 8498593;
srom_1(69170) <= 9072391;
srom_1(69171) <= 9642982;
srom_1(69172) <= 10207691;
srom_1(69173) <= 10763869;
srom_1(69174) <= 11308910;
srom_1(69175) <= 11840255;
srom_1(69176) <= 12355415;
srom_1(69177) <= 12851973;
srom_1(69178) <= 13327601;
srom_1(69179) <= 13780068;
srom_1(69180) <= 14207253;
srom_1(69181) <= 14607152;
srom_1(69182) <= 14977890;
srom_1(69183) <= 15317729;
srom_1(69184) <= 15625075;
srom_1(69185) <= 15898487;
srom_1(69186) <= 16136682;
srom_1(69187) <= 16338543;
srom_1(69188) <= 16503125;
srom_1(69189) <= 16629655;
srom_1(69190) <= 16717540;
srom_1(69191) <= 16766368;
srom_1(69192) <= 16775909;
srom_1(69193) <= 16746120;
srom_1(69194) <= 16677139;
srom_1(69195) <= 16569290;
srom_1(69196) <= 16423080;
srom_1(69197) <= 16239193;
srom_1(69198) <= 16018492;
srom_1(69199) <= 15762011;
srom_1(69200) <= 15470955;
srom_1(69201) <= 15146686;
srom_1(69202) <= 14790727;
srom_1(69203) <= 14404746;
srom_1(69204) <= 13990554;
srom_1(69205) <= 13550092;
srom_1(69206) <= 13085425;
srom_1(69207) <= 12598734;
srom_1(69208) <= 12092301;
srom_1(69209) <= 11568499;
srom_1(69210) <= 11029785;
srom_1(69211) <= 10478687;
srom_1(69212) <= 9917787;
srom_1(69213) <= 9349716;
srom_1(69214) <= 8777138;
srom_1(69215) <= 8202739;
srom_1(69216) <= 7629211;
srom_1(69217) <= 7059244;
srom_1(69218) <= 6495511;
srom_1(69219) <= 5940655;
srom_1(69220) <= 5397279;
srom_1(69221) <= 4867929;
srom_1(69222) <= 4355090;
srom_1(69223) <= 3861165;
srom_1(69224) <= 3388471;
srom_1(69225) <= 2939224;
srom_1(69226) <= 2515531;
srom_1(69227) <= 2119379;
srom_1(69228) <= 1752626;
srom_1(69229) <= 1416991;
srom_1(69230) <= 1114048;
srom_1(69231) <= 845219;
srom_1(69232) <= 611762;
srom_1(69233) <= 414775;
srom_1(69234) <= 255179;
srom_1(69235) <= 133723;
srom_1(69236) <= 50978;
srom_1(69237) <= 7330;
srom_1(69238) <= 2985;
srom_1(69239) <= 37964;
srom_1(69240) <= 112101;
srom_1(69241) <= 225050;
srom_1(69242) <= 376280;
srom_1(69243) <= 565083;
srom_1(69244) <= 790573;
srom_1(69245) <= 1051693;
srom_1(69246) <= 1347218;
srom_1(69247) <= 1675763;
srom_1(69248) <= 2035787;
srom_1(69249) <= 2425601;
srom_1(69250) <= 2843378;
srom_1(69251) <= 3287158;
srom_1(69252) <= 3754860;
srom_1(69253) <= 4244292;
srom_1(69254) <= 4753158;
srom_1(69255) <= 5279072;
srom_1(69256) <= 5819568;
srom_1(69257) <= 6372110;
srom_1(69258) <= 6934109;
srom_1(69259) <= 7502928;
srom_1(69260) <= 8075901;
srom_1(69261) <= 8650340;
srom_1(69262) <= 9223551;
srom_1(69263) <= 9792847;
srom_1(69264) <= 10355559;
srom_1(69265) <= 10909046;
srom_1(69266) <= 11450715;
srom_1(69267) <= 11978024;
srom_1(69268) <= 12488501;
srom_1(69269) <= 12979752;
srom_1(69270) <= 13449474;
srom_1(69271) <= 13895463;
srom_1(69272) <= 14315629;
srom_1(69273) <= 14708002;
srom_1(69274) <= 15070740;
srom_1(69275) <= 15402144;
srom_1(69276) <= 15700658;
srom_1(69277) <= 15964885;
srom_1(69278) <= 16193583;
srom_1(69279) <= 16385681;
srom_1(69280) <= 16540278;
srom_1(69281) <= 16656649;
srom_1(69282) <= 16734248;
srom_1(69283) <= 16772712;
srom_1(69284) <= 16771860;
srom_1(69285) <= 16731695;
srom_1(69286) <= 16652408;
srom_1(69287) <= 16534368;
srom_1(69288) <= 16378130;
srom_1(69289) <= 16184427;
srom_1(69290) <= 15954166;
srom_1(69291) <= 15688428;
srom_1(69292) <= 15388458;
srom_1(69293) <= 15055664;
srom_1(69294) <= 14691605;
srom_1(69295) <= 14297990;
srom_1(69296) <= 13876663;
srom_1(69297) <= 13429601;
srom_1(69298) <= 12958901;
srom_1(69299) <= 12466768;
srom_1(69300) <= 11955512;
srom_1(69301) <= 11427529;
srom_1(69302) <= 10885295;
srom_1(69303) <= 10331354;
srom_1(69304) <= 9768303;
srom_1(69305) <= 9198781;
srom_1(69306) <= 8625461;
srom_1(69307) <= 8051029;
srom_1(69308) <= 7478181;
srom_1(69309) <= 6909602;
srom_1(69310) <= 6347959;
srom_1(69311) <= 5795885;
srom_1(69312) <= 5255969;
srom_1(69313) <= 4730743;
srom_1(69314) <= 4222670;
srom_1(69315) <= 3734133;
srom_1(69316) <= 3267422;
srom_1(69317) <= 2824726;
srom_1(69318) <= 2408121;
srom_1(69319) <= 2019560;
srom_1(69320) <= 1660867;
srom_1(69321) <= 1333721;
srom_1(69322) <= 1039659;
srom_1(69323) <= 780058;
srom_1(69324) <= 556137;
srom_1(69325) <= 368944;
srom_1(69326) <= 219359;
srom_1(69327) <= 108082;
srom_1(69328) <= 35635;
srom_1(69329) <= 2358;
srom_1(69330) <= 8407;
srom_1(69331) <= 53754;
srom_1(69332) <= 138186;
srom_1(69333) <= 261307;
srom_1(69334) <= 422539;
srom_1(69335) <= 621128;
srom_1(69336) <= 856140;
srom_1(69337) <= 1126475;
srom_1(69338) <= 1430864;
srom_1(69339) <= 1767881;
srom_1(69340) <= 2135945;
srom_1(69341) <= 2533329;
srom_1(69342) <= 2958171;
srom_1(69343) <= 3408478;
srom_1(69344) <= 3882139;
srom_1(69345) <= 4376932;
srom_1(69346) <= 4890537;
srom_1(69347) <= 5420545;
srom_1(69348) <= 5964472;
srom_1(69349) <= 6519767;
srom_1(69350) <= 7083825;
srom_1(69351) <= 7654002;
srom_1(69352) <= 8227623;
srom_1(69353) <= 8802000;
srom_1(69354) <= 9374438;
srom_1(69355) <= 9942253;
srom_1(69356) <= 10502782;
srom_1(69357) <= 11053398;
srom_1(69358) <= 11591517;
srom_1(69359) <= 12114617;
srom_1(69360) <= 12620244;
srom_1(69361) <= 13106027;
srom_1(69362) <= 13569689;
srom_1(69363) <= 14009056;
srom_1(69364) <= 14422065;
srom_1(69365) <= 14806782;
srom_1(69366) <= 15161402;
srom_1(69367) <= 15484262;
srom_1(69368) <= 15773848;
srom_1(69369) <= 16028802;
srom_1(69370) <= 16247928;
srom_1(69371) <= 16430200;
srom_1(69372) <= 16574762;
srom_1(69373) <= 16680935;
srom_1(69374) <= 16748224;
srom_1(69375) <= 16776311;
srom_1(69376) <= 16765065;
srom_1(69377) <= 16714540;
srom_1(69378) <= 16624971;
srom_1(69379) <= 16496779;
srom_1(69380) <= 16330565;
srom_1(69381) <= 16127108;
srom_1(69382) <= 15887363;
srom_1(69383) <= 15612454;
srom_1(69384) <= 15303670;
srom_1(69385) <= 14962458;
srom_1(69386) <= 14590420;
srom_1(69387) <= 14189299;
srom_1(69388) <= 13760976;
srom_1(69389) <= 13307461;
srom_1(69390) <= 12830879;
srom_1(69391) <= 12333467;
srom_1(69392) <= 11817555;
srom_1(69393) <= 11285564;
srom_1(69394) <= 10739988;
srom_1(69395) <= 10183385;
srom_1(69396) <= 9618366;
srom_1(69397) <= 9047581;
srom_1(69398) <= 8473705;
srom_1(69399) <= 7899430;
srom_1(69400) <= 7327450;
srom_1(69401) <= 6760445;
srom_1(69402) <= 6201075;
srom_1(69403) <= 5651964;
srom_1(69404) <= 5115685;
srom_1(69405) <= 4594754;
srom_1(69406) <= 4091614;
srom_1(69407) <= 3608624;
srom_1(69408) <= 3148049;
srom_1(69409) <= 2712049;
srom_1(69410) <= 2302668;
srom_1(69411) <= 1921826;
srom_1(69412) <= 1571310;
srom_1(69413) <= 1252761;
srom_1(69414) <= 967676;
srom_1(69415) <= 717389;
srom_1(69416) <= 503076;
srom_1(69417) <= 325740;
srom_1(69418) <= 186214;
srom_1(69419) <= 85152;
srom_1(69420) <= 23027;
srom_1(69421) <= 132;
srom_1(69422) <= 16573;
srom_1(69423) <= 72274;
srom_1(69424) <= 166972;
srom_1(69425) <= 300225;
srom_1(69426) <= 471407;
srom_1(69427) <= 679715;
srom_1(69428) <= 924173;
srom_1(69429) <= 1203634;
srom_1(69430) <= 1516788;
srom_1(69431) <= 1862167;
srom_1(69432) <= 2238150;
srom_1(69433) <= 2642974;
srom_1(69434) <= 3074742;
srom_1(69435) <= 3531429;
srom_1(69436) <= 4010892;
srom_1(69437) <= 4510884;
srom_1(69438) <= 5029060;
srom_1(69439) <= 5562990;
srom_1(69440) <= 6110171;
srom_1(69441) <= 6668036;
srom_1(69442) <= 7233969;
srom_1(69443) <= 7805316;
srom_1(69444) <= 8379399;
srom_1(69445) <= 8953525;
srom_1(69446) <= 9525002;
srom_1(69447) <= 10091150;
srom_1(69448) <= 10649314;
srom_1(69449) <= 11196877;
srom_1(69450) <= 11731271;
srom_1(69451) <= 12249990;
srom_1(69452) <= 12750602;
srom_1(69453) <= 13230759;
srom_1(69454) <= 13688209;
srom_1(69455) <= 14120808;
srom_1(69456) <= 14526526;
srom_1(69457) <= 14903462;
srom_1(69458) <= 15249847;
srom_1(69459) <= 15564057;
srom_1(69460) <= 15844620;
srom_1(69461) <= 16090218;
srom_1(69462) <= 16299701;
srom_1(69463) <= 16472086;
srom_1(69464) <= 16606565;
srom_1(69465) <= 16702507;
srom_1(69466) <= 16759463;
srom_1(69467) <= 16777164;
srom_1(69468) <= 16755529;
srom_1(69469) <= 16694658;
srom_1(69470) <= 16594838;
srom_1(69471) <= 16456535;
srom_1(69472) <= 16280400;
srom_1(69473) <= 16067257;
srom_1(69474) <= 15818106;
srom_1(69475) <= 15534116;
srom_1(69476) <= 15216617;
srom_1(69477) <= 14867100;
srom_1(69478) <= 14487204;
srom_1(69479) <= 14078708;
srom_1(69480) <= 13643530;
srom_1(69481) <= 13183710;
srom_1(69482) <= 12701404;
srom_1(69483) <= 12198874;
srom_1(69484) <= 11678476;
srom_1(69485) <= 11142650;
srom_1(69486) <= 10593910;
srom_1(69487) <= 10034829;
srom_1(69488) <= 9468028;
srom_1(69489) <= 8896165;
srom_1(69490) <= 8321922;
srom_1(69491) <= 7747992;
srom_1(69492) <= 7177065;
srom_1(69493) <= 6611821;
srom_1(69494) <= 6054908;
srom_1(69495) <= 5508938;
srom_1(69496) <= 4976473;
srom_1(69497) <= 4460008;
srom_1(69498) <= 3961965;
srom_1(69499) <= 3484681;
srom_1(69500) <= 3030393;
srom_1(69501) <= 2601231;
srom_1(69502) <= 2199208;
srom_1(69503) <= 1826210;
srom_1(69504) <= 1483985;
srom_1(69505) <= 1174138;
srom_1(69506) <= 898122;
srom_1(69507) <= 657231;
srom_1(69508) <= 452596;
srom_1(69509) <= 285175;
srom_1(69510) <= 155754;
srom_1(69511) <= 64940;
srom_1(69512) <= 13158;
srom_1(69513) <= 652;
srom_1(69514) <= 27480;
srom_1(69515) <= 93516;
srom_1(69516) <= 198450;
srom_1(69517) <= 341791;
srom_1(69518) <= 522866;
srom_1(69519) <= 740826;
srom_1(69520) <= 994650;
srom_1(69521) <= 1283146;
srom_1(69522) <= 1604962;
srom_1(69523) <= 1958589;
srom_1(69524) <= 2342368;
srom_1(69525) <= 2754501;
srom_1(69526) <= 3193053;
srom_1(69527) <= 3655970;
srom_1(69528) <= 4141079;
srom_1(69529) <= 4646107;
srom_1(69530) <= 5168684;
srom_1(69531) <= 5706361;
srom_1(69532) <= 6256615;
srom_1(69533) <= 6816867;
srom_1(69534) <= 7384490;
srom_1(69535) <= 7956821;
srom_1(69536) <= 8531178;
srom_1(69537) <= 9104865;
srom_1(69538) <= 9675194;
srom_1(69539) <= 10239489;
srom_1(69540) <= 10795106;
srom_1(69541) <= 11339437;
srom_1(69542) <= 11869931;
srom_1(69543) <= 12384099;
srom_1(69544) <= 12879532;
srom_1(69545) <= 13353904;
srom_1(69546) <= 13804993;
srom_1(69547) <= 14230683;
srom_1(69548) <= 14628977;
srom_1(69549) <= 14998008;
srom_1(69550) <= 15336045;
srom_1(69551) <= 15641503;
srom_1(69552) <= 15912950;
srom_1(69553) <= 16149113;
srom_1(69554) <= 16348884;
srom_1(69555) <= 16511326;
srom_1(69556) <= 16635678;
srom_1(69557) <= 16721357;
srom_1(69558) <= 16767961;
srom_1(69559) <= 16775271;
srom_1(69560) <= 16743253;
srom_1(69561) <= 16672058;
srom_1(69562) <= 16562018;
srom_1(69563) <= 16413650;
srom_1(69564) <= 16227651;
srom_1(69565) <= 16004891;
srom_1(69566) <= 15746416;
srom_1(69567) <= 15453438;
srom_1(69568) <= 15127330;
srom_1(69569) <= 14769622;
srom_1(69570) <= 14381991;
srom_1(69571) <= 13966255;
srom_1(69572) <= 13524364;
srom_1(69573) <= 13058389;
srom_1(69574) <= 12570516;
srom_1(69575) <= 12063033;
srom_1(69576) <= 11538319;
srom_1(69577) <= 10998835;
srom_1(69578) <= 10447111;
srom_1(69579) <= 9885734;
srom_1(69580) <= 9317336;
srom_1(69581) <= 8744583;
srom_1(69582) <= 8170161;
srom_1(69583) <= 7596763;
srom_1(69584) <= 7027078;
srom_1(69585) <= 6463778;
srom_1(69586) <= 5909504;
srom_1(69587) <= 5366856;
srom_1(69588) <= 4838377;
srom_1(69589) <= 4326547;
srom_1(69590) <= 3833765;
srom_1(69591) <= 3362343;
srom_1(69592) <= 2914490;
srom_1(69593) <= 2492307;
srom_1(69594) <= 2097774;
srom_1(69595) <= 1732741;
srom_1(69596) <= 1398920;
srom_1(69597) <= 1097876;
srom_1(69598) <= 831020;
srom_1(69599) <= 599605;
srom_1(69600) <= 404714;
srom_1(69601) <= 247263;
srom_1(69602) <= 127990;
srom_1(69603) <= 47453;
srom_1(69604) <= 6031;
srom_1(69605) <= 3918;
srom_1(69606) <= 41124;
srom_1(69607) <= 117473;
srom_1(69608) <= 232609;
srom_1(69609) <= 385991;
srom_1(69610) <= 576900;
srom_1(69611) <= 804441;
srom_1(69612) <= 1067547;
srom_1(69613) <= 1364984;
srom_1(69614) <= 1695356;
srom_1(69615) <= 2057116;
srom_1(69616) <= 2448566;
srom_1(69617) <= 2867872;
srom_1(69618) <= 3313065;
srom_1(69619) <= 3782060;
srom_1(69620) <= 4272657;
srom_1(69621) <= 4782554;
srom_1(69622) <= 5309362;
srom_1(69623) <= 5850609;
srom_1(69624) <= 6403758;
srom_1(69625) <= 6966214;
srom_1(69626) <= 7535340;
srom_1(69627) <= 8108468;
srom_1(69628) <= 8682909;
srom_1(69629) <= 9255971;
srom_1(69630) <= 9824965;
srom_1(69631) <= 10387223;
srom_1(69632) <= 10940109;
srom_1(69633) <= 11481030;
srom_1(69634) <= 12007450;
srom_1(69635) <= 12516900;
srom_1(69636) <= 13006991;
srom_1(69637) <= 13475425;
srom_1(69638) <= 13920004;
srom_1(69639) <= 14338646;
srom_1(69640) <= 14729385;
srom_1(69641) <= 15090390;
srom_1(69642) <= 15419969;
srom_1(69643) <= 15716575;
srom_1(69644) <= 15978817;
srom_1(69645) <= 16205467;
srom_1(69646) <= 16395460;
srom_1(69647) <= 16547907;
srom_1(69648) <= 16662092;
srom_1(69649) <= 16737479;
srom_1(69650) <= 16773716;
srom_1(69651) <= 16770632;
srom_1(69652) <= 16728242;
srom_1(69653) <= 16646745;
srom_1(69654) <= 16526522;
srom_1(69655) <= 16368138;
srom_1(69656) <= 16172335;
srom_1(69657) <= 15940032;
srom_1(69658) <= 15672317;
srom_1(69659) <= 15370447;
srom_1(69660) <= 15035836;
srom_1(69661) <= 14670054;
srom_1(69662) <= 14274816;
srom_1(69663) <= 13851976;
srom_1(69664) <= 13403516;
srom_1(69665) <= 12931540;
srom_1(69666) <= 12438260;
srom_1(69667) <= 11925990;
srom_1(69668) <= 11397132;
srom_1(69669) <= 10854165;
srom_1(69670) <= 10299638;
srom_1(69671) <= 9736148;
srom_1(69672) <= 9166340;
srom_1(69673) <= 8592884;
srom_1(69674) <= 8018471;
srom_1(69675) <= 7445793;
srom_1(69676) <= 6877536;
srom_1(69677) <= 6316366;
srom_1(69678) <= 5764912;
srom_1(69679) <= 5225762;
srom_1(69680) <= 4701444;
srom_1(69681) <= 4194416;
srom_1(69682) <= 3707057;
srom_1(69683) <= 3241650;
srom_1(69684) <= 2800380;
srom_1(69685) <= 2385314;
srom_1(69686) <= 1998400;
srom_1(69687) <= 1641452;
srom_1(69688) <= 1316144;
srom_1(69689) <= 1024001;
srom_1(69690) <= 766393;
srom_1(69691) <= 544528;
srom_1(69692) <= 359447;
srom_1(69693) <= 212017;
srom_1(69694) <= 102930;
srom_1(69695) <= 32698;
srom_1(69696) <= 1649;
srom_1(69697) <= 9929;
srom_1(69698) <= 57500;
srom_1(69699) <= 144139;
srom_1(69700) <= 269439;
srom_1(69701) <= 432812;
srom_1(69702) <= 633492;
srom_1(69703) <= 870539;
srom_1(69704) <= 1142841;
srom_1(69705) <= 1449121;
srom_1(69706) <= 1787942;
srom_1(69707) <= 2157716;
srom_1(69708) <= 2556709;
srom_1(69709) <= 2983050;
srom_1(69710) <= 3434739;
srom_1(69711) <= 3909659;
srom_1(69712) <= 4405582;
srom_1(69713) <= 4920182;
srom_1(69714) <= 5451047;
srom_1(69715) <= 5995688;
srom_1(69716) <= 6551550;
srom_1(69717) <= 7116026;
srom_1(69718) <= 7686470;
srom_1(69719) <= 8260206;
srom_1(69720) <= 8834545;
srom_1(69721) <= 9406792;
srom_1(69722) <= 9974265;
srom_1(69723) <= 10534302;
srom_1(69724) <= 11084277;
srom_1(69725) <= 11621612;
srom_1(69726) <= 12143785;
srom_1(69727) <= 12648350;
srom_1(69728) <= 13132938;
srom_1(69729) <= 13595280;
srom_1(69730) <= 14033205;
srom_1(69731) <= 14444660;
srom_1(69732) <= 14827717;
srom_1(69733) <= 15180579;
srom_1(69734) <= 15501591;
srom_1(69735) <= 15789247;
srom_1(69736) <= 16042199;
srom_1(69737) <= 16259261;
srom_1(69738) <= 16439415;
srom_1(69739) <= 16581816;
srom_1(69740) <= 16685796;
srom_1(69741) <= 16750868;
srom_1(69742) <= 16776726;
srom_1(69743) <= 16763249;
srom_1(69744) <= 16710501;
srom_1(69745) <= 16618728;
srom_1(69746) <= 16488362;
srom_1(69747) <= 16320013;
srom_1(69748) <= 16114471;
srom_1(69749) <= 15872700;
srom_1(69750) <= 15595834;
srom_1(69751) <= 15285170;
srom_1(69752) <= 14942166;
srom_1(69753) <= 14568430;
srom_1(69754) <= 14165714;
srom_1(69755) <= 13735908;
srom_1(69756) <= 13281026;
srom_1(69757) <= 12803203;
srom_1(69758) <= 12304677;
srom_1(69759) <= 11787788;
srom_1(69760) <= 11254959;
srom_1(69761) <= 10708689;
srom_1(69762) <= 10151539;
srom_1(69763) <= 9586122;
srom_1(69764) <= 9015089;
srom_1(69765) <= 8441119;
srom_1(69766) <= 7866902;
srom_1(69767) <= 7295132;
srom_1(69768) <= 6728489;
srom_1(69769) <= 6169632;
srom_1(69770) <= 5621179;
srom_1(69771) <= 5085705;
srom_1(69772) <= 4565718;
srom_1(69773) <= 4063659;
srom_1(69774) <= 3581881;
srom_1(69775) <= 3122643;
srom_1(69776) <= 2688099;
srom_1(69777) <= 2280287;
srom_1(69778) <= 1901118;
srom_1(69779) <= 1552372;
srom_1(69780) <= 1235683;
srom_1(69781) <= 952537;
srom_1(69782) <= 704261;
srom_1(69783) <= 492020;
srom_1(69784) <= 316808;
srom_1(69785) <= 179448;
srom_1(69786) <= 80583;
srom_1(69787) <= 20678;
srom_1(69788) <= 12;
srom_1(69789) <= 18684;
srom_1(69790) <= 76605;
srom_1(69791) <= 173504;
srom_1(69792) <= 308926;
srom_1(69793) <= 482237;
srom_1(69794) <= 692623;
srom_1(69795) <= 939099;
srom_1(69796) <= 1220508;
srom_1(69797) <= 1535530;
srom_1(69798) <= 1882689;
srom_1(69799) <= 2260356;
srom_1(69800) <= 2666761;
srom_1(69801) <= 3099998;
srom_1(69802) <= 3558035;
srom_1(69803) <= 4038724;
srom_1(69804) <= 4539811;
srom_1(69805) <= 5058946;
srom_1(69806) <= 5593695;
srom_1(69807) <= 6141551;
srom_1(69808) <= 6699943;
srom_1(69809) <= 7266255;
srom_1(69810) <= 7837829;
srom_1(69811) <= 8411987;
srom_1(69812) <= 8986035;
srom_1(69813) <= 9557281;
srom_1(69814) <= 10123047;
srom_1(69815) <= 10680679;
srom_1(69816) <= 11227563;
srom_1(69817) <= 11761135;
srom_1(69818) <= 12278891;
srom_1(69819) <= 12778404;
srom_1(69820) <= 13257333;
srom_1(69821) <= 13713430;
srom_1(69822) <= 14144557;
srom_1(69823) <= 14548692;
srom_1(69824) <= 14923941;
srom_1(69825) <= 15268544;
srom_1(69826) <= 15580884;
srom_1(69827) <= 15859496;
srom_1(69828) <= 16103076;
srom_1(69829) <= 16310479;
srom_1(69830) <= 16480734;
srom_1(69831) <= 16613043;
srom_1(69832) <= 16706784;
srom_1(69833) <= 16761518;
srom_1(69834) <= 16776989;
srom_1(69835) <= 16753124;
srom_1(69836) <= 16690035;
srom_1(69837) <= 16588018;
srom_1(69838) <= 16447550;
srom_1(69839) <= 16269292;
srom_1(69840) <= 16054078;
srom_1(69841) <= 15802918;
srom_1(69842) <= 15516991;
srom_1(69843) <= 15197635;
srom_1(69844) <= 14846350;
srom_1(69845) <= 14464782;
srom_1(69846) <= 14054721;
srom_1(69847) <= 13618089;
srom_1(69848) <= 13156935;
srom_1(69849) <= 12673420;
srom_1(69850) <= 12169813;
srom_1(69851) <= 11648474;
srom_1(69852) <= 11111848;
srom_1(69853) <= 10562452;
srom_1(69854) <= 10002862;
srom_1(69855) <= 9435703;
srom_1(69856) <= 8863633;
srom_1(69857) <= 8289336;
srom_1(69858) <= 7715504;
srom_1(69859) <= 7144829;
srom_1(69860) <= 6579986;
srom_1(69861) <= 6023624;
srom_1(69862) <= 5478353;
srom_1(69863) <= 4946728;
srom_1(69864) <= 4431244;
srom_1(69865) <= 3934317;
srom_1(69866) <= 3458278;
srom_1(69867) <= 3005360;
srom_1(69868) <= 2577684;
srom_1(69869) <= 2177259;
srom_1(69870) <= 1805960;
srom_1(69871) <= 1465530;
srom_1(69872) <= 1157564;
srom_1(69873) <= 883508;
srom_1(69874) <= 644645;
srom_1(69875) <= 442096;
srom_1(69876) <= 276812;
srom_1(69877) <= 149566;
srom_1(69878) <= 60956;
srom_1(69879) <= 11397;
srom_1(69880) <= 1122;
srom_1(69881) <= 30178;
srom_1(69882) <= 98431;
srom_1(69883) <= 205558;
srom_1(69884) <= 351059;
srom_1(69885) <= 534250;
srom_1(69886) <= 754274;
srom_1(69887) <= 1010097;
srom_1(69888) <= 1300521;
srom_1(69889) <= 1624183;
srom_1(69890) <= 1979566;
srom_1(69891) <= 2365003;
srom_1(69892) <= 2778687;
srom_1(69893) <= 3218677;
srom_1(69894) <= 3682912;
srom_1(69895) <= 4169213;
srom_1(69896) <= 4675300;
srom_1(69897) <= 5198800;
srom_1(69898) <= 5737258;
srom_1(69899) <= 6288149;
srom_1(69900) <= 6848890;
srom_1(69901) <= 7416851;
srom_1(69902) <= 7989369;
srom_1(69903) <= 8563760;
srom_1(69904) <= 9137328;
srom_1(69905) <= 9707386;
srom_1(69906) <= 10271260;
srom_1(69907) <= 10826305;
srom_1(69908) <= 11369920;
srom_1(69909) <= 11899553;
srom_1(69910) <= 12412723;
srom_1(69911) <= 12907022;
srom_1(69912) <= 13380133;
srom_1(69913) <= 13829837;
srom_1(69914) <= 14254025;
srom_1(69915) <= 14650708;
srom_1(69916) <= 15018026;
srom_1(69917) <= 15354256;
srom_1(69918) <= 15657822;
srom_1(69919) <= 15927300;
srom_1(69920) <= 16161427;
srom_1(69921) <= 16359104;
srom_1(69922) <= 16519404;
srom_1(69923) <= 16641577;
srom_1(69924) <= 16725049;
srom_1(69925) <= 16769428;
srom_1(69926) <= 16774507;
srom_1(69927) <= 16740261;
srom_1(69928) <= 16666851;
srom_1(69929) <= 16554622;
srom_1(69930) <= 16404100;
srom_1(69931) <= 16215990;
srom_1(69932) <= 15991175;
srom_1(69933) <= 15730709;
srom_1(69934) <= 15435814;
srom_1(69935) <= 15107871;
srom_1(69936) <= 14748420;
srom_1(69937) <= 14359145;
srom_1(69938) <= 13941872;
srom_1(69939) <= 13498559;
srom_1(69940) <= 13031282;
srom_1(69941) <= 12542235;
srom_1(69942) <= 12033710;
srom_1(69943) <= 11508092;
srom_1(69944) <= 10967845;
srom_1(69945) <= 10415504;
srom_1(69946) <= 9853658;
srom_1(69947) <= 9284941;
srom_1(69948) <= 8712022;
srom_1(69949) <= 8137585;
srom_1(69950) <= 7564326;
srom_1(69951) <= 6994933;
srom_1(69952) <= 6432074;
srom_1(69953) <= 5878391;
srom_1(69954) <= 5336478;
srom_1(69955) <= 4808879;
srom_1(69956) <= 4298066;
srom_1(69957) <= 3806434;
srom_1(69958) <= 3336290;
srom_1(69959) <= 2889839;
srom_1(69960) <= 2469172;
srom_1(69961) <= 2076264;
srom_1(69962) <= 1712957;
srom_1(69963) <= 1380954;
srom_1(69964) <= 1081813;
srom_1(69965) <= 816935;
srom_1(69966) <= 587564;
srom_1(69967) <= 394775;
srom_1(69968) <= 239471;
srom_1(69969) <= 122381;
srom_1(69970) <= 44055;
srom_1(69971) <= 4859;
srom_1(69972) <= 4977;
srom_1(69973) <= 44409;
srom_1(69974) <= 122970;
srom_1(69975) <= 240292;
srom_1(69976) <= 395823;
srom_1(69977) <= 588835;
srom_1(69978) <= 818424;
srom_1(69979) <= 1083511;
srom_1(69980) <= 1382855;
srom_1(69981) <= 1715051;
srom_1(69982) <= 2078541;
srom_1(69983) <= 2471622;
srom_1(69984) <= 2892449;
srom_1(69985) <= 3339050;
srom_1(69986) <= 3809329;
srom_1(69987) <= 4301083;
srom_1(69988) <= 4812004;
srom_1(69989) <= 5339698;
srom_1(69990) <= 5881688;
srom_1(69991) <= 6435435;
srom_1(69992) <= 6998341;
srom_1(69993) <= 7567766;
srom_1(69994) <= 8141040;
srom_1(69995) <= 8715475;
srom_1(69996) <= 9288377;
srom_1(69997) <= 9857060;
srom_1(69998) <= 10418857;
srom_1(69999) <= 10971134;
srom_1(70000) <= 11511300;
srom_1(70001) <= 12036822;
srom_1(70002) <= 12545237;
srom_1(70003) <= 13034160;
srom_1(70004) <= 13501299;
srom_1(70005) <= 13944462;
srom_1(70006) <= 14361572;
srom_1(70007) <= 14750673;
srom_1(70008) <= 15109940;
srom_1(70009) <= 15437688;
srom_1(70010) <= 15732380;
srom_1(70011) <= 15992635;
srom_1(70012) <= 16217233;
srom_1(70013) <= 16405119;
srom_1(70014) <= 16555412;
srom_1(70015) <= 16667409;
srom_1(70016) <= 16740584;
srom_1(70017) <= 16774594;
srom_1(70018) <= 16769278;
srom_1(70019) <= 16724663;
srom_1(70020) <= 16640957;
srom_1(70021) <= 16518554;
srom_1(70022) <= 16358026;
srom_1(70023) <= 16160126;
srom_1(70024) <= 15925784;
srom_1(70025) <= 15656096;
srom_1(70026) <= 15352330;
srom_1(70027) <= 15015908;
srom_1(70028) <= 14648408;
srom_1(70029) <= 14251554;
srom_1(70030) <= 13827206;
srom_1(70031) <= 13377355;
srom_1(70032) <= 12904110;
srom_1(70033) <= 12409690;
srom_1(70034) <= 11896414;
srom_1(70035) <= 11366689;
srom_1(70036) <= 10822999;
srom_1(70037) <= 10267892;
srom_1(70038) <= 9703973;
srom_1(70039) <= 9133886;
srom_1(70040) <= 8560304;
srom_1(70041) <= 7985917;
srom_1(70042) <= 7413419;
srom_1(70043) <= 6845493;
srom_1(70044) <= 6284803;
srom_1(70045) <= 5733979;
srom_1(70046) <= 5195604;
srom_1(70047) <= 4672201;
srom_1(70048) <= 4166226;
srom_1(70049) <= 3680051;
srom_1(70050) <= 3215956;
srom_1(70051) <= 2776118;
srom_1(70052) <= 2362598;
srom_1(70053) <= 1977337;
srom_1(70054) <= 1622140;
srom_1(70055) <= 1298673;
srom_1(70056) <= 1008454;
srom_1(70057) <= 752842;
srom_1(70058) <= 533038;
srom_1(70059) <= 350070;
srom_1(70060) <= 204798;
srom_1(70061) <= 97903;
srom_1(70062) <= 29886;
srom_1(70063) <= 1066;
srom_1(70064) <= 11578;
srom_1(70065) <= 61372;
srom_1(70066) <= 150216;
srom_1(70067) <= 277693;
srom_1(70068) <= 443204;
srom_1(70069) <= 645974;
srom_1(70070) <= 885052;
srom_1(70071) <= 1159317;
srom_1(70072) <= 1467482;
srom_1(70073) <= 1808103;
srom_1(70074) <= 2179582;
srom_1(70075) <= 2580177;
srom_1(70076) <= 3008010;
srom_1(70077) <= 3461075;
srom_1(70078) <= 3937246;
srom_1(70079) <= 4434292;
srom_1(70080) <= 4949880;
srom_1(70081) <= 5481594;
srom_1(70082) <= 6026940;
srom_1(70083) <= 6583360;
srom_1(70084) <= 7148246;
srom_1(70085) <= 7718949;
srom_1(70086) <= 8292791;
srom_1(70087) <= 8867083;
srom_1(70088) <= 9439132;
srom_1(70089) <= 10006254;
srom_1(70090) <= 10565790;
srom_1(70091) <= 11115116;
srom_1(70092) <= 11651658;
srom_1(70093) <= 12172897;
srom_1(70094) <= 12676391;
srom_1(70095) <= 13159778;
srom_1(70096) <= 13620791;
srom_1(70097) <= 14057269;
srom_1(70098) <= 14467164;
srom_1(70099) <= 14848555;
srom_1(70100) <= 15199653;
srom_1(70101) <= 15518812;
srom_1(70102) <= 15804534;
srom_1(70103) <= 16055481;
srom_1(70104) <= 16270475;
srom_1(70105) <= 16448509;
srom_1(70106) <= 16588747;
srom_1(70107) <= 16690531;
srom_1(70108) <= 16753385;
srom_1(70109) <= 16777014;
srom_1(70110) <= 16761306;
srom_1(70111) <= 16706336;
srom_1(70112) <= 16612362;
srom_1(70113) <= 16479823;
srom_1(70114) <= 16309342;
srom_1(70115) <= 16101718;
srom_1(70116) <= 15857924;
srom_1(70117) <= 15579104;
srom_1(70118) <= 15266566;
srom_1(70119) <= 14921774;
srom_1(70120) <= 14546346;
srom_1(70121) <= 14142042;
srom_1(70122) <= 13710759;
srom_1(70123) <= 13254518;
srom_1(70124) <= 12775459;
srom_1(70125) <= 12275829;
srom_1(70126) <= 11757970;
srom_1(70127) <= 11224311;
srom_1(70128) <= 10677355;
srom_1(70129) <= 10119665;
srom_1(70130) <= 9553858;
srom_1(70131) <= 8982587;
srom_1(70132) <= 8408531;
srom_1(70133) <= 7834381;
srom_1(70134) <= 7262830;
srom_1(70135) <= 6696558;
srom_1(70136) <= 6138221;
srom_1(70137) <= 5590437;
srom_1(70138) <= 5055774;
srom_1(70139) <= 4536740;
srom_1(70140) <= 4035769;
srom_1(70141) <= 3555210;
srom_1(70142) <= 3097316;
srom_1(70143) <= 2664235;
srom_1(70144) <= 2257997;
srom_1(70145) <= 1880508;
srom_1(70146) <= 1533538;
srom_1(70147) <= 1218713;
srom_1(70148) <= 937511;
srom_1(70149) <= 691249;
srom_1(70150) <= 481083;
srom_1(70151) <= 307998;
srom_1(70152) <= 172805;
srom_1(70153) <= 76140;
srom_1(70154) <= 18454;
srom_1(70155) <= 19;
srom_1(70156) <= 20921;
srom_1(70157) <= 81062;
srom_1(70158) <= 180159;
srom_1(70159) <= 317749;
srom_1(70160) <= 493186;
srom_1(70161) <= 705648;
srom_1(70162) <= 954137;
srom_1(70163) <= 1237489;
srom_1(70164) <= 1554375;
srom_1(70165) <= 1903310;
srom_1(70166) <= 2282656;
srom_1(70167) <= 2690635;
srom_1(70168) <= 3125333;
srom_1(70169) <= 3584713;
srom_1(70170) <= 4066620;
srom_1(70171) <= 4568795;
srom_1(70172) <= 5088882;
srom_1(70173) <= 5624442;
srom_1(70174) <= 6172964;
srom_1(70175) <= 6731877;
srom_1(70176) <= 7298558;
srom_1(70177) <= 7870351;
srom_1(70178) <= 8444574;
srom_1(70179) <= 9018535;
srom_1(70180) <= 9589542;
srom_1(70181) <= 10154917;
srom_1(70182) <= 10712009;
srom_1(70183) <= 11258207;
srom_1(70184) <= 11790947;
srom_1(70185) <= 12307733;
srom_1(70186) <= 12806141;
srom_1(70187) <= 13283833;
srom_1(70188) <= 13738570;
srom_1(70189) <= 14168219;
srom_1(70190) <= 14570766;
srom_1(70191) <= 14944322;
srom_1(70192) <= 15287137;
srom_1(70193) <= 15597601;
srom_1(70194) <= 15874261;
srom_1(70195) <= 16115817;
srom_1(70196) <= 16321138;
srom_1(70197) <= 16489261;
srom_1(70198) <= 16619396;
srom_1(70199) <= 16710935;
srom_1(70200) <= 16763448;
srom_1(70201) <= 16776688;
srom_1(70202) <= 16750593;
srom_1(70203) <= 16685286;
srom_1(70204) <= 16581074;
srom_1(70205) <= 16438444;
srom_1(70206) <= 16258065;
srom_1(70207) <= 16040784;
srom_1(70208) <= 15787619;
srom_1(70209) <= 15499758;
srom_1(70210) <= 15178550;
srom_1(70211) <= 14825502;
srom_1(70212) <= 14442269;
srom_1(70213) <= 14030648;
srom_1(70214) <= 13592569;
srom_1(70215) <= 13130088;
srom_1(70216) <= 12645372;
srom_1(70217) <= 12140695;
srom_1(70218) <= 11618423;
srom_1(70219) <= 11081005;
srom_1(70220) <= 10530961;
srom_1(70221) <= 9970872;
srom_1(70222) <= 9403362;
srom_1(70223) <= 8831094;
srom_1(70224) <= 8256751;
srom_1(70225) <= 7683026;
srom_1(70226) <= 7112610;
srom_1(70227) <= 6548178;
srom_1(70228) <= 5992376;
srom_1(70229) <= 5447811;
srom_1(70230) <= 4917036;
srom_1(70231) <= 4402540;
srom_1(70232) <= 3906737;
srom_1(70233) <= 3431951;
srom_1(70234) <= 2980408;
srom_1(70235) <= 2554226;
srom_1(70236) <= 2155403;
srom_1(70237) <= 1785810;
srom_1(70238) <= 1447180;
srom_1(70239) <= 1141100;
srom_1(70240) <= 869007;
srom_1(70241) <= 632176;
srom_1(70242) <= 431717;
srom_1(70243) <= 268570;
srom_1(70244) <= 143502;
srom_1(70245) <= 57097;
srom_1(70246) <= 9762;
srom_1(70247) <= 1718;
srom_1(70248) <= 33003;
srom_1(70249) <= 103471;
srom_1(70250) <= 212790;
srom_1(70251) <= 360448;
srom_1(70252) <= 545753;
srom_1(70253) <= 767837;
srom_1(70254) <= 1025656;
srom_1(70255) <= 1318003;
srom_1(70256) <= 1643506;
srom_1(70257) <= 2000640;
srom_1(70258) <= 2387729;
srom_1(70259) <= 2802958;
srom_1(70260) <= 3244380;
srom_1(70261) <= 3709925;
srom_1(70262) <= 4197410;
srom_1(70263) <= 4704549;
srom_1(70264) <= 5228964;
srom_1(70265) <= 5768195;
srom_1(70266) <= 6319714;
srom_1(70267) <= 6880936;
srom_1(70268) <= 7449227;
srom_1(70269) <= 8021923;
srom_1(70270) <= 8596339;
srom_1(70271) <= 9169781;
srom_1(70272) <= 9739559;
srom_1(70273) <= 10303002;
srom_1(70274) <= 10857468;
srom_1(70275) <= 11400357;
srom_1(70276) <= 11929123;
srom_1(70277) <= 12441286;
srom_1(70278) <= 12934444;
srom_1(70279) <= 13406286;
srom_1(70280) <= 13854598;
srom_1(70281) <= 14277278;
srom_1(70282) <= 14672344;
srom_1(70283) <= 15037943;
srom_1(70284) <= 15372362;
srom_1(70285) <= 15674031;
srom_1(70286) <= 15941536;
srom_1(70287) <= 16173623;
srom_1(70288) <= 16369203;
srom_1(70289) <= 16527360;
srom_1(70290) <= 16647351;
srom_1(70291) <= 16728614;
srom_1(70292) <= 16770768;
srom_1(70293) <= 16773616;
srom_1(70294) <= 16737142;
srom_1(70295) <= 16661520;
srom_1(70296) <= 16547103;
srom_1(70297) <= 16394429;
srom_1(70298) <= 16204212;
srom_1(70299) <= 15977345;
srom_1(70300) <= 15714892;
srom_1(70301) <= 15418084;
srom_1(70302) <= 15088311;
srom_1(70303) <= 14727122;
srom_1(70304) <= 14336209;
srom_1(70305) <= 13917406;
srom_1(70306) <= 13472676;
srom_1(70307) <= 13004106;
srom_1(70308) <= 12513891;
srom_1(70309) <= 12004332;
srom_1(70310) <= 11477818;
srom_1(70311) <= 10936817;
srom_1(70312) <= 10383867;
srom_1(70313) <= 9821560;
srom_1(70314) <= 9252533;
srom_1(70315) <= 8679456;
srom_1(70316) <= 8105014;
srom_1(70317) <= 7531903;
srom_1(70318) <= 6962808;
srom_1(70319) <= 6400400;
srom_1(70320) <= 5847315;
srom_1(70321) <= 5306147;
srom_1(70322) <= 4779434;
srom_1(70323) <= 4269646;
srom_1(70324) <= 3779172;
srom_1(70325) <= 3310314;
srom_1(70326) <= 2865270;
srom_1(70327) <= 2446127;
srom_1(70328) <= 2054850;
srom_1(70329) <= 1693274;
srom_1(70330) <= 1363095;
srom_1(70331) <= 1065860;
srom_1(70332) <= 802965;
srom_1(70333) <= 575642;
srom_1(70334) <= 384956;
srom_1(70335) <= 231802;
srom_1(70336) <= 116898;
srom_1(70337) <= 40783;
srom_1(70338) <= 3813;
srom_1(70339) <= 6163;
srom_1(70340) <= 47821;
srom_1(70341) <= 128592;
srom_1(70342) <= 248097;
srom_1(70343) <= 405776;
srom_1(70344) <= 600888;
srom_1(70345) <= 832520;
srom_1(70346) <= 1099586;
srom_1(70347) <= 1400831;
srom_1(70348) <= 1734845;
srom_1(70349) <= 2100061;
srom_1(70350) <= 2494766;
srom_1(70351) <= 2917109;
srom_1(70352) <= 3365110;
srom_1(70353) <= 3836668;
srom_1(70354) <= 4329571;
srom_1(70355) <= 4841509;
srom_1(70356) <= 5370080;
srom_1(70357) <= 5912806;
srom_1(70358) <= 6467142;
srom_1(70359) <= 7030488;
srom_1(70360) <= 7600203;
srom_1(70361) <= 8173615;
srom_1(70362) <= 8748035;
srom_1(70363) <= 9320770;
srom_1(70364) <= 9889134;
srom_1(70365) <= 10450461;
srom_1(70366) <= 11002119;
srom_1(70367) <= 11541522;
srom_1(70368) <= 12066139;
srom_1(70369) <= 12573512;
srom_1(70370) <= 13061260;
srom_1(70371) <= 13527096;
srom_1(70372) <= 13968836;
srom_1(70373) <= 14384408;
srom_1(70374) <= 14771864;
srom_1(70375) <= 15129387;
srom_1(70376) <= 15455300;
srom_1(70377) <= 15748075;
srom_1(70378) <= 16006339;
srom_1(70379) <= 16228880;
srom_1(70380) <= 16414656;
srom_1(70381) <= 16562795;
srom_1(70382) <= 16672602;
srom_1(70383) <= 16743563;
srom_1(70384) <= 16775345;
srom_1(70385) <= 16767798;
srom_1(70386) <= 16720958;
srom_1(70387) <= 16635046;
srom_1(70388) <= 16510462;
srom_1(70389) <= 16347793;
srom_1(70390) <= 16147800;
srom_1(70391) <= 15911422;
srom_1(70392) <= 15639766;
srom_1(70393) <= 15334108;
srom_1(70394) <= 14995879;
srom_1(70395) <= 14626667;
srom_1(70396) <= 14228202;
srom_1(70397) <= 13802354;
srom_1(70398) <= 13351119;
srom_1(70399) <= 12876612;
srom_1(70400) <= 12381060;
srom_1(70401) <= 11866786;
srom_1(70402) <= 11336202;
srom_1(70403) <= 10791795;
srom_1(70404) <= 10236119;
srom_1(70405) <= 9671779;
srom_1(70406) <= 9101422;
srom_1(70407) <= 8527722;
srom_1(70408) <= 7953370;
srom_1(70409) <= 7381059;
srom_1(70410) <= 6813473;
srom_1(70411) <= 6253273;
srom_1(70412) <= 5703086;
srom_1(70413) <= 5165493;
srom_1(70414) <= 4643014;
srom_1(70415) <= 4138099;
srom_1(70416) <= 3653117;
srom_1(70417) <= 3190341;
srom_1(70418) <= 2751941;
srom_1(70419) <= 2339973;
srom_1(70420) <= 1956370;
srom_1(70421) <= 1602929;
srom_1(70422) <= 1281309;
srom_1(70423) <= 993018;
srom_1(70424) <= 739407;
srom_1(70425) <= 521666;
srom_1(70426) <= 340815;
srom_1(70427) <= 197703;
srom_1(70428) <= 93002;
srom_1(70429) <= 27201;
srom_1(70430) <= 610;
srom_1(70431) <= 13353;
srom_1(70432) <= 65370;
srom_1(70433) <= 156418;
srom_1(70434) <= 286069;
srom_1(70435) <= 453716;
srom_1(70436) <= 658573;
srom_1(70437) <= 899678;
srom_1(70438) <= 1175901;
srom_1(70439) <= 1485948;
srom_1(70440) <= 1828363;
srom_1(70441) <= 2201541;
srom_1(70442) <= 2603733;
srom_1(70443) <= 3033052;
srom_1(70444) <= 3487485;
srom_1(70445) <= 3964901;
srom_1(70446) <= 4463061;
srom_1(70447) <= 4979630;
srom_1(70448) <= 5512184;
srom_1(70449) <= 6058227;
srom_1(70450) <= 6615198;
srom_1(70451) <= 7180485;
srom_1(70452) <= 7751437;
srom_1(70453) <= 8325378;
srom_1(70454) <= 8899614;
srom_1(70455) <= 9471455;
srom_1(70456) <= 10038217;
srom_1(70457) <= 10597244;
srom_1(70458) <= 11145914;
srom_1(70459) <= 11681654;
srom_1(70460) <= 12201952;
srom_1(70461) <= 12704368;
srom_1(70462) <= 13186545;
srom_1(70463) <= 13646224;
srom_1(70464) <= 14081247;
srom_1(70465) <= 14489576;
srom_1(70466) <= 14869295;
srom_1(70467) <= 15218624;
srom_1(70468) <= 15535925;
srom_1(70469) <= 15819710;
srom_1(70470) <= 16068647;
srom_1(70471) <= 16281571;
srom_1(70472) <= 16457481;
srom_1(70473) <= 16595554;
srom_1(70474) <= 16695141;
srom_1(70475) <= 16755777;
srom_1(70476) <= 16777175;
srom_1(70477) <= 16759237;
srom_1(70478) <= 16702046;
srom_1(70479) <= 16605871;
srom_1(70480) <= 16471162;
srom_1(70481) <= 16298551;
srom_1(70482) <= 16088848;
srom_1(70483) <= 15843035;
srom_1(70484) <= 15562266;
srom_1(70485) <= 15247858;
srom_1(70486) <= 14901284;
srom_1(70487) <= 14524170;
srom_1(70488) <= 14118284;
srom_1(70489) <= 13685530;
srom_1(70490) <= 13227936;
srom_1(70491) <= 12747650;
srom_1(70492) <= 12246922;
srom_1(70493) <= 11728101;
srom_1(70494) <= 11193620;
srom_1(70495) <= 10645986;
srom_1(70496) <= 10087766;
srom_1(70497) <= 9521578;
srom_1(70498) <= 8950077;
srom_1(70499) <= 8375943;
srom_1(70500) <= 7801869;
srom_1(70501) <= 7230546;
srom_1(70502) <= 6664653;
srom_1(70503) <= 6106845;
srom_1(70504) <= 5559737;
srom_1(70505) <= 5025894;
srom_1(70506) <= 4507820;
srom_1(70507) <= 4007945;
srom_1(70508) <= 3528612;
srom_1(70509) <= 3072069;
srom_1(70510) <= 2640457;
srom_1(70511) <= 2235800;
srom_1(70512) <= 1859996;
srom_1(70513) <= 1514807;
srom_1(70514) <= 1201851;
srom_1(70515) <= 922597;
srom_1(70516) <= 678353;
srom_1(70517) <= 470265;
srom_1(70518) <= 299309;
srom_1(70519) <= 166287;
srom_1(70520) <= 71822;
srom_1(70521) <= 16357;
srom_1(70522) <= 152;
srom_1(70523) <= 23284;
srom_1(70524) <= 85644;
srom_1(70525) <= 186939;
srom_1(70526) <= 326694;
srom_1(70527) <= 504255;
srom_1(70528) <= 718788;
srom_1(70529) <= 969288;
srom_1(70530) <= 1254579;
srom_1(70531) <= 1573324;
srom_1(70532) <= 1924028;
srom_1(70533) <= 2305047;
srom_1(70534) <= 2714594;
srom_1(70535) <= 3150748;
srom_1(70536) <= 3611465;
srom_1(70537) <= 4094583;
srom_1(70538) <= 4597837;
srom_1(70539) <= 5118867;
srom_1(70540) <= 5655231;
srom_1(70541) <= 6204412;
srom_1(70542) <= 6763835;
srom_1(70543) <= 7330878;
srom_1(70544) <= 7902880;
srom_1(70545) <= 8477161;
srom_1(70546) <= 9051026;
srom_1(70547) <= 9621785;
srom_1(70548) <= 10186761;
srom_1(70549) <= 10743305;
srom_1(70550) <= 11288807;
srom_1(70551) <= 11820709;
srom_1(70552) <= 12336516;
srom_1(70553) <= 12833811;
srom_1(70554) <= 13310260;
srom_1(70555) <= 13763630;
srom_1(70556) <= 14191795;
srom_1(70557) <= 14592746;
srom_1(70558) <= 14964604;
srom_1(70559) <= 15305625;
srom_1(70560) <= 15614210;
srom_1(70561) <= 15888912;
srom_1(70562) <= 16128442;
srom_1(70563) <= 16331677;
srom_1(70564) <= 16497664;
srom_1(70565) <= 16625626;
srom_1(70566) <= 16714961;
srom_1(70567) <= 16765251;
srom_1(70568) <= 16776260;
srom_1(70569) <= 16747936;
srom_1(70570) <= 16680413;
srom_1(70571) <= 16574006;
srom_1(70572) <= 16429216;
srom_1(70573) <= 16246720;
srom_1(70574) <= 16027374;
srom_1(70575) <= 15772208;
srom_1(70576) <= 15482418;
srom_1(70577) <= 15159362;
srom_1(70578) <= 14804556;
srom_1(70579) <= 14419664;
srom_1(70580) <= 14006490;
srom_1(70581) <= 13566971;
srom_1(70582) <= 13103169;
srom_1(70583) <= 12617260;
srom_1(70584) <= 12111520;
srom_1(70585) <= 11588323;
srom_1(70586) <= 11050121;
srom_1(70587) <= 10499438;
srom_1(70588) <= 9938857;
srom_1(70589) <= 9371006;
srom_1(70590) <= 8798548;
srom_1(70591) <= 8224168;
srom_1(70592) <= 7650559;
srom_1(70593) <= 7080411;
srom_1(70594) <= 6516398;
srom_1(70595) <= 5961164;
srom_1(70596) <= 5417313;
srom_1(70597) <= 4887396;
srom_1(70598) <= 4373897;
srom_1(70599) <= 3879224;
srom_1(70600) <= 3405698;
srom_1(70601) <= 2955537;
srom_1(70602) <= 2530855;
srom_1(70603) <= 2133641;
srom_1(70604) <= 1765760;
srom_1(70605) <= 1428934;
srom_1(70606) <= 1124746;
srom_1(70607) <= 854620;
srom_1(70608) <= 619823;
srom_1(70609) <= 421457;
srom_1(70610) <= 260452;
srom_1(70611) <= 137562;
srom_1(70612) <= 53364;
srom_1(70613) <= 8254;
srom_1(70614) <= 2441;
srom_1(70615) <= 35954;
srom_1(70616) <= 108636;
srom_1(70617) <= 220145;
srom_1(70618) <= 369959;
srom_1(70619) <= 557375;
srom_1(70620) <= 781514;
srom_1(70621) <= 1041326;
srom_1(70622) <= 1335592;
srom_1(70623) <= 1662931;
srom_1(70624) <= 2021810;
srom_1(70625) <= 2410545;
srom_1(70626) <= 2827313;
srom_1(70627) <= 3270159;
srom_1(70628) <= 3737008;
srom_1(70629) <= 4225670;
srom_1(70630) <= 4733853;
srom_1(70631) <= 5259175;
srom_1(70632) <= 5799172;
srom_1(70633) <= 6351311;
srom_1(70634) <= 6913004;
srom_1(70635) <= 7481617;
srom_1(70636) <= 8054482;
srom_1(70637) <= 8628915;
srom_1(70638) <= 9202221;
srom_1(70639) <= 9771711;
srom_1(70640) <= 10334716;
srom_1(70641) <= 10888594;
srom_1(70642) <= 11430750;
srom_1(70643) <= 11958639;
srom_1(70644) <= 12469788;
srom_1(70645) <= 12961798;
srom_1(70646) <= 13432363;
srom_1(70647) <= 13879277;
srom_1(70648) <= 14300442;
srom_1(70649) <= 14693885;
srom_1(70650) <= 15057761;
srom_1(70651) <= 15390362;
srom_1(70652) <= 15690130;
srom_1(70653) <= 15955658;
srom_1(70654) <= 16185702;
srom_1(70655) <= 16379183;
srom_1(70656) <= 16535193;
srom_1(70657) <= 16653001;
srom_1(70658) <= 16732054;
srom_1(70659) <= 16771982;
srom_1(70660) <= 16772598;
srom_1(70661) <= 16733898;
srom_1(70662) <= 16656064;
srom_1(70663) <= 16539462;
srom_1(70664) <= 16384637;
srom_1(70665) <= 16192316;
srom_1(70666) <= 15963400;
srom_1(70667) <= 15698964;
srom_1(70668) <= 15400247;
srom_1(70669) <= 15068650;
srom_1(70670) <= 14705728;
srom_1(70671) <= 14313183;
srom_1(70672) <= 13892856;
srom_1(70673) <= 13446717;
srom_1(70674) <= 12976859;
srom_1(70675) <= 12485485;
srom_1(70676) <= 11974900;
srom_1(70677) <= 11447497;
srom_1(70678) <= 10905750;
srom_1(70679) <= 10352199;
srom_1(70680) <= 9789440;
srom_1(70681) <= 9220112;
srom_1(70682) <= 8646885;
srom_1(70683) <= 8072447;
srom_1(70684) <= 7499492;
srom_1(70685) <= 6930705;
srom_1(70686) <= 6368756;
srom_1(70687) <= 5816278;
srom_1(70688) <= 5275863;
srom_1(70689) <= 4750044;
srom_1(70690) <= 4241288;
srom_1(70691) <= 3751980;
srom_1(70692) <= 3284415;
srom_1(70693) <= 2840785;
srom_1(70694) <= 2423171;
srom_1(70695) <= 2033530;
srom_1(70696) <= 1673691;
srom_1(70697) <= 1345341;
srom_1(70698) <= 1050018;
srom_1(70699) <= 789109;
srom_1(70700) <= 563837;
srom_1(70701) <= 375257;
srom_1(70702) <= 224255;
srom_1(70703) <= 111539;
srom_1(70704) <= 37636;
srom_1(70705) <= 2894;
srom_1(70706) <= 7475;
srom_1(70707) <= 51359;
srom_1(70708) <= 134339;
srom_1(70709) <= 256025;
srom_1(70710) <= 415848;
srom_1(70711) <= 613059;
srom_1(70712) <= 846731;
srom_1(70713) <= 1115770;
srom_1(70714) <= 1418914;
srom_1(70715) <= 1754741;
srom_1(70716) <= 2121676;
srom_1(70717) <= 2517999;
srom_1(70718) <= 2941852;
srom_1(70719) <= 3391246;
srom_1(70720) <= 3864075;
srom_1(70721) <= 4358120;
srom_1(70722) <= 4871066;
srom_1(70723) <= 5400507;
srom_1(70724) <= 5943961;
srom_1(70725) <= 6498878;
srom_1(70726) <= 7062656;
srom_1(70727) <= 7632653;
srom_1(70728) <= 8206194;
srom_1(70729) <= 8780591;
srom_1(70730) <= 9353149;
srom_1(70731) <= 9921185;
srom_1(70732) <= 10482033;
srom_1(70733) <= 11033065;
srom_1(70734) <= 11571696;
srom_1(70735) <= 12095401;
srom_1(70736) <= 12601723;
srom_1(70737) <= 13088288;
srom_1(70738) <= 13552815;
srom_1(70739) <= 13993126;
srom_1(70740) <= 14407154;
srom_1(70741) <= 14792960;
srom_1(70742) <= 15148733;
srom_1(70743) <= 15472806;
srom_1(70744) <= 15763659;
srom_1(70745) <= 16019927;
srom_1(70746) <= 16240410;
srom_1(70747) <= 16424072;
srom_1(70748) <= 16570054;
srom_1(70749) <= 16677670;
srom_1(70750) <= 16746416;
srom_1(70751) <= 16775969;
srom_1(70752) <= 16766191;
srom_1(70753) <= 16717128;
srom_1(70754) <= 16629009;
srom_1(70755) <= 16502248;
srom_1(70756) <= 16337440;
srom_1(70757) <= 16135357;
srom_1(70758) <= 15896946;
srom_1(70759) <= 15623327;
srom_1(70760) <= 15315781;
srom_1(70761) <= 14975751;
srom_1(70762) <= 14604832;
srom_1(70763) <= 14204763;
srom_1(70764) <= 13777420;
srom_1(70765) <= 13324807;
srom_1(70766) <= 12849047;
srom_1(70767) <= 12352370;
srom_1(70768) <= 11837105;
srom_1(70769) <= 11305670;
srom_1(70770) <= 10760555;
srom_1(70771) <= 10204317;
srom_1(70772) <= 9639565;
srom_1(70773) <= 9068947;
srom_1(70774) <= 8495138;
srom_1(70775) <= 7920830;
srom_1(70776) <= 7348715;
srom_1(70777) <= 6781477;
srom_1(70778) <= 6221775;
srom_1(70779) <= 5672234;
srom_1(70780) <= 5135431;
srom_1(70781) <= 4613883;
srom_1(70782) <= 4110037;
srom_1(70783) <= 3626254;
srom_1(70784) <= 3164803;
srom_1(70785) <= 2727849;
srom_1(70786) <= 2317440;
srom_1(70787) <= 1935500;
srom_1(70788) <= 1583822;
srom_1(70789) <= 1264053;
srom_1(70790) <= 977694;
srom_1(70791) <= 726087;
srom_1(70792) <= 510412;
srom_1(70793) <= 331681;
srom_1(70794) <= 190732;
srom_1(70795) <= 88225;
srom_1(70796) <= 24642;
srom_1(70797) <= 280;
srom_1(70798) <= 15254;
srom_1(70799) <= 69493;
srom_1(70800) <= 162744;
srom_1(70801) <= 294568;
srom_1(70802) <= 464348;
srom_1(70803) <= 671288;
srom_1(70804) <= 914417;
srom_1(70805) <= 1192595;
srom_1(70806) <= 1504518;
srom_1(70807) <= 1848722;
srom_1(70808) <= 2223594;
srom_1(70809) <= 2627376;
srom_1(70810) <= 3058175;
srom_1(70811) <= 3513969;
srom_1(70812) <= 3992623;
srom_1(70813) <= 4491890;
srom_1(70814) <= 5009431;
srom_1(70815) <= 5542818;
srom_1(70816) <= 6089550;
srom_1(70817) <= 6647063;
srom_1(70818) <= 7212742;
srom_1(70819) <= 7783936;
srom_1(70820) <= 8357965;
srom_1(70821) <= 8932138;
srom_1(70822) <= 9503762;
srom_1(70823) <= 10070156;
srom_1(70824) <= 10628666;
srom_1(70825) <= 11176671;
srom_1(70826) <= 11711601;
srom_1(70827) <= 12230949;
srom_1(70828) <= 12732279;
srom_1(70829) <= 13213240;
srom_1(70830) <= 13671577;
srom_1(70831) <= 14105140;
srom_1(70832) <= 14511896;
srom_1(70833) <= 14889938;
srom_1(70834) <= 15237493;
srom_1(70835) <= 15552931;
srom_1(70836) <= 15834773;
srom_1(70837) <= 16081698;
srom_1(70838) <= 16292547;
srom_1(70839) <= 16466331;
srom_1(70840) <= 16602237;
srom_1(70841) <= 16699626;
srom_1(70842) <= 16758042;
srom_1(70843) <= 16777210;
srom_1(70844) <= 16757042;
srom_1(70845) <= 16697631;
srom_1(70846) <= 16599256;
srom_1(70847) <= 16462379;
srom_1(70848) <= 16287641;
srom_1(70849) <= 16075861;
srom_1(70850) <= 15828034;
srom_1(70851) <= 15545320;
srom_1(70852) <= 15229047;
srom_1(70853) <= 14880696;
srom_1(70854) <= 14501901;
srom_1(70855) <= 14094439;
srom_1(70856) <= 13660220;
srom_1(70857) <= 13201281;
srom_1(70858) <= 12719774;
srom_1(70859) <= 12217957;
srom_1(70860) <= 11698182;
srom_1(70861) <= 11162887;
srom_1(70862) <= 10614583;
srom_1(70863) <= 10055841;
srom_1(70864) <= 9489280;
srom_1(70865) <= 8917558;
srom_1(70866) <= 8343356;
srom_1(70867) <= 7769365;
srom_1(70868) <= 7198279;
srom_1(70869) <= 6632774;
srom_1(70870) <= 6075503;
srom_1(70871) <= 5529079;
srom_1(70872) <= 4996065;
srom_1(70873) <= 4478959;
srom_1(70874) <= 3980186;
srom_1(70875) <= 3502087;
srom_1(70876) <= 3046902;
srom_1(70877) <= 2616766;
srom_1(70878) <= 2213696;
srom_1(70879) <= 1839582;
srom_1(70880) <= 1496180;
srom_1(70881) <= 1185098;
srom_1(70882) <= 907795;
srom_1(70883) <= 665573;
srom_1(70884) <= 459567;
srom_1(70885) <= 290743;
srom_1(70886) <= 159892;
srom_1(70887) <= 67629;
srom_1(70888) <= 14386;
srom_1(70889) <= 412;
srom_1(70890) <= 25773;
srom_1(70891) <= 90351;
srom_1(70892) <= 193842;
srom_1(70893) <= 335761;
srom_1(70894) <= 515443;
srom_1(70895) <= 732044;
srom_1(70896) <= 984550;
srom_1(70897) <= 1271776;
srom_1(70898) <= 1592375;
srom_1(70899) <= 1944844;
srom_1(70900) <= 2327530;
srom_1(70901) <= 2738639;
srom_1(70902) <= 3176242;
srom_1(70903) <= 3638288;
srom_1(70904) <= 4122610;
srom_1(70905) <= 4626936;
srom_1(70906) <= 5148902;
srom_1(70907) <= 5686060;
srom_1(70908) <= 6235892;
srom_1(70909) <= 6795818;
srom_1(70910) <= 7363213;
srom_1(70911) <= 7935417;
srom_1(70912) <= 8509746;
srom_1(70913) <= 9083507;
srom_1(70914) <= 9654009;
srom_1(70915) <= 10218578;
srom_1(70916) <= 10774565;
srom_1(70917) <= 11319363;
srom_1(70918) <= 11850418;
srom_1(70919) <= 12365239;
srom_1(70920) <= 12861413;
srom_1(70921) <= 13336612;
srom_1(70922) <= 13788608;
srom_1(70923) <= 14215282;
srom_1(70924) <= 14614633;
srom_1(70925) <= 14984787;
srom_1(70926) <= 15324010;
srom_1(70927) <= 15630710;
srom_1(70928) <= 15903450;
srom_1(70929) <= 16140950;
srom_1(70930) <= 16342096;
srom_1(70931) <= 16505946;
srom_1(70932) <= 16631731;
srom_1(70933) <= 16718861;
srom_1(70934) <= 16766927;
srom_1(70935) <= 16775705;
srom_1(70936) <= 16745153;
srom_1(70937) <= 16675414;
srom_1(70938) <= 16566815;
srom_1(70939) <= 16419866;
srom_1(70940) <= 16235256;
srom_1(70941) <= 16013850;
srom_1(70942) <= 15756686;
srom_1(70943) <= 15464971;
srom_1(70944) <= 15140073;
srom_1(70945) <= 14783514;
srom_1(70946) <= 14396968;
srom_1(70947) <= 13982247;
srom_1(70948) <= 13541295;
srom_1(70949) <= 13076180;
srom_1(70950) <= 12589083;
srom_1(70951) <= 12082290;
srom_1(70952) <= 11558175;
srom_1(70953) <= 11019197;
srom_1(70954) <= 10467883;
srom_1(70955) <= 9906819;
srom_1(70956) <= 9338635;
srom_1(70957) <= 8765996;
srom_1(70958) <= 8191588;
srom_1(70959) <= 7618104;
srom_1(70960) <= 7048232;
srom_1(70961) <= 6484646;
srom_1(70962) <= 5929989;
srom_1(70963) <= 5386861;
srom_1(70964) <= 4857809;
srom_1(70965) <= 4345314;
srom_1(70966) <= 3851779;
srom_1(70967) <= 3379520;
srom_1(70968) <= 2930749;
srom_1(70969) <= 2507573;
srom_1(70970) <= 2111974;
srom_1(70971) <= 1745809;
srom_1(70972) <= 1410794;
srom_1(70973) <= 1108501;
srom_1(70974) <= 840346;
srom_1(70975) <= 607588;
srom_1(70976) <= 411318;
srom_1(70977) <= 252456;
srom_1(70978) <= 131747;
srom_1(70979) <= 49757;
srom_1(70980) <= 6871;
srom_1(70981) <= 3290;
srom_1(70982) <= 39031;
srom_1(70983) <= 113926;
srom_1(70984) <= 227623;
srom_1(70985) <= 379590;
srom_1(70986) <= 569114;
srom_1(70987) <= 795307;
srom_1(70988) <= 1057107;
srom_1(70989) <= 1353287;
srom_1(70990) <= 1682458;
srom_1(70991) <= 2043076;
srom_1(70992) <= 2433451;
srom_1(70993) <= 2851752;
srom_1(70994) <= 3296016;
srom_1(70995) <= 3764162;
srom_1(70996) <= 4253993;
srom_1(70997) <= 4763213;
srom_1(70998) <= 5289434;
srom_1(70999) <= 5830188;
srom_1(71000) <= 6382939;
srom_1(71001) <= 6945095;
srom_1(71002) <= 7514020;
srom_1(71003) <= 8087047;
srom_1(71004) <= 8661488;
srom_1(71005) <= 9234649;
srom_1(71006) <= 9803842;
srom_1(71007) <= 10366400;
srom_1(71008) <= 10919682;
srom_1(71009) <= 11461096;
srom_1(71010) <= 11988102;
srom_1(71011) <= 12498228;
srom_1(71012) <= 12989083;
srom_1(71013) <= 13458364;
srom_1(71014) <= 13903872;
srom_1(71015) <= 14323517;
srom_1(71016) <= 14715331;
srom_1(71017) <= 15077477;
srom_1(71018) <= 15408257;
srom_1(71019) <= 15706119;
srom_1(71020) <= 15969666;
srom_1(71021) <= 16197663;
srom_1(71022) <= 16389041;
srom_1(71023) <= 16542903;
srom_1(71024) <= 16658526;
srom_1(71025) <= 16735368;
srom_1(71026) <= 16773070;
srom_1(71027) <= 16771454;
srom_1(71028) <= 16730528;
srom_1(71029) <= 16650483;
srom_1(71030) <= 16531697;
srom_1(71031) <= 16374724;
srom_1(71032) <= 16180301;
srom_1(71033) <= 15949341;
srom_1(71034) <= 15682926;
srom_1(71035) <= 15382305;
srom_1(71036) <= 15048889;
srom_1(71037) <= 14684240;
srom_1(71038) <= 14290068;
srom_1(71039) <= 13868223;
srom_1(71040) <= 13420682;
srom_1(71041) <= 12949544;
srom_1(71042) <= 12457017;
srom_1(71043) <= 11945413;
srom_1(71044) <= 11417130;
srom_1(71045) <= 10874645;
srom_1(71046) <= 10320502;
srom_1(71047) <= 9757299;
srom_1(71048) <= 9187679;
srom_1(71049) <= 8614311;
srom_1(71050) <= 8039885;
srom_1(71051) <= 7467094;
srom_1(71052) <= 6898625;
srom_1(71053) <= 6337142;
srom_1(71054) <= 5785280;
srom_1(71055) <= 5245625;
srom_1(71056) <= 4720709;
srom_1(71057) <= 4212993;
srom_1(71058) <= 3724858;
srom_1(71059) <= 3258592;
srom_1(71060) <= 2816384;
srom_1(71061) <= 2400305;
srom_1(71062) <= 2012307;
srom_1(71063) <= 1654210;
srom_1(71064) <= 1327693;
srom_1(71065) <= 1034287;
srom_1(71066) <= 775368;
srom_1(71067) <= 552150;
srom_1(71068) <= 365680;
srom_1(71069) <= 216832;
srom_1(71070) <= 106305;
srom_1(71071) <= 34616;
srom_1(71072) <= 2101;
srom_1(71073) <= 8914;
srom_1(71074) <= 55022;
srom_1(71075) <= 140209;
srom_1(71076) <= 264076;
srom_1(71077) <= 426042;
srom_1(71078) <= 625346;
srom_1(71079) <= 861056;
srom_1(71080) <= 1132064;
srom_1(71081) <= 1437101;
srom_1(71082) <= 1774736;
srom_1(71083) <= 2143386;
srom_1(71084) <= 2541321;
srom_1(71085) <= 2966677;
srom_1(71086) <= 3417458;
srom_1(71087) <= 3891550;
srom_1(71088) <= 4386731;
srom_1(71089) <= 4900677;
srom_1(71090) <= 5430980;
srom_1(71091) <= 5975152;
srom_1(71092) <= 6530642;
srom_1(71093) <= 7094844;
srom_1(71094) <= 7665113;
srom_1(71095) <= 8238775;
srom_1(71096) <= 8813140;
srom_1(71097) <= 9385513;
srom_1(71098) <= 9953212;
srom_1(71099) <= 10513574;
srom_1(71100) <= 11063971;
srom_1(71101) <= 11601823;
srom_1(71102) <= 12124607;
srom_1(71103) <= 12629871;
srom_1(71104) <= 13115246;
srom_1(71105) <= 13578457;
srom_1(71106) <= 14017331;
srom_1(71107) <= 14429809;
srom_1(71108) <= 14813959;
srom_1(71109) <= 15167977;
srom_1(71110) <= 15490205;
srom_1(71111) <= 15779131;
srom_1(71112) <= 16033400;
srom_1(71113) <= 16251821;
srom_1(71114) <= 16433368;
srom_1(71115) <= 16577190;
srom_1(71116) <= 16682613;
srom_1(71117) <= 16749143;
srom_1(71118) <= 16776467;
srom_1(71119) <= 16764458;
srom_1(71120) <= 16713172;
srom_1(71121) <= 16622848;
srom_1(71122) <= 16493912;
srom_1(71123) <= 16326967;
srom_1(71124) <= 16122796;
srom_1(71125) <= 15882357;
srom_1(71126) <= 15606778;
srom_1(71127) <= 15297350;
srom_1(71128) <= 14955524;
srom_1(71129) <= 14582904;
srom_1(71130) <= 14181236;
srom_1(71131) <= 13752405;
srom_1(71132) <= 13298422;
srom_1(71133) <= 12821414;
srom_1(71134) <= 12323620;
srom_1(71135) <= 11807373;
srom_1(71136) <= 11275094;
srom_1(71137) <= 10729279;
srom_1(71138) <= 10172488;
srom_1(71139) <= 9607332;
srom_1(71140) <= 9036461;
srom_1(71141) <= 8462552;
srom_1(71142) <= 7888296;
srom_1(71143) <= 7316386;
srom_1(71144) <= 6749505;
srom_1(71145) <= 6190309;
srom_1(71146) <= 5641423;
srom_1(71147) <= 5105418;
srom_1(71148) <= 4584810;
srom_1(71149) <= 4082039;
srom_1(71150) <= 3599463;
srom_1(71151) <= 3139345;
srom_1(71152) <= 2703842;
srom_1(71153) <= 2294997;
srom_1(71154) <= 1914728;
srom_1(71155) <= 1564816;
srom_1(71156) <= 1246904;
srom_1(71157) <= 962482;
srom_1(71158) <= 712883;
srom_1(71159) <= 499278;
srom_1(71160) <= 322669;
srom_1(71161) <= 183884;
srom_1(71162) <= 83574;
srom_1(71163) <= 22209;
srom_1(71164) <= 77;
srom_1(71165) <= 17281;
srom_1(71166) <= 73742;
srom_1(71167) <= 169194;
srom_1(71168) <= 303189;
srom_1(71169) <= 475100;
srom_1(71170) <= 684120;
srom_1(71171) <= 929269;
srom_1(71172) <= 1209397;
srom_1(71173) <= 1523191;
srom_1(71174) <= 1869180;
srom_1(71175) <= 2245740;
srom_1(71176) <= 2651106;
srom_1(71177) <= 3083377;
srom_1(71178) <= 3540527;
srom_1(71179) <= 4020411;
srom_1(71180) <= 4520778;
srom_1(71181) <= 5039283;
srom_1(71182) <= 5573495;
srom_1(71183) <= 6120907;
srom_1(71184) <= 6678954;
srom_1(71185) <= 7245017;
srom_1(71186) <= 7816443;
srom_1(71187) <= 8390553;
srom_1(71188) <= 8964653;
srom_1(71189) <= 9536052;
srom_1(71190) <= 10102070;
srom_1(71191) <= 10660053;
srom_1(71192) <= 11207385;
srom_1(71193) <= 11741498;
srom_1(71194) <= 12259888;
srom_1(71195) <= 12760125;
srom_1(71196) <= 13239862;
srom_1(71197) <= 13696850;
srom_1(71198) <= 14128946;
srom_1(71199) <= 14534123;
srom_1(71200) <= 14910482;
srom_1(71201) <= 15256258;
srom_1(71202) <= 15569828;
srom_1(71203) <= 15849724;
srom_1(71204) <= 16094632;
srom_1(71205) <= 16303404;
srom_1(71206) <= 16475060;
srom_1(71207) <= 16608796;
srom_1(71208) <= 16703985;
srom_1(71209) <= 16760181;
srom_1(71210) <= 16777119;
srom_1(71211) <= 16754720;
srom_1(71212) <= 16693090;
srom_1(71213) <= 16592517;
srom_1(71214) <= 16453474;
srom_1(71215) <= 16276611;
srom_1(71216) <= 16062759;
srom_1(71217) <= 15812920;
srom_1(71218) <= 15528266;
srom_1(71219) <= 15210132;
srom_1(71220) <= 14860009;
srom_1(71221) <= 14479540;
srom_1(71222) <= 14070508;
srom_1(71223) <= 13634832;
srom_1(71224) <= 13174554;
srom_1(71225) <= 12691833;
srom_1(71226) <= 12188933;
srom_1(71227) <= 11668212;
srom_1(71228) <= 11132112;
srom_1(71229) <= 10583147;
srom_1(71230) <= 10023891;
srom_1(71231) <= 9456966;
srom_1(71232) <= 8885031;
srom_1(71233) <= 8310769;
srom_1(71234) <= 7736871;
srom_1(71235) <= 7166030;
srom_1(71236) <= 6600922;
srom_1(71237) <= 6044196;
srom_1(71238) <= 5498465;
srom_1(71239) <= 4966286;
srom_1(71240) <= 4450156;
srom_1(71241) <= 3952495;
srom_1(71242) <= 3475636;
srom_1(71243) <= 3021815;
srom_1(71244) <= 2593162;
srom_1(71245) <= 2191685;
srom_1(71246) <= 1819268;
srom_1(71247) <= 1477656;
srom_1(71248) <= 1168453;
srom_1(71249) <= 893107;
srom_1(71250) <= 652910;
srom_1(71251) <= 448989;
srom_1(71252) <= 282299;
srom_1(71253) <= 153622;
srom_1(71254) <= 63562;
srom_1(71255) <= 12541;
srom_1(71256) <= 799;
srom_1(71257) <= 28389;
srom_1(71258) <= 95184;
srom_1(71259) <= 200869;
srom_1(71260) <= 344949;
srom_1(71261) <= 526749;
srom_1(71262) <= 745416;
srom_1(71263) <= 999924;
srom_1(71264) <= 1289081;
srom_1(71265) <= 1611529;
srom_1(71266) <= 1965758;
srom_1(71267) <= 2350105;
srom_1(71268) <= 2762769;
srom_1(71269) <= 3201815;
srom_1(71270) <= 3665183;
srom_1(71271) <= 4150701;
srom_1(71272) <= 4656092;
srom_1(71273) <= 5178986;
srom_1(71274) <= 5716931;
srom_1(71275) <= 6267405;
srom_1(71276) <= 6827825;
srom_1(71277) <= 7395565;
srom_1(71278) <= 7967961;
srom_1(71279) <= 8542330;
srom_1(71280) <= 9115978;
srom_1(71281) <= 9686215;
srom_1(71282) <= 10250367;
srom_1(71283) <= 10805788;
srom_1(71284) <= 11349875;
srom_1(71285) <= 11880075;
srom_1(71286) <= 12393903;
srom_1(71287) <= 12888948;
srom_1(71288) <= 13362890;
srom_1(71289) <= 13813506;
srom_1(71290) <= 14238682;
srom_1(71291) <= 14636425;
srom_1(71292) <= 15004871;
srom_1(71293) <= 15342290;
srom_1(71294) <= 15647101;
srom_1(71295) <= 15917874;
srom_1(71296) <= 16153340;
srom_1(71297) <= 16352395;
srom_1(71298) <= 16514105;
srom_1(71299) <= 16637711;
srom_1(71300) <= 16722635;
srom_1(71301) <= 16768477;
srom_1(71302) <= 16775024;
srom_1(71303) <= 16742243;
srom_1(71304) <= 16670290;
srom_1(71305) <= 16559501;
srom_1(71306) <= 16410395;
srom_1(71307) <= 16223673;
srom_1(71308) <= 16000210;
srom_1(71309) <= 15741053;
srom_1(71310) <= 15447417;
srom_1(71311) <= 15120681;
srom_1(71312) <= 14762376;
srom_1(71313) <= 14374182;
srom_1(71314) <= 13957919;
srom_1(71315) <= 13515540;
srom_1(71316) <= 13049119;
srom_1(71317) <= 12560844;
srom_1(71318) <= 12053003;
srom_1(71319) <= 11527979;
srom_1(71320) <= 10988233;
srom_1(71321) <= 10436296;
srom_1(71322) <= 9874758;
srom_1(71323) <= 9306250;
srom_1(71324) <= 8733439;
srom_1(71325) <= 8159011;
srom_1(71326) <= 7585659;
srom_1(71327) <= 7016073;
srom_1(71328) <= 6452924;
srom_1(71329) <= 5898851;
srom_1(71330) <= 5356453;
srom_1(71331) <= 4828275;
srom_1(71332) <= 4316792;
srom_1(71333) <= 3824403;
srom_1(71334) <= 3353417;
srom_1(71335) <= 2906043;
srom_1(71336) <= 2484379;
srom_1(71337) <= 2090402;
srom_1(71338) <= 1725959;
srom_1(71339) <= 1392759;
srom_1(71340) <= 1092366;
srom_1(71341) <= 826187;
srom_1(71342) <= 595470;
srom_1(71343) <= 401299;
srom_1(71344) <= 244583;
srom_1(71345) <= 126056;
srom_1(71346) <= 46276;
srom_1(71347) <= 5616;
srom_1(71348) <= 4266;
srom_1(71349) <= 42234;
srom_1(71350) <= 119341;
srom_1(71351) <= 235225;
srom_1(71352) <= 389343;
srom_1(71353) <= 580972;
srom_1(71354) <= 809214;
srom_1(71355) <= 1072998;
srom_1(71356) <= 1371088;
srom_1(71357) <= 1702086;
srom_1(71358) <= 2064438;
srom_1(71359) <= 2456447;
srom_1(71360) <= 2876274;
srom_1(71361) <= 3321950;
srom_1(71362) <= 3791386;
srom_1(71363) <= 4282379;
srom_1(71364) <= 4792628;
srom_1(71365) <= 5319739;
srom_1(71366) <= 5861242;
srom_1(71367) <= 6414596;
srom_1(71368) <= 6977207;
srom_1(71369) <= 7546437;
srom_1(71370) <= 8119616;
srom_1(71371) <= 8694056;
srom_1(71372) <= 9267064;
srom_1(71373) <= 9835952;
srom_1(71374) <= 10398054;
srom_1(71375) <= 10950732;
srom_1(71376) <= 11491396;
srom_1(71377) <= 12017510;
srom_1(71378) <= 12526606;
srom_1(71379) <= 13016298;
srom_1(71380) <= 13484289;
srom_1(71381) <= 13928385;
srom_1(71382) <= 14346503;
srom_1(71383) <= 14736682;
srom_1(71384) <= 15097093;
srom_1(71385) <= 15426045;
srom_1(71386) <= 15721997;
srom_1(71387) <= 15983560;
srom_1(71388) <= 16209507;
srom_1(71389) <= 16398779;
srom_1(71390) <= 16550490;
srom_1(71391) <= 16663926;
srom_1(71392) <= 16738556;
srom_1(71393) <= 16774031;
srom_1(71394) <= 16770183;
srom_1(71395) <= 16727031;
srom_1(71396) <= 16644778;
srom_1(71397) <= 16523809;
srom_1(71398) <= 16364690;
srom_1(71399) <= 16168170;
srom_1(71400) <= 15935168;
srom_1(71401) <= 15666778;
srom_1(71402) <= 15364258;
srom_1(71403) <= 15029026;
srom_1(71404) <= 14662656;
srom_1(71405) <= 14266864;
srom_1(71406) <= 13843507;
srom_1(71407) <= 13394570;
srom_1(71408) <= 12922159;
srom_1(71409) <= 12428488;
srom_1(71410) <= 11915873;
srom_1(71411) <= 11386717;
srom_1(71412) <= 10843502;
srom_1(71413) <= 10288775;
srom_1(71414) <= 9725138;
srom_1(71415) <= 9155233;
srom_1(71416) <= 8581733;
srom_1(71417) <= 8007328;
srom_1(71418) <= 7434711;
srom_1(71419) <= 6866566;
srom_1(71420) <= 6305559;
srom_1(71421) <= 5754320;
srom_1(71422) <= 5215435;
srom_1(71423) <= 4691429;
srom_1(71424) <= 4184761;
srom_1(71425) <= 3697806;
srom_1(71426) <= 3232847;
srom_1(71427) <= 2792066;
srom_1(71428) <= 2377529;
srom_1(71429) <= 1991180;
srom_1(71430) <= 1634831;
srom_1(71431) <= 1310152;
srom_1(71432) <= 1018667;
srom_1(71433) <= 761742;
srom_1(71434) <= 540582;
srom_1(71435) <= 356224;
srom_1(71436) <= 209532;
srom_1(71437) <= 101196;
srom_1(71438) <= 31721;
srom_1(71439) <= 1435;
srom_1(71440) <= 10479;
srom_1(71441) <= 58812;
srom_1(71442) <= 146205;
srom_1(71443) <= 272250;
srom_1(71444) <= 436355;
srom_1(71445) <= 637751;
srom_1(71446) <= 875494;
srom_1(71447) <= 1148468;
srom_1(71448) <= 1455394;
srom_1(71449) <= 1794831;
srom_1(71450) <= 2165190;
srom_1(71451) <= 2564732;
srom_1(71452) <= 2991584;
srom_1(71453) <= 3443745;
srom_1(71454) <= 3919093;
srom_1(71455) <= 4415401;
srom_1(71456) <= 4930341;
srom_1(71457) <= 5461498;
srom_1(71458) <= 6006380;
srom_1(71459) <= 6562434;
srom_1(71460) <= 7127052;
srom_1(71461) <= 7697585;
srom_1(71462) <= 8271359;
srom_1(71463) <= 8845683;
srom_1(71464) <= 9417863;
srom_1(71465) <= 9985216;
srom_1(71466) <= 10545083;
srom_1(71467) <= 11094837;
srom_1(71468) <= 11631901;
srom_1(71469) <= 12153756;
srom_1(71470) <= 12657954;
srom_1(71471) <= 13142133;
srom_1(71472) <= 13604020;
srom_1(71473) <= 14041451;
srom_1(71474) <= 14452373;
srom_1(71475) <= 14834860;
srom_1(71476) <= 15187119;
srom_1(71477) <= 15507497;
srom_1(71478) <= 15794492;
srom_1(71479) <= 16046758;
srom_1(71480) <= 16263113;
srom_1(71481) <= 16442541;
srom_1(71482) <= 16584202;
srom_1(71483) <= 16687431;
srom_1(71484) <= 16751744;
srom_1(71485) <= 16776839;
srom_1(71486) <= 16762598;
srom_1(71487) <= 16709090;
srom_1(71488) <= 16616563;
srom_1(71489) <= 16485453;
srom_1(71490) <= 16316374;
srom_1(71491) <= 16110119;
srom_1(71492) <= 15867656;
srom_1(71493) <= 15590120;
srom_1(71494) <= 15278814;
srom_1(71495) <= 14935197;
srom_1(71496) <= 14560882;
srom_1(71497) <= 14157622;
srom_1(71498) <= 13727309;
srom_1(71499) <= 13271962;
srom_1(71500) <= 12793714;
srom_1(71501) <= 12294810;
srom_1(71502) <= 11777588;
srom_1(71503) <= 11244474;
srom_1(71504) <= 10697968;
srom_1(71505) <= 10140632;
srom_1(71506) <= 9575081;
srom_1(71507) <= 9003966;
srom_1(71508) <= 8429965;
srom_1(71509) <= 7855770;
srom_1(71510) <= 7284074;
srom_1(71511) <= 6717558;
srom_1(71512) <= 6158877;
srom_1(71513) <= 5610653;
srom_1(71514) <= 5075455;
srom_1(71515) <= 4555794;
srom_1(71516) <= 4054106;
srom_1(71517) <= 3572744;
srom_1(71518) <= 3113965;
srom_1(71519) <= 2679921;
srom_1(71520) <= 2272647;
srom_1(71521) <= 1894053;
srom_1(71522) <= 1545914;
srom_1(71523) <= 1229863;
srom_1(71524) <= 947381;
srom_1(71525) <= 699794;
srom_1(71526) <= 488263;
srom_1(71527) <= 313779;
srom_1(71528) <= 177160;
srom_1(71529) <= 79048;
srom_1(71530) <= 19902;
srom_1(71531) <= 0;
srom_1(71532) <= 19435;
srom_1(71533) <= 78116;
srom_1(71534) <= 175768;
srom_1(71535) <= 311932;
srom_1(71536) <= 485971;
srom_1(71537) <= 697068;
srom_1(71538) <= 944233;
srom_1(71539) <= 1226308;
srom_1(71540) <= 1541969;
srom_1(71541) <= 1889736;
srom_1(71542) <= 2267978;
srom_1(71543) <= 2674923;
srom_1(71544) <= 3108660;
srom_1(71545) <= 3567158;
srom_1(71546) <= 4048264;
srom_1(71547) <= 4549724;
srom_1(71548) <= 5069186;
srom_1(71549) <= 5604214;
srom_1(71550) <= 6152299;
srom_1(71551) <= 6710870;
srom_1(71552) <= 7277309;
srom_1(71553) <= 7848960;
srom_1(71554) <= 8423140;
srom_1(71555) <= 8997159;
srom_1(71556) <= 9568325;
srom_1(71557) <= 10133958;
srom_1(71558) <= 10691406;
srom_1(71559) <= 11238056;
srom_1(71560) <= 11771344;
srom_1(71561) <= 12288769;
srom_1(71562) <= 12787905;
srom_1(71563) <= 13266411;
srom_1(71564) <= 13722044;
srom_1(71565) <= 14152666;
srom_1(71566) <= 14556258;
srom_1(71567) <= 14930928;
srom_1(71568) <= 15274919;
srom_1(71569) <= 15586618;
srom_1(71570) <= 15864562;
srom_1(71571) <= 16107450;
srom_1(71572) <= 16314141;
srom_1(71573) <= 16483666;
srom_1(71574) <= 16615231;
srom_1(71575) <= 16708219;
srom_1(71576) <= 16762193;
srom_1(71577) <= 16776900;
srom_1(71578) <= 16752272;
srom_1(71579) <= 16688424;
srom_1(71580) <= 16585655;
srom_1(71581) <= 16444447;
srom_1(71582) <= 16265463;
srom_1(71583) <= 16049541;
srom_1(71584) <= 15797695;
srom_1(71585) <= 15511104;
srom_1(71586) <= 15191114;
srom_1(71587) <= 14839225;
srom_1(71588) <= 14457087;
srom_1(71589) <= 14046491;
srom_1(71590) <= 13609364;
srom_1(71591) <= 13147754;
srom_1(71592) <= 12663828;
srom_1(71593) <= 12159853;
srom_1(71594) <= 11638194;
srom_1(71595) <= 11101296;
srom_1(71596) <= 10551678;
srom_1(71597) <= 9991916;
srom_1(71598) <= 9424635;
srom_1(71599) <= 8852497;
srom_1(71600) <= 8278183;
srom_1(71601) <= 7704387;
srom_1(71602) <= 7133799;
srom_1(71603) <= 6569096;
srom_1(71604) <= 6012925;
srom_1(71605) <= 5467894;
srom_1(71606) <= 4936560;
srom_1(71607) <= 4421413;
srom_1(71608) <= 3924870;
srom_1(71609) <= 3449259;
srom_1(71610) <= 2996810;
srom_1(71611) <= 2569645;
srom_1(71612) <= 2169768;
srom_1(71613) <= 1799052;
srom_1(71614) <= 1459238;
srom_1(71615) <= 1151917;
srom_1(71616) <= 878532;
srom_1(71617) <= 640364;
srom_1(71618) <= 438530;
srom_1(71619) <= 273977;
srom_1(71620) <= 147476;
srom_1(71621) <= 59621;
srom_1(71622) <= 10823;
srom_1(71623) <= 1312;
srom_1(71624) <= 31131;
srom_1(71625) <= 100141;
srom_1(71626) <= 208019;
srom_1(71627) <= 354259;
srom_1(71628) <= 538174;
srom_1(71629) <= 758903;
srom_1(71630) <= 1015410;
srom_1(71631) <= 1306492;
srom_1(71632) <= 1630785;
srom_1(71633) <= 1986768;
srom_1(71634) <= 2372771;
srom_1(71635) <= 2786984;
srom_1(71636) <= 3227466;
srom_1(71637) <= 3692149;
srom_1(71638) <= 4178856;
srom_1(71639) <= 4685304;
srom_1(71640) <= 5209118;
srom_1(71641) <= 5747842;
srom_1(71642) <= 6298949;
srom_1(71643) <= 6859855;
srom_1(71644) <= 7427931;
srom_1(71645) <= 8000511;
srom_1(71646) <= 8574911;
srom_1(71647) <= 9148437;
srom_1(71648) <= 9718400;
srom_1(71649) <= 10282128;
srom_1(71650) <= 10836976;
srom_1(71651) <= 11380342;
srom_1(71652) <= 11909680;
srom_1(71653) <= 12422506;
srom_1(71654) <= 12916415;
srom_1(71655) <= 13389093;
srom_1(71656) <= 13838321;
srom_1(71657) <= 14261993;
srom_1(71658) <= 14658124;
srom_1(71659) <= 15024854;
srom_1(71660) <= 15360465;
srom_1(71661) <= 15663382;
srom_1(71662) <= 15932185;
srom_1(71663) <= 16165614;
srom_1(71664) <= 16362574;
srom_1(71665) <= 16522141;
srom_1(71666) <= 16643567;
srom_1(71667) <= 16726283;
srom_1(71668) <= 16769901;
srom_1(71669) <= 16774216;
srom_1(71670) <= 16739208;
srom_1(71671) <= 16665041;
srom_1(71672) <= 16552063;
srom_1(71673) <= 16400804;
srom_1(71674) <= 16211972;
srom_1(71675) <= 15986455;
srom_1(71676) <= 15725308;
srom_1(71677) <= 15429757;
srom_1(71678) <= 15101188;
srom_1(71679) <= 14741141;
srom_1(71680) <= 14351305;
srom_1(71681) <= 13933508;
srom_1(71682) <= 13489709;
srom_1(71683) <= 13021989;
srom_1(71684) <= 12532541;
srom_1(71685) <= 12023661;
srom_1(71686) <= 11497735;
srom_1(71687) <= 10957230;
srom_1(71688) <= 10404679;
srom_1(71689) <= 9842674;
srom_1(71690) <= 9273851;
srom_1(71691) <= 8700876;
srom_1(71692) <= 8126437;
srom_1(71693) <= 7553227;
srom_1(71694) <= 6983935;
srom_1(71695) <= 6421230;
srom_1(71696) <= 5867750;
srom_1(71697) <= 5326092;
srom_1(71698) <= 4798795;
srom_1(71699) <= 4288331;
srom_1(71700) <= 3797096;
srom_1(71701) <= 3327391;
srom_1(71702) <= 2881420;
srom_1(71703) <= 2461275;
srom_1(71704) <= 2068924;
srom_1(71705) <= 1706209;
srom_1(71706) <= 1374830;
srom_1(71707) <= 1076341;
srom_1(71708) <= 812141;
srom_1(71709) <= 583470;
srom_1(71710) <= 391400;
srom_1(71711) <= 236832;
srom_1(71712) <= 120490;
srom_1(71713) <= 42921;
srom_1(71714) <= 4487;
srom_1(71715) <= 5369;
srom_1(71716) <= 45563;
srom_1(71717) <= 124880;
srom_1(71718) <= 242949;
srom_1(71719) <= 399216;
srom_1(71720) <= 592948;
srom_1(71721) <= 823236;
srom_1(71722) <= 1089000;
srom_1(71723) <= 1388996;
srom_1(71724) <= 1721814;
srom_1(71725) <= 2085896;
srom_1(71726) <= 2479533;
srom_1(71727) <= 2900880;
srom_1(71728) <= 3347961;
srom_1(71729) <= 3818679;
srom_1(71730) <= 4310827;
srom_1(71731) <= 4822097;
srom_1(71732) <= 5350091;
srom_1(71733) <= 5892335;
srom_1(71734) <= 6446284;
srom_1(71735) <= 7009341;
srom_1(71736) <= 7578866;
srom_1(71737) <= 8152189;
srom_1(71738) <= 8726620;
srom_1(71739) <= 9299466;
srom_1(71740) <= 9868041;
srom_1(71741) <= 10429678;
srom_1(71742) <= 10981743;
srom_1(71743) <= 11521649;
srom_1(71744) <= 12046863;
srom_1(71745) <= 12554922;
srom_1(71746) <= 13043443;
srom_1(71747) <= 13510137;
srom_1(71748) <= 13952814;
srom_1(71749) <= 14369398;
srom_1(71750) <= 14757937;
srom_1(71751) <= 15116607;
srom_1(71752) <= 15443728;
srom_1(71753) <= 15737765;
srom_1(71754) <= 15997338;
srom_1(71755) <= 16221232;
srom_1(71756) <= 16408397;
srom_1(71757) <= 16557953;
srom_1(71758) <= 16669201;
srom_1(71759) <= 16741618;
srom_1(71760) <= 16774865;
srom_1(71761) <= 16768786;
srom_1(71762) <= 16723409;
srom_1(71763) <= 16638948;
srom_1(71764) <= 16515798;
srom_1(71765) <= 16354537;
srom_1(71766) <= 16155921;
srom_1(71767) <= 15920881;
srom_1(71768) <= 15650520;
srom_1(71769) <= 15346105;
srom_1(71770) <= 15009064;
srom_1(71771) <= 14640977;
srom_1(71772) <= 14243571;
srom_1(71773) <= 13818709;
srom_1(71774) <= 13368384;
srom_1(71775) <= 12894706;
srom_1(71776) <= 12399898;
srom_1(71777) <= 11886279;
srom_1(71778) <= 11356259;
srom_1(71779) <= 10812323;
srom_1(71780) <= 10257020;
srom_1(71781) <= 9692957;
srom_1(71782) <= 9122776;
srom_1(71783) <= 8549153;
srom_1(71784) <= 7974777;
srom_1(71785) <= 7402341;
srom_1(71786) <= 6834531;
srom_1(71787) <= 6274008;
srom_1(71788) <= 5723401;
srom_1(71789) <= 5185292;
srom_1(71790) <= 4662205;
srom_1(71791) <= 4156592;
srom_1(71792) <= 3670824;
srom_1(71793) <= 3207180;
srom_1(71794) <= 2767833;
srom_1(71795) <= 2354844;
srom_1(71796) <= 1970150;
srom_1(71797) <= 1615553;
srom_1(71798) <= 1292718;
srom_1(71799) <= 1003158;
srom_1(71800) <= 748231;
srom_1(71801) <= 529132;
srom_1(71802) <= 346889;
srom_1(71803) <= 202356;
srom_1(71804) <= 96212;
srom_1(71805) <= 28953;
srom_1(71806) <= 896;
srom_1(71807) <= 12171;
srom_1(71808) <= 62726;
srom_1(71809) <= 152325;
srom_1(71810) <= 280546;
srom_1(71811) <= 446789;
srom_1(71812) <= 650273;
srom_1(71813) <= 890045;
srom_1(71814) <= 1164981;
srom_1(71815) <= 1473790;
srom_1(71816) <= 1815026;
srom_1(71817) <= 2187087;
srom_1(71818) <= 2588230;
srom_1(71819) <= 3016572;
srom_1(71820) <= 3470106;
srom_1(71821) <= 3946704;
srom_1(71822) <= 4444132;
srom_1(71823) <= 4960057;
srom_1(71824) <= 5492059;
srom_1(71825) <= 6037644;
srom_1(71826) <= 6594254;
srom_1(71827) <= 7159278;
srom_1(71828) <= 7730067;
srom_1(71829) <= 8303944;
srom_1(71830) <= 8878218;
srom_1(71831) <= 9450197;
srom_1(71832) <= 10017196;
srom_1(71833) <= 10576559;
srom_1(71834) <= 11125662;
srom_1(71835) <= 11661930;
srom_1(71836) <= 12182848;
srom_1(71837) <= 12685974;
srom_1(71838) <= 13168948;
srom_1(71839) <= 13629505;
srom_1(71840) <= 14065485;
srom_1(71841) <= 14474845;
srom_1(71842) <= 14855665;
srom_1(71843) <= 15206158;
srom_1(71844) <= 15524681;
srom_1(71845) <= 15809741;
srom_1(71846) <= 16060001;
srom_1(71847) <= 16274286;
srom_1(71848) <= 16451594;
srom_1(71849) <= 16591091;
srom_1(71850) <= 16692123;
srom_1(71851) <= 16754218;
srom_1(71852) <= 16777083;
srom_1(71853) <= 16760612;
srom_1(71854) <= 16704882;
srom_1(71855) <= 16610154;
srom_1(71856) <= 16476872;
srom_1(71857) <= 16305662;
srom_1(71858) <= 16097326;
srom_1(71859) <= 15852841;
srom_1(71860) <= 15573353;
srom_1(71861) <= 15260174;
srom_1(71862) <= 14914772;
srom_1(71863) <= 14538766;
srom_1(71864) <= 14133920;
srom_1(71865) <= 13702133;
srom_1(71866) <= 13245428;
srom_1(71867) <= 12765948;
srom_1(71868) <= 12265942;
srom_1(71869) <= 11747753;
srom_1(71870) <= 11213811;
srom_1(71871) <= 10666622;
srom_1(71872) <= 10108750;
srom_1(71873) <= 9542812;
srom_1(71874) <= 8971461;
srom_1(71875) <= 8397377;
srom_1(71876) <= 7823252;
srom_1(71877) <= 7251778;
srom_1(71878) <= 6685635;
srom_1(71879) <= 6127478;
srom_1(71880) <= 5579925;
srom_1(71881) <= 5045542;
srom_1(71882) <= 4526835;
srom_1(71883) <= 4026238;
srom_1(71884) <= 3546098;
srom_1(71885) <= 3088666;
srom_1(71886) <= 2656087;
srom_1(71887) <= 2250389;
srom_1(71888) <= 1873476;
srom_1(71889) <= 1527115;
srom_1(71890) <= 1212930;
srom_1(71891) <= 932393;
srom_1(71892) <= 686822;
srom_1(71893) <= 477367;
srom_1(71894) <= 305010;
srom_1(71895) <= 170560;
srom_1(71896) <= 74648;
srom_1(71897) <= 17722;
srom_1(71898) <= 50;
srom_1(71899) <= 21715;
srom_1(71900) <= 82616;
srom_1(71901) <= 182466;
srom_1(71902) <= 320797;
srom_1(71903) <= 496961;
srom_1(71904) <= 710132;
srom_1(71905) <= 959310;
srom_1(71906) <= 1243326;
srom_1(71907) <= 1560849;
srom_1(71908) <= 1910390;
srom_1(71909) <= 2290309;
srom_1(71910) <= 2698826;
srom_1(71911) <= 3134023;
srom_1(71912) <= 3593861;
srom_1(71913) <= 4076184;
srom_1(71914) <= 4578728;
srom_1(71915) <= 5099139;
srom_1(71916) <= 5634975;
srom_1(71917) <= 6183724;
srom_1(71918) <= 6742812;
srom_1(71919) <= 7309618;
srom_1(71920) <= 7881484;
srom_1(71921) <= 8455728;
srom_1(71922) <= 9029657;
srom_1(71923) <= 9600580;
srom_1(71924) <= 10165819;
srom_1(71925) <= 10722725;
srom_1(71926) <= 11268685;
srom_1(71927) <= 11801139;
srom_1(71928) <= 12317591;
srom_1(71929) <= 12815619;
srom_1(71930) <= 13292886;
srom_1(71931) <= 13747156;
srom_1(71932) <= 14176298;
srom_1(71933) <= 14578300;
srom_1(71934) <= 14951275;
srom_1(71935) <= 15293476;
srom_1(71936) <= 15603298;
srom_1(71937) <= 15879288;
srom_1(71938) <= 16120151;
srom_1(71939) <= 16324759;
srom_1(71940) <= 16492151;
srom_1(71941) <= 16621542;
srom_1(71942) <= 16712327;
srom_1(71943) <= 16764079;
srom_1(71944) <= 16776556;
srom_1(71945) <= 16749698;
srom_1(71946) <= 16683632;
srom_1(71947) <= 16578669;
srom_1(71948) <= 16435299;
srom_1(71949) <= 16254195;
srom_1(71950) <= 16036207;
srom_1(71951) <= 15782357;
srom_1(71952) <= 15493835;
srom_1(71953) <= 15171994;
srom_1(71954) <= 14818344;
srom_1(71955) <= 14434542;
srom_1(71956) <= 14022389;
srom_1(71957) <= 13583817;
srom_1(71958) <= 13120883;
srom_1(71959) <= 12635757;
srom_1(71960) <= 12130716;
srom_1(71961) <= 11608126;
srom_1(71962) <= 11070439;
srom_1(71963) <= 10520176;
srom_1(71964) <= 9959917;
srom_1(71965) <= 9392289;
srom_1(71966) <= 8819955;
srom_1(71967) <= 8245599;
srom_1(71968) <= 7671913;
srom_1(71969) <= 7101588;
srom_1(71970) <= 6537298;
srom_1(71971) <= 5981689;
srom_1(71972) <= 5437367;
srom_1(71973) <= 4906885;
srom_1(71974) <= 4392730;
srom_1(71975) <= 3897313;
srom_1(71976) <= 3422957;
srom_1(71977) <= 2971886;
srom_1(71978) <= 2546217;
srom_1(71979) <= 2147944;
srom_1(71980) <= 1778936;
srom_1(71981) <= 1440923;
srom_1(71982) <= 1135490;
srom_1(71983) <= 864070;
srom_1(71984) <= 627935;
srom_1(71985) <= 428192;
srom_1(71986) <= 265778;
srom_1(71987) <= 141455;
srom_1(71988) <= 55805;
srom_1(71989) <= 9231;
srom_1(71990) <= 1951;
srom_1(71991) <= 33999;
srom_1(71992) <= 105224;
srom_1(71993) <= 215293;
srom_1(71994) <= 363690;
srom_1(71995) <= 549718;
srom_1(71996) <= 772505;
srom_1(71997) <= 1031007;
srom_1(71998) <= 1324011;
srom_1(71999) <= 1650143;
srom_1(72000) <= 2007875;
srom_1(72001) <= 2395528;
srom_1(72002) <= 2811284;
srom_1(72003) <= 3253194;
srom_1(72004) <= 3719187;
srom_1(72005) <= 4207075;
srom_1(72006) <= 4714572;
srom_1(72007) <= 5239299;
srom_1(72008) <= 5778793;
srom_1(72009) <= 6330525;
srom_1(72010) <= 6891909;
srom_1(72011) <= 7460311;
srom_1(72012) <= 8033066;
srom_1(72013) <= 8607489;
srom_1(72014) <= 9180885;
srom_1(72015) <= 9750566;
srom_1(72016) <= 10313860;
srom_1(72017) <= 10868126;
srom_1(72018) <= 11410765;
srom_1(72019) <= 11939231;
srom_1(72020) <= 12451048;
srom_1(72021) <= 12943814;
srom_1(72022) <= 13415220;
srom_1(72023) <= 13863054;
srom_1(72024) <= 14285216;
srom_1(72025) <= 14679727;
srom_1(72026) <= 15044737;
srom_1(72027) <= 15378534;
srom_1(72028) <= 15679553;
srom_1(72029) <= 15946382;
srom_1(72030) <= 16177771;
srom_1(72031) <= 16372633;
srom_1(72032) <= 16530055;
srom_1(72033) <= 16649299;
srom_1(72034) <= 16729806;
srom_1(72035) <= 16771198;
srom_1(72036) <= 16773281;
srom_1(72037) <= 16736046;
srom_1(72038) <= 16659667;
srom_1(72039) <= 16544502;
srom_1(72040) <= 16391091;
srom_1(72041) <= 16200153;
srom_1(72042) <= 15972585;
srom_1(72043) <= 15709453;
srom_1(72044) <= 15411991;
srom_1(72045) <= 15081593;
srom_1(72046) <= 14719810;
srom_1(72047) <= 14328338;
srom_1(72048) <= 13909013;
srom_1(72049) <= 13463800;
srom_1(72050) <= 12994788;
srom_1(72051) <= 12504176;
srom_1(72052) <= 11994265;
srom_1(72053) <= 11467445;
srom_1(72054) <= 10926188;
srom_1(72055) <= 10373031;
srom_1(72056) <= 9810569;
srom_1(72057) <= 9241438;
srom_1(72058) <= 8668308;
srom_1(72059) <= 8093867;
srom_1(72060) <= 7520808;
srom_1(72061) <= 6951818;
srom_1(72062) <= 6389566;
srom_1(72063) <= 5836688;
srom_1(72064) <= 5295777;
srom_1(72065) <= 4769369;
srom_1(72066) <= 4259933;
srom_1(72067) <= 3769857;
srom_1(72068) <= 3301441;
srom_1(72069) <= 2856880;
srom_1(72070) <= 2438260;
srom_1(72071) <= 2047542;
srom_1(72072) <= 1686560;
srom_1(72073) <= 1357006;
srom_1(72074) <= 1060426;
srom_1(72075) <= 798210;
srom_1(72076) <= 571588;
srom_1(72077) <= 381623;
srom_1(72078) <= 229205;
srom_1(72079) <= 115049;
srom_1(72080) <= 39691;
srom_1(72081) <= 3484;
srom_1(72082) <= 6598;
srom_1(72083) <= 49018;
srom_1(72084) <= 130545;
srom_1(72085) <= 250797;
srom_1(72086) <= 409210;
srom_1(72087) <= 605041;
srom_1(72088) <= 837371;
srom_1(72089) <= 1105113;
srom_1(72090) <= 1407009;
srom_1(72091) <= 1741644;
srom_1(72092) <= 2107449;
srom_1(72093) <= 2502708;
srom_1(72094) <= 2925568;
srom_1(72095) <= 3374047;
srom_1(72096) <= 3846041;
srom_1(72097) <= 4339336;
srom_1(72098) <= 4851619;
srom_1(72099) <= 5380489;
srom_1(72100) <= 5923465;
srom_1(72101) <= 6478001;
srom_1(72102) <= 7041496;
srom_1(72103) <= 7611308;
srom_1(72104) <= 8184765;
srom_1(72105) <= 8759179;
srom_1(72106) <= 9331854;
srom_1(72107) <= 9900106;
srom_1(72108) <= 10461271;
srom_1(72109) <= 11012715;
srom_1(72110) <= 11551855;
srom_1(72111) <= 12076161;
srom_1(72112) <= 12583175;
srom_1(72113) <= 13070519;
srom_1(72114) <= 13535908;
srom_1(72115) <= 13977159;
srom_1(72116) <= 14392204;
srom_1(72117) <= 14779096;
srom_1(72118) <= 15136020;
srom_1(72119) <= 15461304;
srom_1(72120) <= 15753421;
srom_1(72121) <= 16011003;
srom_1(72122) <= 16232840;
srom_1(72123) <= 16417893;
srom_1(72124) <= 16565293;
srom_1(72125) <= 16674351;
srom_1(72126) <= 16744554;
srom_1(72127) <= 16775573;
srom_1(72128) <= 16767262;
srom_1(72129) <= 16719661;
srom_1(72130) <= 16632993;
srom_1(72131) <= 16507665;
srom_1(72132) <= 16344263;
srom_1(72133) <= 16143554;
srom_1(72134) <= 15906480;
srom_1(72135) <= 15634152;
srom_1(72136) <= 15327847;
srom_1(72137) <= 14989001;
srom_1(72138) <= 14619204;
srom_1(72139) <= 14220190;
srom_1(72140) <= 13793829;
srom_1(72141) <= 13342122;
srom_1(72142) <= 12867185;
srom_1(72143) <= 12371247;
srom_1(72144) <= 11856633;
srom_1(72145) <= 11325756;
srom_1(72146) <= 10781106;
srom_1(72147) <= 10225237;
srom_1(72148) <= 9660755;
srom_1(72149) <= 9090308;
srom_1(72150) <= 8516570;
srom_1(72151) <= 7942232;
srom_1(72152) <= 7369987;
srom_1(72153) <= 6802519;
srom_1(72154) <= 6242489;
srom_1(72155) <= 5692522;
srom_1(72156) <= 5155198;
srom_1(72157) <= 4633037;
srom_1(72158) <= 4128487;
srom_1(72159) <= 3643914;
srom_1(72160) <= 3181591;
srom_1(72161) <= 2743685;
srom_1(72162) <= 2332250;
srom_1(72163) <= 1949216;
srom_1(72164) <= 1596378;
srom_1(72165) <= 1275391;
srom_1(72166) <= 987760;
srom_1(72167) <= 734835;
srom_1(72168) <= 517801;
srom_1(72169) <= 337675;
srom_1(72170) <= 195303;
srom_1(72171) <= 91353;
srom_1(72172) <= 26311;
srom_1(72173) <= 483;
srom_1(72174) <= 13989;
srom_1(72175) <= 66767;
srom_1(72176) <= 158569;
srom_1(72177) <= 288964;
srom_1(72178) <= 457342;
srom_1(72179) <= 662912;
srom_1(72180) <= 904710;
srom_1(72181) <= 1181603;
srom_1(72182) <= 1492292;
srom_1(72183) <= 1835320;
srom_1(72184) <= 2209079;
srom_1(72185) <= 2611815;
srom_1(72186) <= 3041642;
srom_1(72187) <= 3496541;
srom_1(72188) <= 3974382;
srom_1(72189) <= 4472922;
srom_1(72190) <= 4989824;
srom_1(72191) <= 5522664;
srom_1(72192) <= 6068944;
srom_1(72193) <= 6626101;
srom_1(72194) <= 7191524;
srom_1(72195) <= 7762560;
srom_1(72196) <= 8336531;
srom_1(72197) <= 8910747;
srom_1(72198) <= 9482514;
srom_1(72199) <= 10049152;
srom_1(72200) <= 10608003;
srom_1(72201) <= 11156446;
srom_1(72202) <= 11691910;
srom_1(72203) <= 12211883;
srom_1(72204) <= 12713928;
srom_1(72205) <= 13195690;
srom_1(72206) <= 13654910;
srom_1(72207) <= 14089434;
srom_1(72208) <= 14497226;
srom_1(72209) <= 14876372;
srom_1(72210) <= 15225094;
srom_1(72211) <= 15541758;
srom_1(72212) <= 15824878;
srom_1(72213) <= 16073127;
srom_1(72214) <= 16285341;
srom_1(72215) <= 16460524;
srom_1(72216) <= 16597855;
srom_1(72217) <= 16696690;
srom_1(72218) <= 16756566;
srom_1(72219) <= 16777202;
srom_1(72220) <= 16758500;
srom_1(72221) <= 16700549;
srom_1(72222) <= 16603621;
srom_1(72223) <= 16468170;
srom_1(72224) <= 16294830;
srom_1(72225) <= 16084416;
srom_1(72226) <= 15837913;
srom_1(72227) <= 15556479;
srom_1(72228) <= 15241431;
srom_1(72229) <= 14894248;
srom_1(72230) <= 14516558;
srom_1(72231) <= 14110132;
srom_1(72232) <= 13676876;
srom_1(72233) <= 13218821;
srom_1(72234) <= 12738116;
srom_1(72235) <= 12237014;
srom_1(72236) <= 11717866;
srom_1(72237) <= 11183106;
srom_1(72238) <= 10635242;
srom_1(72239) <= 10076842;
srom_1(72240) <= 9510525;
srom_1(72241) <= 8938948;
srom_1(72242) <= 8364790;
srom_1(72243) <= 7790743;
srom_1(72244) <= 7219500;
srom_1(72245) <= 6653739;
srom_1(72246) <= 6096114;
srom_1(72247) <= 5549239;
srom_1(72248) <= 5015679;
srom_1(72249) <= 4497935;
srom_1(72250) <= 3998436;
srom_1(72251) <= 3519525;
srom_1(72252) <= 3063446;
srom_1(72253) <= 2632338;
srom_1(72254) <= 2228224;
srom_1(72255) <= 1852998;
srom_1(72256) <= 1508420;
srom_1(72257) <= 1196105;
srom_1(72258) <= 917518;
srom_1(72259) <= 673966;
srom_1(72260) <= 466590;
srom_1(72261) <= 296363;
srom_1(72262) <= 164084;
srom_1(72263) <= 70373;
srom_1(72264) <= 15668;
srom_1(72265) <= 227;
srom_1(72266) <= 24122;
srom_1(72267) <= 87241;
srom_1(72268) <= 189288;
srom_1(72269) <= 329784;
srom_1(72270) <= 508071;
srom_1(72271) <= 723312;
srom_1(72272) <= 974499;
srom_1(72273) <= 1260453;
srom_1(72274) <= 1579833;
srom_1(72275) <= 1931142;
srom_1(72276) <= 2312732;
srom_1(72277) <= 2722814;
srom_1(72278) <= 3159465;
srom_1(72279) <= 3620637;
srom_1(72280) <= 4104168;
srom_1(72281) <= 4607790;
srom_1(72282) <= 5129142;
srom_1(72283) <= 5665778;
srom_1(72284) <= 6215183;
srom_1(72285) <= 6774779;
srom_1(72286) <= 7341943;
srom_1(72287) <= 7914016;
srom_1(72288) <= 8488314;
srom_1(72289) <= 9062144;
srom_1(72290) <= 9632816;
srom_1(72291) <= 10197654;
srom_1(72292) <= 10754008;
srom_1(72293) <= 11299270;
srom_1(72294) <= 11830883;
srom_1(72295) <= 12346354;
srom_1(72296) <= 12843266;
srom_1(72297) <= 13319288;
srom_1(72298) <= 13772188;
srom_1(72299) <= 14199844;
srom_1(72300) <= 14600248;
srom_1(72301) <= 14971523;
srom_1(72302) <= 15311930;
srom_1(72303) <= 15619870;
srom_1(72304) <= 15893900;
srom_1(72305) <= 16132736;
srom_1(72306) <= 16335257;
srom_1(72307) <= 16500513;
srom_1(72308) <= 16627729;
srom_1(72309) <= 16716310;
srom_1(72310) <= 16765839;
srom_1(72311) <= 16776084;
srom_1(72312) <= 16746998;
srom_1(72313) <= 16678716;
srom_1(72314) <= 16571559;
srom_1(72315) <= 16426029;
srom_1(72316) <= 16242809;
srom_1(72317) <= 16022758;
srom_1(72318) <= 15766908;
srom_1(72319) <= 15476459;
srom_1(72320) <= 15152772;
srom_1(72321) <= 14797365;
srom_1(72322) <= 14411906;
srom_1(72323) <= 13998202;
srom_1(72324) <= 13558192;
srom_1(72325) <= 13093940;
srom_1(72326) <= 12607623;
srom_1(72327) <= 12101522;
srom_1(72328) <= 11578010;
srom_1(72329) <= 11039541;
srom_1(72330) <= 10488641;
srom_1(72331) <= 9927894;
srom_1(72332) <= 9359928;
srom_1(72333) <= 8787408;
srom_1(72334) <= 8213017;
srom_1(72335) <= 7639450;
srom_1(72336) <= 7069395;
srom_1(72337) <= 6505527;
srom_1(72338) <= 5950490;
srom_1(72339) <= 5406885;
srom_1(72340) <= 4877263;
srom_1(72341) <= 4364107;
srom_1(72342) <= 3869823;
srom_1(72343) <= 3396729;
srom_1(72344) <= 2947044;
srom_1(72345) <= 2522876;
srom_1(72346) <= 2126215;
srom_1(72347) <= 1758920;
srom_1(72348) <= 1422714;
srom_1(72349) <= 1119173;
srom_1(72350) <= 849722;
srom_1(72351) <= 615622;
srom_1(72352) <= 417973;
srom_1(72353) <= 257701;
srom_1(72354) <= 135558;
srom_1(72355) <= 52116;
srom_1(72356) <= 7766;
srom_1(72357) <= 2718;
srom_1(72358) <= 36993;
srom_1(72359) <= 110432;
srom_1(72360) <= 222691;
srom_1(72361) <= 373242;
srom_1(72362) <= 561380;
srom_1(72363) <= 786222;
srom_1(72364) <= 1046715;
srom_1(72365) <= 1341636;
srom_1(72366) <= 1669603;
srom_1(72367) <= 2029078;
srom_1(72368) <= 2418375;
srom_1(72369) <= 2835668;
srom_1(72370) <= 3279001;
srom_1(72371) <= 3746294;
srom_1(72372) <= 4235357;
srom_1(72373) <= 4743896;
srom_1(72374) <= 5269526;
srom_1(72375) <= 5809783;
srom_1(72376) <= 6362133;
srom_1(72377) <= 6923985;
srom_1(72378) <= 7492706;
srom_1(72379) <= 8065628;
srom_1(72380) <= 8640064;
srom_1(72381) <= 9213321;
srom_1(72382) <= 9782711;
srom_1(72383) <= 10345563;
srom_1(72384) <= 10899239;
srom_1(72385) <= 11441141;
srom_1(72386) <= 11968729;
srom_1(72387) <= 12479529;
srom_1(72388) <= 12971145;
srom_1(72389) <= 13441271;
srom_1(72390) <= 13887704;
srom_1(72391) <= 14308350;
srom_1(72392) <= 14701236;
srom_1(72393) <= 15064520;
srom_1(72394) <= 15396499;
srom_1(72395) <= 15695615;
srom_1(72396) <= 15960465;
srom_1(72397) <= 16189809;
srom_1(72398) <= 16382571;
srom_1(72399) <= 16537846;
srom_1(72400) <= 16654906;
srom_1(72401) <= 16733203;
srom_1(72402) <= 16772369;
srom_1(72403) <= 16772221;
srom_1(72404) <= 16732759;
srom_1(72405) <= 16654168;
srom_1(72406) <= 16536818;
srom_1(72407) <= 16381257;
srom_1(72408) <= 16188217;
srom_1(72409) <= 15958601;
srom_1(72410) <= 15693487;
srom_1(72411) <= 15394118;
srom_1(72412) <= 15061898;
srom_1(72413) <= 14698384;
srom_1(72414) <= 14305282;
srom_1(72415) <= 13884434;
srom_1(72416) <= 13437815;
srom_1(72417) <= 12967518;
srom_1(72418) <= 12475749;
srom_1(72419) <= 11964814;
srom_1(72420) <= 11437108;
srom_1(72421) <= 10895108;
srom_1(72422) <= 10341353;
srom_1(72423) <= 9778442;
srom_1(72424) <= 9209013;
srom_1(72425) <= 8635737;
srom_1(72426) <= 8061302;
srom_1(72427) <= 7488402;
srom_1(72428) <= 6919723;
srom_1(72429) <= 6357932;
srom_1(72430) <= 5805664;
srom_1(72431) <= 5265508;
srom_1(72432) <= 4739997;
srom_1(72433) <= 4231596;
srom_1(72434) <= 3742689;
srom_1(72435) <= 3275568;
srom_1(72436) <= 2832424;
srom_1(72437) <= 2415334;
srom_1(72438) <= 2026256;
srom_1(72439) <= 1667012;
srom_1(72440) <= 1339289;
srom_1(72441) <= 1044622;
srom_1(72442) <= 784393;
srom_1(72443) <= 559824;
srom_1(72444) <= 371966;
srom_1(72445) <= 221701;
srom_1(72446) <= 109733;
srom_1(72447) <= 36588;
srom_1(72448) <= 2608;
srom_1(72449) <= 7954;
srom_1(72450) <= 52599;
srom_1(72451) <= 136334;
srom_1(72452) <= 258767;
srom_1(72453) <= 419324;
srom_1(72454) <= 617251;
srom_1(72455) <= 851621;
srom_1(72456) <= 1121335;
srom_1(72457) <= 1425127;
srom_1(72458) <= 1761573;
srom_1(72459) <= 2129096;
srom_1(72460) <= 2525972;
srom_1(72461) <= 2950339;
srom_1(72462) <= 3400209;
srom_1(72463) <= 3873471;
srom_1(72464) <= 4367906;
srom_1(72465) <= 4881195;
srom_1(72466) <= 5410932;
srom_1(72467) <= 5954632;
srom_1(72468) <= 6509746;
srom_1(72469) <= 7073671;
srom_1(72470) <= 7643762;
srom_1(72471) <= 8217345;
srom_1(72472) <= 8791732;
srom_1(72473) <= 9364228;
srom_1(72474) <= 9932149;
srom_1(72475) <= 10492832;
srom_1(72476) <= 11043648;
srom_1(72477) <= 11582013;
srom_1(72478) <= 12105403;
srom_1(72479) <= 12611364;
srom_1(72480) <= 13097523;
srom_1(72481) <= 13561600;
srom_1(72482) <= 14001420;
srom_1(72483) <= 14414918;
srom_1(72484) <= 14800158;
srom_1(72485) <= 15155331;
srom_1(72486) <= 15478773;
srom_1(72487) <= 15768967;
srom_1(72488) <= 16024552;
srom_1(72489) <= 16244329;
srom_1(72490) <= 16427268;
srom_1(72491) <= 16572510;
srom_1(72492) <= 16679376;
srom_1(72493) <= 16747364;
srom_1(72494) <= 16776154;
srom_1(72495) <= 16765612;
srom_1(72496) <= 16715788;
srom_1(72497) <= 16626915;
srom_1(72498) <= 16499409;
srom_1(72499) <= 16333869;
srom_1(72500) <= 16131071;
srom_1(72501) <= 15891966;
srom_1(72502) <= 15617675;
srom_1(72503) <= 15309484;
srom_1(72504) <= 14968839;
srom_1(72505) <= 14597337;
srom_1(72506) <= 14196721;
srom_1(72507) <= 13768868;
srom_1(72508) <= 13315785;
srom_1(72509) <= 12839597;
srom_1(72510) <= 12342536;
srom_1(72511) <= 11826935;
srom_1(72512) <= 11295209;
srom_1(72513) <= 10749854;
srom_1(72514) <= 10193426;
srom_1(72515) <= 9628535;
srom_1(72516) <= 9057829;
srom_1(72517) <= 8483985;
srom_1(72518) <= 7909694;
srom_1(72519) <= 7337648;
srom_1(72520) <= 6770531;
srom_1(72521) <= 6211002;
srom_1(72522) <= 5661684;
srom_1(72523) <= 5125153;
srom_1(72524) <= 4603926;
srom_1(72525) <= 4100447;
srom_1(72526) <= 3617076;
srom_1(72527) <= 3156081;
srom_1(72528) <= 2719622;
srom_1(72529) <= 2309748;
srom_1(72530) <= 1928379;
srom_1(72531) <= 1577305;
srom_1(72532) <= 1258171;
srom_1(72533) <= 972475;
srom_1(72534) <= 721555;
srom_1(72535) <= 506588;
srom_1(72536) <= 328583;
srom_1(72537) <= 188374;
srom_1(72538) <= 86619;
srom_1(72539) <= 23795;
srom_1(72540) <= 196;
srom_1(72541) <= 15933;
srom_1(72542) <= 70933;
srom_1(72543) <= 164937;
srom_1(72544) <= 297505;
srom_1(72545) <= 468015;
srom_1(72546) <= 675667;
srom_1(72547) <= 919488;
srom_1(72548) <= 1198334;
srom_1(72549) <= 1510897;
srom_1(72550) <= 1855713;
srom_1(72551) <= 2231163;
srom_1(72552) <= 2635488;
srom_1(72553) <= 3066792;
srom_1(72554) <= 3523051;
srom_1(72555) <= 4002126;
srom_1(72556) <= 4501771;
srom_1(72557) <= 5019643;
srom_1(72558) <= 5553313;
srom_1(72559) <= 6100279;
srom_1(72560) <= 6657975;
srom_1(72561) <= 7223787;
srom_1(72562) <= 7795061;
srom_1(72563) <= 8369119;
srom_1(72564) <= 8943268;
srom_1(72565) <= 9514815;
srom_1(72566) <= 10081082;
srom_1(72567) <= 10639412;
srom_1(72568) <= 11187188;
srom_1(72569) <= 11721840;
srom_1(72570) <= 12240861;
srom_1(72571) <= 12741817;
srom_1(72572) <= 13222360;
srom_1(72573) <= 13680236;
srom_1(72574) <= 14113297;
srom_1(72575) <= 14519514;
srom_1(72576) <= 14896980;
srom_1(72577) <= 15243927;
srom_1(72578) <= 15558727;
srom_1(72579) <= 15839903;
srom_1(72580) <= 16086138;
srom_1(72581) <= 16296276;
srom_1(72582) <= 16469333;
srom_1(72583) <= 16604496;
srom_1(72584) <= 16701132;
srom_1(72585) <= 16758788;
srom_1(72586) <= 16777193;
srom_1(72587) <= 16756261;
srom_1(72588) <= 16696091;
srom_1(72589) <= 16596964;
srom_1(72590) <= 16459345;
srom_1(72591) <= 16283879;
srom_1(72592) <= 16071390;
srom_1(72593) <= 15822874;
srom_1(72594) <= 15539496;
srom_1(72595) <= 15222584;
srom_1(72596) <= 14873626;
srom_1(72597) <= 14494258;
srom_1(72598) <= 14086258;
srom_1(72599) <= 13651540;
srom_1(72600) <= 13192142;
srom_1(72601) <= 12710218;
srom_1(72602) <= 12208029;
srom_1(72603) <= 11687930;
srom_1(72604) <= 11152359;
srom_1(72605) <= 10603827;
srom_1(72606) <= 10044908;
srom_1(72607) <= 9478222;
srom_1(72608) <= 8906426;
srom_1(72609) <= 8332202;
srom_1(72610) <= 7758243;
srom_1(72611) <= 7187239;
srom_1(72612) <= 6621869;
srom_1(72613) <= 6064784;
srom_1(72614) <= 5518596;
srom_1(72615) <= 4985867;
srom_1(72616) <= 4469094;
srom_1(72617) <= 3970701;
srom_1(72618) <= 3493025;
srom_1(72619) <= 3038306;
srom_1(72620) <= 2608677;
srom_1(72621) <= 2206152;
srom_1(72622) <= 1832618;
srom_1(72623) <= 1489828;
srom_1(72624) <= 1179388;
srom_1(72625) <= 902755;
srom_1(72626) <= 661226;
srom_1(72627) <= 455933;
srom_1(72628) <= 287839;
srom_1(72629) <= 157732;
srom_1(72630) <= 66223;
srom_1(72631) <= 13740;
srom_1(72632) <= 530;
srom_1(72633) <= 26655;
srom_1(72634) <= 91991;
srom_1(72635) <= 196233;
srom_1(72636) <= 338892;
srom_1(72637) <= 519299;
srom_1(72638) <= 736608;
srom_1(72639) <= 989799;
srom_1(72640) <= 1277687;
srom_1(72641) <= 1598919;
srom_1(72642) <= 1951991;
srom_1(72643) <= 2335247;
srom_1(72644) <= 2746888;
srom_1(72645) <= 3184986;
srom_1(72646) <= 3647485;
srom_1(72647) <= 4132217;
srom_1(72648) <= 4636909;
srom_1(72649) <= 5159193;
srom_1(72650) <= 5696622;
srom_1(72651) <= 6246674;
srom_1(72652) <= 6806770;
srom_1(72653) <= 7374284;
srom_1(72654) <= 7946555;
srom_1(72655) <= 8520899;
srom_1(72656) <= 9094622;
srom_1(72657) <= 9665034;
srom_1(72658) <= 10229461;
srom_1(72659) <= 10785255;
srom_1(72660) <= 11329811;
srom_1(72661) <= 11860575;
srom_1(72662) <= 12375057;
srom_1(72663) <= 12870845;
srom_1(72664) <= 13345615;
srom_1(72665) <= 13797139;
srom_1(72666) <= 14223301;
srom_1(72667) <= 14622102;
srom_1(72668) <= 14991672;
srom_1(72669) <= 15330278;
srom_1(72670) <= 15636332;
srom_1(72671) <= 15908400;
srom_1(72672) <= 16145204;
srom_1(72673) <= 16345635;
srom_1(72674) <= 16508752;
srom_1(72675) <= 16633792;
srom_1(72676) <= 16720167;
srom_1(72677) <= 16767472;
srom_1(72678) <= 16775486;
srom_1(72679) <= 16744171;
srom_1(72680) <= 16673674;
srom_1(72681) <= 16564325;
srom_1(72682) <= 16416638;
srom_1(72683) <= 16231305;
srom_1(72684) <= 16009194;
srom_1(72685) <= 15751348;
srom_1(72686) <= 15458975;
srom_1(72687) <= 15133447;
srom_1(72688) <= 14776290;
srom_1(72689) <= 14389179;
srom_1(72690) <= 13973930;
srom_1(72691) <= 13532488;
srom_1(72692) <= 13066926;
srom_1(72693) <= 12579425;
srom_1(72694) <= 12072272;
srom_1(72695) <= 11547845;
srom_1(72696) <= 11008603;
srom_1(72697) <= 10457075;
srom_1(72698) <= 9895848;
srom_1(72699) <= 9327552;
srom_1(72700) <= 8754854;
srom_1(72701) <= 8180438;
srom_1(72702) <= 7606998;
srom_1(72703) <= 7037223;
srom_1(72704) <= 6473785;
srom_1(72705) <= 5919327;
srom_1(72706) <= 5376448;
srom_1(72707) <= 4847694;
srom_1(72708) <= 4335545;
srom_1(72709) <= 3842402;
srom_1(72710) <= 3370577;
srom_1(72711) <= 2922284;
srom_1(72712) <= 2499624;
srom_1(72713) <= 2104580;
srom_1(72714) <= 1739004;
srom_1(72715) <= 1404610;
srom_1(72716) <= 1102966;
srom_1(72717) <= 835487;
srom_1(72718) <= 603427;
srom_1(72719) <= 407875;
srom_1(72720) <= 249747;
srom_1(72721) <= 129785;
srom_1(72722) <= 48552;
srom_1(72723) <= 6428;
srom_1(72724) <= 3610;
srom_1(72725) <= 40113;
srom_1(72726) <= 115765;
srom_1(72727) <= 230211;
srom_1(72728) <= 382915;
srom_1(72729) <= 573160;
srom_1(72730) <= 800054;
srom_1(72731) <= 1062534;
srom_1(72732) <= 1359368;
srom_1(72733) <= 1689164;
srom_1(72734) <= 2050377;
srom_1(72735) <= 2441312;
srom_1(72736) <= 2860135;
srom_1(72737) <= 3304884;
srom_1(72738) <= 3773472;
srom_1(72739) <= 4263702;
srom_1(72740) <= 4773275;
srom_1(72741) <= 5299801;
srom_1(72742) <= 5840812;
srom_1(72743) <= 6393771;
srom_1(72744) <= 6956083;
srom_1(72745) <= 7525114;
srom_1(72746) <= 8098194;
srom_1(72747) <= 8672635;
srom_1(72748) <= 9245745;
srom_1(72749) <= 9814835;
srom_1(72750) <= 10377237;
srom_1(72751) <= 10930314;
srom_1(72752) <= 11471472;
srom_1(72753) <= 11998173;
srom_1(72754) <= 12507948;
srom_1(72755) <= 12998405;
srom_1(72756) <= 13467246;
srom_1(72757) <= 13912272;
srom_1(72758) <= 14331394;
srom_1(72759) <= 14722650;
srom_1(72760) <= 15084202;
srom_1(72761) <= 15414357;
srom_1(72762) <= 15711566;
srom_1(72763) <= 15974434;
srom_1(72764) <= 16201730;
srom_1(72765) <= 16392388;
srom_1(72766) <= 16545513;
srom_1(72767) <= 16660388;
srom_1(72768) <= 16736473;
srom_1(72769) <= 16773413;
srom_1(72770) <= 16771033;
srom_1(72771) <= 16729345;
srom_1(72772) <= 16648545;
srom_1(72773) <= 16529011;
srom_1(72774) <= 16371303;
srom_1(72775) <= 16176162;
srom_1(72776) <= 15944503;
srom_1(72777) <= 15677411;
srom_1(72778) <= 15376140;
srom_1(72779) <= 15042102;
srom_1(72780) <= 14676863;
srom_1(72781) <= 14282136;
srom_1(72782) <= 13859773;
srom_1(72783) <= 13411753;
srom_1(72784) <= 12940178;
srom_1(72785) <= 12447260;
srom_1(72786) <= 11935309;
srom_1(72787) <= 11406726;
srom_1(72788) <= 10863990;
srom_1(72789) <= 10309646;
srom_1(72790) <= 9746294;
srom_1(72791) <= 9176575;
srom_1(72792) <= 8603161;
srom_1(72793) <= 8028741;
srom_1(72794) <= 7456009;
srom_1(72795) <= 6887650;
srom_1(72796) <= 6326329;
srom_1(72797) <= 5774679;
srom_1(72798) <= 5235286;
srom_1(72799) <= 4710681;
srom_1(72800) <= 4203323;
srom_1(72801) <= 3715591;
srom_1(72802) <= 3249772;
srom_1(72803) <= 2808051;
srom_1(72804) <= 2392499;
srom_1(72805) <= 2005065;
srom_1(72806) <= 1647566;
srom_1(72807) <= 1321678;
srom_1(72808) <= 1028928;
srom_1(72809) <= 770691;
srom_1(72810) <= 548177;
srom_1(72811) <= 362430;
srom_1(72812) <= 214320;
srom_1(72813) <= 104542;
srom_1(72814) <= 33611;
srom_1(72815) <= 1859;
srom_1(72816) <= 9436;
srom_1(72817) <= 56305;
srom_1(72818) <= 142248;
srom_1(72819) <= 266860;
srom_1(72820) <= 429558;
srom_1(72821) <= 629579;
srom_1(72822) <= 865985;
srom_1(72823) <= 1137666;
srom_1(72824) <= 1443350;
srom_1(72825) <= 1781603;
srom_1(72826) <= 2150838;
srom_1(72827) <= 2549324;
srom_1(72828) <= 2975193;
srom_1(72829) <= 3426446;
srom_1(72830) <= 3900970;
srom_1(72831) <= 4396537;
srom_1(72832) <= 4910824;
srom_1(72833) <= 5441420;
srom_1(72834) <= 5985837;
srom_1(72835) <= 6541520;
srom_1(72836) <= 7105866;
srom_1(72837) <= 7676226;
srom_1(72838) <= 8249927;
srom_1(72839) <= 8824279;
srom_1(72840) <= 9396587;
srom_1(72841) <= 9964169;
srom_1(72842) <= 10524362;
srom_1(72843) <= 11074540;
srom_1(72844) <= 11612123;
srom_1(72845) <= 12134590;
srom_1(72846) <= 12639490;
srom_1(72847) <= 13124457;
srom_1(72848) <= 13587215;
srom_1(72849) <= 14025596;
srom_1(72850) <= 14437542;
srom_1(72851) <= 14821123;
srom_1(72852) <= 15174540;
srom_1(72853) <= 15496136;
srom_1(72854) <= 15784401;
srom_1(72855) <= 16037985;
srom_1(72856) <= 16255699;
srom_1(72857) <= 16436521;
srom_1(72858) <= 16579604;
srom_1(72859) <= 16684276;
srom_1(72860) <= 16750047;
srom_1(72861) <= 16776609;
srom_1(72862) <= 16763836;
srom_1(72863) <= 16711789;
srom_1(72864) <= 16620711;
srom_1(72865) <= 16491031;
srom_1(72866) <= 16323355;
srom_1(72867) <= 16118471;
srom_1(72868) <= 15877338;
srom_1(72869) <= 15601089;
srom_1(72870) <= 15291017;
srom_1(72871) <= 14948578;
srom_1(72872) <= 14575377;
srom_1(72873) <= 14173164;
srom_1(72874) <= 13743825;
srom_1(72875) <= 13289374;
srom_1(72876) <= 12811941;
srom_1(72877) <= 12313766;
srom_1(72878) <= 11797184;
srom_1(72879) <= 11264618;
srom_1(72880) <= 10718566;
srom_1(72881) <= 10161588;
srom_1(72882) <= 9596296;
srom_1(72883) <= 9025340;
srom_1(72884) <= 8451399;
srom_1(72885) <= 7877163;
srom_1(72886) <= 7305325;
srom_1(72887) <= 6738567;
srom_1(72888) <= 6179547;
srom_1(72889) <= 5630886;
srom_1(72890) <= 5095157;
srom_1(72891) <= 4574872;
srom_1(72892) <= 4072471;
srom_1(72893) <= 3590310;
srom_1(72894) <= 3130649;
srom_1(72895) <= 2695645;
srom_1(72896) <= 2287337;
srom_1(72897) <= 1907640;
srom_1(72898) <= 1558335;
srom_1(72899) <= 1241059;
srom_1(72900) <= 957301;
srom_1(72901) <= 708390;
srom_1(72902) <= 495494;
srom_1(72903) <= 319612;
srom_1(72904) <= 181569;
srom_1(72905) <= 82011;
srom_1(72906) <= 21405;
srom_1(72907) <= 36;
srom_1(72908) <= 18004;
srom_1(72909) <= 75225;
srom_1(72910) <= 171430;
srom_1(72911) <= 306168;
srom_1(72912) <= 478807;
srom_1(72913) <= 688539;
srom_1(72914) <= 934378;
srom_1(72915) <= 1215173;
srom_1(72916) <= 1529606;
srom_1(72917) <= 1876204;
srom_1(72918) <= 2253341;
srom_1(72919) <= 2659248;
srom_1(72920) <= 3092022;
srom_1(72921) <= 3549633;
srom_1(72922) <= 4029937;
srom_1(72923) <= 4530679;
srom_1(72924) <= 5049512;
srom_1(72925) <= 5584004;
srom_1(72926) <= 6131648;
srom_1(72927) <= 6689875;
srom_1(72928) <= 7256068;
srom_1(72929) <= 7827572;
srom_1(72930) <= 8401706;
srom_1(72931) <= 8975780;
srom_1(72932) <= 9547100;
srom_1(72933) <= 10112987;
srom_1(72934) <= 10670788;
srom_1(72935) <= 11217887;
srom_1(72936) <= 11751719;
srom_1(72937) <= 12269780;
srom_1(72938) <= 12769641;
srom_1(72939) <= 13248957;
srom_1(72940) <= 13705482;
srom_1(72941) <= 14137074;
srom_1(72942) <= 14541710;
srom_1(72943) <= 14917491;
srom_1(72944) <= 15262657;
srom_1(72945) <= 15575587;
srom_1(72946) <= 15854815;
srom_1(72947) <= 16099032;
srom_1(72948) <= 16307092;
srom_1(72949) <= 16478019;
srom_1(72950) <= 16611013;
srom_1(72951) <= 16705448;
srom_1(72952) <= 16760884;
srom_1(72953) <= 16777058;
srom_1(72954) <= 16753897;
srom_1(72955) <= 16691507;
srom_1(72956) <= 16590183;
srom_1(72957) <= 16450398;
srom_1(72958) <= 16272809;
srom_1(72959) <= 16058248;
srom_1(72960) <= 15807722;
srom_1(72961) <= 15522405;
srom_1(72962) <= 15203635;
srom_1(72963) <= 14852907;
srom_1(72964) <= 14471865;
srom_1(72965) <= 14062297;
srom_1(72966) <= 13626124;
srom_1(72967) <= 13165389;
srom_1(72968) <= 12682255;
srom_1(72969) <= 12178987;
srom_1(72970) <= 11657944;
srom_1(72971) <= 11121570;
srom_1(72972) <= 10572380;
srom_1(72973) <= 10012949;
srom_1(72974) <= 9445902;
srom_1(72975) <= 8873897;
srom_1(72976) <= 8299615;
srom_1(72977) <= 7725752;
srom_1(72978) <= 7154996;
srom_1(72979) <= 6590026;
srom_1(72980) <= 6033489;
srom_1(72981) <= 5487997;
srom_1(72982) <= 4956106;
srom_1(72983) <= 4440312;
srom_1(72984) <= 3943032;
srom_1(72985) <= 3466600;
srom_1(72986) <= 3013248;
srom_1(72987) <= 2585103;
srom_1(72988) <= 2184173;
srom_1(72989) <= 1812338;
srom_1(72990) <= 1471341;
srom_1(72991) <= 1162781;
srom_1(72992) <= 888106;
srom_1(72993) <= 648603;
srom_1(72994) <= 445396;
srom_1(72995) <= 279437;
srom_1(72996) <= 151505;
srom_1(72997) <= 62199;
srom_1(72998) <= 11939;
srom_1(72999) <= 960;
srom_1(73000) <= 29313;
srom_1(73001) <= 96866;
srom_1(73002) <= 203302;
srom_1(73003) <= 348122;
srom_1(73004) <= 530646;
srom_1(73005) <= 750019;
srom_1(73006) <= 1005212;
srom_1(73007) <= 1295028;
srom_1(73008) <= 1618108;
srom_1(73009) <= 1972938;
srom_1(73010) <= 2357853;
srom_1(73011) <= 2771048;
srom_1(73012) <= 3210585;
srom_1(73013) <= 3674405;
srom_1(73014) <= 4160330;
srom_1(73015) <= 4666084;
srom_1(73016) <= 5189294;
srom_1(73017) <= 5727506;
srom_1(73018) <= 6278198;
srom_1(73019) <= 6838785;
srom_1(73020) <= 7406641;
srom_1(73021) <= 7979101;
srom_1(73022) <= 8553481;
srom_1(73023) <= 9127089;
srom_1(73024) <= 9697233;
srom_1(73025) <= 10261241;
srom_1(73026) <= 10816467;
srom_1(73027) <= 11360308;
srom_1(73028) <= 11890214;
srom_1(73029) <= 12403700;
srom_1(73030) <= 12898357;
srom_1(73031) <= 13371867;
srom_1(73032) <= 13822008;
srom_1(73033) <= 14246671;
srom_1(73034) <= 14643863;
srom_1(73035) <= 15011721;
srom_1(73036) <= 15348522;
srom_1(73037) <= 15652686;
srom_1(73038) <= 15922785;
srom_1(73039) <= 16157555;
srom_1(73040) <= 16355893;
srom_1(73041) <= 16516869;
srom_1(73042) <= 16639730;
srom_1(73043) <= 16723898;
srom_1(73044) <= 16768979;
srom_1(73045) <= 16774761;
srom_1(73046) <= 16741218;
srom_1(73047) <= 16668507;
srom_1(73048) <= 16556969;
srom_1(73049) <= 16407126;
srom_1(73050) <= 16219682;
srom_1(73051) <= 15995515;
srom_1(73052) <= 15735676;
srom_1(73053) <= 15441385;
srom_1(73054) <= 15114021;
srom_1(73055) <= 14755119;
srom_1(73056) <= 14366362;
srom_1(73057) <= 13949573;
srom_1(73058) <= 13506708;
srom_1(73059) <= 13039841;
srom_1(73060) <= 12551164;
srom_1(73061) <= 12042967;
srom_1(73062) <= 11517633;
srom_1(73063) <= 10977626;
srom_1(73064) <= 10425478;
srom_1(73065) <= 9863779;
srom_1(73066) <= 9295162;
srom_1(73067) <= 8722294;
srom_1(73068) <= 8147861;
srom_1(73069) <= 7574558;
srom_1(73070) <= 7005071;
srom_1(73071) <= 6442073;
srom_1(73072) <= 5888202;
srom_1(73073) <= 5346057;
srom_1(73074) <= 4818179;
srom_1(73075) <= 4307044;
srom_1(73076) <= 3815049;
srom_1(73077) <= 3344501;
srom_1(73078) <= 2897606;
srom_1(73079) <= 2476461;
srom_1(73080) <= 2083040;
srom_1(73081) <= 1719188;
srom_1(73082) <= 1386611;
srom_1(73083) <= 1086868;
srom_1(73084) <= 821366;
srom_1(73085) <= 591350;
srom_1(73086) <= 397897;
srom_1(73087) <= 241916;
srom_1(73088) <= 124137;
srom_1(73089) <= 45114;
srom_1(73090) <= 5215;
srom_1(73091) <= 4630;
srom_1(73092) <= 43359;
srom_1(73093) <= 121223;
srom_1(73094) <= 237855;
srom_1(73095) <= 392708;
srom_1(73096) <= 585058;
srom_1(73097) <= 814000;
srom_1(73098) <= 1078463;
srom_1(73099) <= 1377205;
srom_1(73100) <= 1708827;
srom_1(73101) <= 2071772;
srom_1(73102) <= 2464339;
srom_1(73103) <= 2884687;
srom_1(73104) <= 3330844;
srom_1(73105) <= 3800719;
srom_1(73106) <= 4292109;
srom_1(73107) <= 4802708;
srom_1(73108) <= 5330123;
srom_1(73109) <= 5871880;
srom_1(73110) <= 6425439;
srom_1(73111) <= 6988203;
srom_1(73112) <= 7557535;
srom_1(73113) <= 8130764;
srom_1(73114) <= 8705202;
srom_1(73115) <= 9278156;
srom_1(73116) <= 9846938;
srom_1(73117) <= 10408881;
srom_1(73118) <= 10961351;
srom_1(73119) <= 11501756;
srom_1(73120) <= 12027562;
srom_1(73121) <= 12536305;
srom_1(73122) <= 13025597;
srom_1(73123) <= 13493145;
srom_1(73124) <= 13936756;
srom_1(73125) <= 14354349;
srom_1(73126) <= 14743968;
srom_1(73127) <= 15103783;
srom_1(73128) <= 15432109;
srom_1(73129) <= 15727406;
srom_1(73130) <= 15988289;
srom_1(73131) <= 16213534;
srom_1(73132) <= 16402085;
srom_1(73133) <= 16553058;
srom_1(73134) <= 16665745;
srom_1(73135) <= 16739618;
srom_1(73136) <= 16774330;
srom_1(73137) <= 16769719;
srom_1(73138) <= 16725806;
srom_1(73139) <= 16642797;
srom_1(73140) <= 16521081;
srom_1(73141) <= 16361229;
srom_1(73142) <= 16163990;
srom_1(73143) <= 15930291;
srom_1(73144) <= 15661225;
srom_1(73145) <= 15358056;
srom_1(73146) <= 15022205;
srom_1(73147) <= 14655247;
srom_1(73148) <= 14258902;
srom_1(73149) <= 13835029;
srom_1(73150) <= 13385616;
srom_1(73151) <= 12912770;
srom_1(73152) <= 12418710;
srom_1(73153) <= 11905750;
srom_1(73154) <= 11376298;
srom_1(73155) <= 10832835;
srom_1(73156) <= 10277910;
srom_1(73157) <= 9714126;
srom_1(73158) <= 9144126;
srom_1(73159) <= 8570583;
srom_1(73160) <= 7996186;
srom_1(73161) <= 7423630;
srom_1(73162) <= 6855599;
srom_1(73163) <= 6294757;
srom_1(73164) <= 5743733;
srom_1(73165) <= 5205113;
srom_1(73166) <= 4681420;
srom_1(73167) <= 4175112;
srom_1(73168) <= 3688563;
srom_1(73169) <= 3224054;
srom_1(73170) <= 2783763;
srom_1(73171) <= 2369755;
srom_1(73172) <= 1983971;
srom_1(73173) <= 1628221;
srom_1(73174) <= 1304173;
srom_1(73175) <= 1013346;
srom_1(73176) <= 757105;
srom_1(73177) <= 536650;
srom_1(73178) <= 353015;
srom_1(73179) <= 207062;
srom_1(73180) <= 99476;
srom_1(73181) <= 30760;
srom_1(73182) <= 1236;
srom_1(73183) <= 11044;
srom_1(73184) <= 60137;
srom_1(73185) <= 148286;
srom_1(73186) <= 275076;
srom_1(73187) <= 439913;
srom_1(73188) <= 642024;
srom_1(73189) <= 880462;
srom_1(73190) <= 1154107;
srom_1(73191) <= 1461678;
srom_1(73192) <= 1801732;
srom_1(73193) <= 2172674;
srom_1(73194) <= 2572764;
srom_1(73195) <= 3000127;
srom_1(73196) <= 3452759;
srom_1(73197) <= 3928536;
srom_1(73198) <= 4425228;
srom_1(73199) <= 4940506;
srom_1(73200) <= 5471953;
srom_1(73201) <= 6017077;
srom_1(73202) <= 6573322;
srom_1(73203) <= 7138080;
srom_1(73204) <= 7708702;
srom_1(73205) <= 8282512;
srom_1(73206) <= 8856819;
srom_1(73207) <= 9428931;
srom_1(73208) <= 9996165;
srom_1(73209) <= 10555860;
srom_1(73210) <= 11105392;
srom_1(73211) <= 11642184;
srom_1(73212) <= 12163720;
srom_1(73213) <= 12667552;
srom_1(73214) <= 13151319;
srom_1(73215) <= 13612751;
srom_1(73216) <= 14049687;
srom_1(73217) <= 14460075;
srom_1(73218) <= 14841992;
srom_1(73219) <= 15193647;
srom_1(73220) <= 15513391;
srom_1(73221) <= 15799724;
srom_1(73222) <= 16051304;
srom_1(73223) <= 16266951;
srom_1(73224) <= 16445653;
srom_1(73225) <= 16586574;
srom_1(73226) <= 16689051;
srom_1(73227) <= 16752605;
srom_1(73228) <= 16776937;
srom_1(73229) <= 16761933;
srom_1(73230) <= 16707664;
srom_1(73231) <= 16614384;
srom_1(73232) <= 16482530;
srom_1(73233) <= 16312721;
srom_1(73234) <= 16105754;
srom_1(73235) <= 15862598;
srom_1(73236) <= 15584394;
srom_1(73237) <= 15272446;
srom_1(73238) <= 14928218;
srom_1(73239) <= 14553323;
srom_1(73240) <= 14149519;
srom_1(73241) <= 13718701;
srom_1(73242) <= 13262888;
srom_1(73243) <= 12784218;
srom_1(73244) <= 12284936;
srom_1(73245) <= 11767382;
srom_1(73246) <= 11233984;
srom_1(73247) <= 10687243;
srom_1(73248) <= 10129723;
srom_1(73249) <= 9564038;
srom_1(73250) <= 8992842;
srom_1(73251) <= 8418811;
srom_1(73252) <= 7844639;
srom_1(73253) <= 7273018;
srom_1(73254) <= 6706629;
srom_1(73255) <= 6148127;
srom_1(73256) <= 5600131;
srom_1(73257) <= 5065211;
srom_1(73258) <= 4545876;
srom_1(73259) <= 4044560;
srom_1(73260) <= 3563616;
srom_1(73261) <= 3105297;
srom_1(73262) <= 2671754;
srom_1(73263) <= 2265019;
srom_1(73264) <= 1886999;
srom_1(73265) <= 1539468;
srom_1(73266) <= 1224055;
srom_1(73267) <= 942239;
srom_1(73268) <= 695341;
srom_1(73269) <= 484520;
srom_1(73270) <= 310764;
srom_1(73271) <= 174887;
srom_1(73272) <= 77528;
srom_1(73273) <= 19142;
srom_1(73274) <= 3;
srom_1(73275) <= 20201;
srom_1(73276) <= 79642;
srom_1(73277) <= 178046;
srom_1(73278) <= 314953;
srom_1(73279) <= 489719;
srom_1(73280) <= 701526;
srom_1(73281) <= 949381;
srom_1(73282) <= 1232120;
srom_1(73283) <= 1548419;
srom_1(73284) <= 1896794;
srom_1(73285) <= 2275611;
srom_1(73286) <= 2683094;
srom_1(73287) <= 3117332;
srom_1(73288) <= 3576289;
srom_1(73289) <= 4057813;
srom_1(73290) <= 4559645;
srom_1(73291) <= 5079432;
srom_1(73292) <= 5614738;
srom_1(73293) <= 6163051;
srom_1(73294) <= 6721800;
srom_1(73295) <= 7288366;
srom_1(73296) <= 7860091;
srom_1(73297) <= 8434294;
srom_1(73298) <= 9008283;
srom_1(73299) <= 9579366;
srom_1(73300) <= 10144866;
srom_1(73301) <= 10702130;
srom_1(73302) <= 11248544;
srom_1(73303) <= 11781548;
srom_1(73304) <= 12298641;
srom_1(73305) <= 12797398;
srom_1(73306) <= 13275481;
srom_1(73307) <= 13730648;
srom_1(73308) <= 14160764;
srom_1(73309) <= 14563813;
srom_1(73310) <= 14937903;
srom_1(73311) <= 15281282;
srom_1(73312) <= 15592339;
srom_1(73313) <= 15869615;
srom_1(73314) <= 16111810;
srom_1(73315) <= 16317788;
srom_1(73316) <= 16486584;
srom_1(73317) <= 16617405;
srom_1(73318) <= 16709639;
srom_1(73319) <= 16762853;
srom_1(73320) <= 16776797;
srom_1(73321) <= 16751405;
srom_1(73322) <= 16686798;
srom_1(73323) <= 16583278;
srom_1(73324) <= 16441330;
srom_1(73325) <= 16261620;
srom_1(73326) <= 16044990;
srom_1(73327) <= 15792458;
srom_1(73328) <= 15505206;
srom_1(73329) <= 15184582;
srom_1(73330) <= 14832089;
srom_1(73331) <= 14449381;
srom_1(73332) <= 14038251;
srom_1(73333) <= 13600629;
srom_1(73334) <= 13138565;
srom_1(73335) <= 12654227;
srom_1(73336) <= 12149887;
srom_1(73337) <= 11627908;
srom_1(73338) <= 11090739;
srom_1(73339) <= 10540899;
srom_1(73340) <= 9980966;
srom_1(73341) <= 9413566;
srom_1(73342) <= 8841360;
srom_1(73343) <= 8267030;
srom_1(73344) <= 7693271;
srom_1(73345) <= 7122772;
srom_1(73346) <= 6558209;
srom_1(73347) <= 6002230;
srom_1(73348) <= 5457441;
srom_1(73349) <= 4926397;
srom_1(73350) <= 4411589;
srom_1(73351) <= 3915430;
srom_1(73352) <= 3440248;
srom_1(73353) <= 2988270;
srom_1(73354) <= 2561617;
srom_1(73355) <= 2162288;
srom_1(73356) <= 1792156;
srom_1(73357) <= 1452957;
srom_1(73358) <= 1146282;
srom_1(73359) <= 873569;
srom_1(73360) <= 636097;
srom_1(73361) <= 434978;
srom_1(73362) <= 271157;
srom_1(73363) <= 145401;
srom_1(73364) <= 58301;
srom_1(73365) <= 10264;
srom_1(73366) <= 1516;
srom_1(73367) <= 32098;
srom_1(73368) <= 101867;
srom_1(73369) <= 210495;
srom_1(73370) <= 357473;
srom_1(73371) <= 542112;
srom_1(73372) <= 763545;
srom_1(73373) <= 1020736;
srom_1(73374) <= 1312476;
srom_1(73375) <= 1637399;
srom_1(73376) <= 1993981;
srom_1(73377) <= 2380550;
srom_1(73378) <= 2795292;
srom_1(73379) <= 3236263;
srom_1(73380) <= 3701395;
srom_1(73381) <= 4188508;
srom_1(73382) <= 4695316;
srom_1(73383) <= 5219443;
srom_1(73384) <= 5758431;
srom_1(73385) <= 6309753;
srom_1(73386) <= 6870824;
srom_1(73387) <= 7439012;
srom_1(73388) <= 8011653;
srom_1(73389) <= 8586061;
srom_1(73390) <= 9159544;
srom_1(73391) <= 9729412;
srom_1(73392) <= 10292992;
srom_1(73393) <= 10847642;
srom_1(73394) <= 11390760;
srom_1(73395) <= 11919800;
srom_1(73396) <= 12432282;
srom_1(73397) <= 12925801;
srom_1(73398) <= 13398044;
srom_1(73399) <= 13846795;
srom_1(73400) <= 14269952;
srom_1(73401) <= 14665529;
srom_1(73402) <= 15031671;
srom_1(73403) <= 15366661;
srom_1(73404) <= 15668929;
srom_1(73405) <= 15937057;
srom_1(73406) <= 16169788;
srom_1(73407) <= 16366030;
srom_1(73408) <= 16524864;
srom_1(73409) <= 16645543;
srom_1(73410) <= 16727503;
srom_1(73411) <= 16770359;
srom_1(73412) <= 16773910;
srom_1(73413) <= 16738140;
srom_1(73414) <= 16663216;
srom_1(73415) <= 16549489;
srom_1(73416) <= 16397493;
srom_1(73417) <= 16207940;
srom_1(73418) <= 15981720;
srom_1(73419) <= 15719894;
srom_1(73420) <= 15423688;
srom_1(73421) <= 15094493;
srom_1(73422) <= 14733851;
srom_1(73423) <= 14343454;
srom_1(73424) <= 13925133;
srom_1(73425) <= 13480850;
srom_1(73426) <= 13012687;
srom_1(73427) <= 12522840;
srom_1(73428) <= 12013606;
srom_1(73429) <= 11487373;
srom_1(73430) <= 10946610;
srom_1(73431) <= 10393850;
srom_1(73432) <= 9831688;
srom_1(73433) <= 9262758;
srom_1(73434) <= 8689730;
srom_1(73435) <= 8115289;
srom_1(73436) <= 7542130;
srom_1(73437) <= 6972940;
srom_1(73438) <= 6410389;
srom_1(73439) <= 5857114;
srom_1(73440) <= 5315711;
srom_1(73441) <= 4788717;
srom_1(73442) <= 4278604;
srom_1(73443) <= 3787765;
srom_1(73444) <= 3318501;
srom_1(73445) <= 2873012;
srom_1(73446) <= 2453387;
srom_1(73447) <= 2061595;
srom_1(73448) <= 1699472;
srom_1(73449) <= 1368717;
srom_1(73450) <= 1070881;
srom_1(73451) <= 807360;
srom_1(73452) <= 579390;
srom_1(73453) <= 388040;
srom_1(73454) <= 234208;
srom_1(73455) <= 118614;
srom_1(73456) <= 41801;
srom_1(73457) <= 4130;
srom_1(73458) <= 5775;
srom_1(73459) <= 46731;
srom_1(73460) <= 126805;
srom_1(73461) <= 245621;
srom_1(73462) <= 402623;
srom_1(73463) <= 597073;
srom_1(73464) <= 828061;
srom_1(73465) <= 1094503;
srom_1(73466) <= 1395149;
srom_1(73467) <= 1728590;
srom_1(73468) <= 2093262;
srom_1(73469) <= 2487455;
srom_1(73470) <= 2909321;
srom_1(73471) <= 3356881;
srom_1(73472) <= 3828036;
srom_1(73473) <= 4320577;
srom_1(73474) <= 4832195;
srom_1(73475) <= 5360490;
srom_1(73476) <= 5902985;
srom_1(73477) <= 6457136;
srom_1(73478) <= 7020344;
srom_1(73479) <= 7589969;
srom_1(73480) <= 8163338;
srom_1(73481) <= 8737764;
srom_1(73482) <= 9310553;
srom_1(73483) <= 9879018;
srom_1(73484) <= 10440494;
srom_1(73485) <= 10992349;
srom_1(73486) <= 11531993;
srom_1(73487) <= 12056897;
srom_1(73488) <= 12564599;
srom_1(73489) <= 13052718;
srom_1(73490) <= 13518966;
srom_1(73491) <= 13961156;
srom_1(73492) <= 14377214;
srom_1(73493) <= 14765190;
srom_1(73494) <= 15123263;
srom_1(73495) <= 15449756;
srom_1(73496) <= 15743136;
srom_1(73497) <= 16002028;
srom_1(73498) <= 16225219;
srom_1(73499) <= 16411660;
srom_1(73500) <= 16560479;
srom_1(73501) <= 16670978;
srom_1(73502) <= 16742637;
srom_1(73503) <= 16775121;
srom_1(73504) <= 16768279;
srom_1(73505) <= 16722141;
srom_1(73506) <= 16636924;
srom_1(73507) <= 16513028;
srom_1(73508) <= 16351034;
srom_1(73509) <= 16151701;
srom_1(73510) <= 15915965;
srom_1(73511) <= 15644930;
srom_1(73512) <= 15339867;
srom_1(73513) <= 15002208;
srom_1(73514) <= 14633536;
srom_1(73515) <= 14235578;
srom_1(73516) <= 13810203;
srom_1(73517) <= 13359403;
srom_1(73518) <= 12885294;
srom_1(73519) <= 12390099;
srom_1(73520) <= 11876138;
srom_1(73521) <= 11345824;
srom_1(73522) <= 10801642;
srom_1(73523) <= 10246145;
srom_1(73524) <= 9681937;
srom_1(73525) <= 9111665;
srom_1(73526) <= 8538001;
srom_1(73527) <= 7963637;
srom_1(73528) <= 7391266;
srom_1(73529) <= 6823572;
srom_1(73530) <= 6263216;
srom_1(73531) <= 5712828;
srom_1(73532) <= 5174987;
srom_1(73533) <= 4652215;
srom_1(73534) <= 4146965;
srom_1(73535) <= 3661606;
srom_1(73536) <= 3198413;
srom_1(73537) <= 2759559;
srom_1(73538) <= 2347101;
srom_1(73539) <= 1962974;
srom_1(73540) <= 1608979;
srom_1(73541) <= 1286776;
srom_1(73542) <= 997875;
srom_1(73543) <= 743633;
srom_1(73544) <= 525240;
srom_1(73545) <= 343722;
srom_1(73546) <= 199928;
srom_1(73547) <= 94534;
srom_1(73548) <= 28034;
srom_1(73549) <= 740;
srom_1(73550) <= 12779;
srom_1(73551) <= 64095;
srom_1(73552) <= 154448;
srom_1(73553) <= 283414;
srom_1(73554) <= 450387;
srom_1(73555) <= 654586;
srom_1(73556) <= 895052;
srom_1(73557) <= 1170658;
srom_1(73558) <= 1480111;
srom_1(73559) <= 1821961;
srom_1(73560) <= 2194604;
srom_1(73561) <= 2596293;
srom_1(73562) <= 3025143;
srom_1(73563) <= 3479145;
srom_1(73564) <= 3956170;
srom_1(73565) <= 4453979;
srom_1(73566) <= 4970239;
srom_1(73567) <= 5502529;
srom_1(73568) <= 6048353;
srom_1(73569) <= 6605151;
srom_1(73570) <= 7170313;
srom_1(73571) <= 7741187;
srom_1(73572) <= 8315098;
srom_1(73573) <= 8889353;
srom_1(73574) <= 9461260;
srom_1(73575) <= 10028137;
srom_1(73576) <= 10587325;
srom_1(73577) <= 11136203;
srom_1(73578) <= 11672197;
srom_1(73579) <= 12192792;
srom_1(73580) <= 12695549;
srom_1(73581) <= 13178109;
srom_1(73582) <= 13638209;
srom_1(73583) <= 14073692;
srom_1(73584) <= 14482516;
srom_1(73585) <= 14862763;
srom_1(73586) <= 15212651;
srom_1(73587) <= 15530538;
srom_1(73588) <= 15814935;
srom_1(73589) <= 16064506;
srom_1(73590) <= 16278083;
srom_1(73591) <= 16454664;
srom_1(73592) <= 16593420;
srom_1(73593) <= 16693701;
srom_1(73594) <= 16755036;
srom_1(73595) <= 16777138;
srom_1(73596) <= 16759904;
srom_1(73597) <= 16703413;
srom_1(73598) <= 16607932;
srom_1(73599) <= 16473907;
srom_1(73600) <= 16301968;
srom_1(73601) <= 16092920;
srom_1(73602) <= 15847744;
srom_1(73603) <= 15567590;
srom_1(73604) <= 15253771;
srom_1(73605) <= 14907759;
srom_1(73606) <= 14531176;
srom_1(73607) <= 14125788;
srom_1(73608) <= 13693497;
srom_1(73609) <= 13236330;
srom_1(73610) <= 12756430;
srom_1(73611) <= 12256047;
srom_1(73612) <= 11737529;
srom_1(73613) <= 11203307;
srom_1(73614) <= 10655885;
srom_1(73615) <= 10097832;
srom_1(73616) <= 9531763;
srom_1(73617) <= 8960334;
srom_1(73618) <= 8386224;
srom_1(73619) <= 7812124;
srom_1(73620) <= 7240729;
srom_1(73621) <= 6674716;
srom_1(73622) <= 6116740;
srom_1(73623) <= 5569417;
srom_1(73624) <= 5035315;
srom_1(73625) <= 4516937;
srom_1(73626) <= 4016715;
srom_1(73627) <= 3536995;
srom_1(73628) <= 3080025;
srom_1(73629) <= 2647949;
srom_1(73630) <= 2242793;
srom_1(73631) <= 1866456;
srom_1(73632) <= 1520705;
srom_1(73633) <= 1207159;
srom_1(73634) <= 927289;
srom_1(73635) <= 682409;
srom_1(73636) <= 473665;
srom_1(73637) <= 302037;
srom_1(73638) <= 168330;
srom_1(73639) <= 73170;
srom_1(73640) <= 17005;
srom_1(73641) <= 96;
srom_1(73642) <= 22525;
srom_1(73643) <= 84185;
srom_1(73644) <= 184787;
srom_1(73645) <= 323859;
srom_1(73646) <= 500750;
srom_1(73647) <= 714630;
srom_1(73648) <= 964496;
srom_1(73649) <= 1249176;
srom_1(73650) <= 1567335;
srom_1(73651) <= 1917482;
srom_1(73652) <= 2297973;
srom_1(73653) <= 2707026;
srom_1(73654) <= 3142722;
srom_1(73655) <= 3603018;
srom_1(73656) <= 4085755;
srom_1(73657) <= 4588669;
srom_1(73658) <= 5109402;
srom_1(73659) <= 5645513;
srom_1(73660) <= 6194488;
srom_1(73661) <= 6753751;
srom_1(73662) <= 7320680;
srom_1(73663) <= 7892618;
srom_1(73664) <= 8466881;
srom_1(73665) <= 9040777;
srom_1(73666) <= 9611615;
srom_1(73667) <= 10176718;
srom_1(73668) <= 10733436;
srom_1(73669) <= 11279158;
srom_1(73670) <= 11811325;
srom_1(73671) <= 12327442;
srom_1(73672) <= 12825089;
srom_1(73673) <= 13301931;
srom_1(73674) <= 13755733;
srom_1(73675) <= 14184367;
srom_1(73676) <= 14585822;
srom_1(73677) <= 14958217;
srom_1(73678) <= 15299804;
srom_1(73679) <= 15608982;
srom_1(73680) <= 15884302;
srom_1(73681) <= 16124472;
srom_1(73682) <= 16328365;
srom_1(73683) <= 16495026;
srom_1(73684) <= 16623674;
srom_1(73685) <= 16713704;
srom_1(73686) <= 16764696;
srom_1(73687) <= 16776408;
srom_1(73688) <= 16748788;
srom_1(73689) <= 16681964;
srom_1(73690) <= 16576249;
srom_1(73691) <= 16432140;
srom_1(73692) <= 16250312;
srom_1(73693) <= 16031617;
srom_1(73694) <= 15777082;
srom_1(73695) <= 15487900;
srom_1(73696) <= 15165427;
srom_1(73697) <= 14811174;
srom_1(73698) <= 14426805;
srom_1(73699) <= 14014120;
srom_1(73700) <= 13575055;
srom_1(73701) <= 13111669;
srom_1(73702) <= 12626135;
srom_1(73703) <= 12120730;
srom_1(73704) <= 11597824;
srom_1(73705) <= 11059868;
srom_1(73706) <= 10509386;
srom_1(73707) <= 9948959;
srom_1(73708) <= 9381215;
srom_1(73709) <= 8808816;
srom_1(73710) <= 8234447;
srom_1(73711) <= 7660800;
srom_1(73712) <= 7090567;
srom_1(73713) <= 6526421;
srom_1(73714) <= 5971007;
srom_1(73715) <= 5426929;
srom_1(73716) <= 4896741;
srom_1(73717) <= 4382926;
srom_1(73718) <= 3887896;
srom_1(73719) <= 3413971;
srom_1(73720) <= 2963374;
srom_1(73721) <= 2538218;
srom_1(73722) <= 2140496;
srom_1(73723) <= 1772074;
srom_1(73724) <= 1434679;
srom_1(73725) <= 1129893;
srom_1(73726) <= 859146;
srom_1(73727) <= 623707;
srom_1(73728) <= 424681;
srom_1(73729) <= 263000;
srom_1(73730) <= 139422;
srom_1(73731) <= 54528;
srom_1(73732) <= 8716;
srom_1(73733) <= 2199;
srom_1(73734) <= 35010;
srom_1(73735) <= 106993;
srom_1(73736) <= 217811;
srom_1(73737) <= 366945;
srom_1(73738) <= 553696;
srom_1(73739) <= 777187;
srom_1(73740) <= 1036371;
srom_1(73741) <= 1330031;
srom_1(73742) <= 1656792;
srom_1(73743) <= 2015121;
srom_1(73744) <= 2403337;
srom_1(73745) <= 2819620;
srom_1(73746) <= 3262018;
srom_1(73747) <= 3728457;
srom_1(73748) <= 4216748;
srom_1(73749) <= 4724603;
srom_1(73750) <= 5249639;
srom_1(73751) <= 5789395;
srom_1(73752) <= 6341340;
srom_1(73753) <= 6902885;
srom_1(73754) <= 7471397;
srom_1(73755) <= 8044210;
srom_1(73756) <= 8618639;
srom_1(73757) <= 9191988;
srom_1(73758) <= 9761570;
srom_1(73759) <= 10324714;
srom_1(73760) <= 10878779;
srom_1(73761) <= 11421167;
srom_1(73762) <= 11949334;
srom_1(73763) <= 12460803;
srom_1(73764) <= 12953176;
srom_1(73765) <= 13424145;
srom_1(73766) <= 13871500;
srom_1(73767) <= 14293144;
srom_1(73768) <= 14687100;
srom_1(73769) <= 15051520;
srom_1(73770) <= 15384695;
srom_1(73771) <= 15685063;
srom_1(73772) <= 15951215;
srom_1(73773) <= 16181904;
srom_1(73774) <= 16376048;
srom_1(73775) <= 16532735;
srom_1(73776) <= 16651232;
srom_1(73777) <= 16730983;
srom_1(73778) <= 16771613;
srom_1(73779) <= 16772933;
srom_1(73780) <= 16734935;
srom_1(73781) <= 16657799;
srom_1(73782) <= 16541886;
srom_1(73783) <= 16387739;
srom_1(73784) <= 16196081;
srom_1(73785) <= 15967812;
srom_1(73786) <= 15704001;
srom_1(73787) <= 15405885;
srom_1(73788) <= 15074864;
srom_1(73789) <= 14712488;
srom_1(73790) <= 14320457;
srom_1(73791) <= 13900610;
srom_1(73792) <= 13454915;
srom_1(73793) <= 12985462;
srom_1(73794) <= 12494453;
srom_1(73795) <= 11984191;
srom_1(73796) <= 11457067;
srom_1(73797) <= 10915555;
srom_1(73798) <= 10362192;
srom_1(73799) <= 9799575;
srom_1(73800) <= 9230342;
srom_1(73801) <= 8657161;
srom_1(73802) <= 8082721;
srom_1(73803) <= 7509715;
srom_1(73804) <= 6940830;
srom_1(73805) <= 6378735;
srom_1(73806) <= 5826065;
srom_1(73807) <= 5285411;
srom_1(73808) <= 4759310;
srom_1(73809) <= 4250227;
srom_1(73810) <= 3760551;
srom_1(73811) <= 3292577;
srom_1(73812) <= 2848500;
srom_1(73813) <= 2430403;
srom_1(73814) <= 2040246;
srom_1(73815) <= 1679858;
srom_1(73816) <= 1350930;
srom_1(73817) <= 1055004;
srom_1(73818) <= 793468;
srom_1(73819) <= 567548;
srom_1(73820) <= 378304;
srom_1(73821) <= 226623;
srom_1(73822) <= 113216;
srom_1(73823) <= 38615;
srom_1(73824) <= 3170;
srom_1(73825) <= 7048;
srom_1(73826) <= 50229;
srom_1(73827) <= 132512;
srom_1(73828) <= 253511;
srom_1(73829) <= 412658;
srom_1(73830) <= 609207;
srom_1(73831) <= 842236;
srom_1(73832) <= 1110652;
srom_1(73833) <= 1413198;
srom_1(73834) <= 1748454;
srom_1(73835) <= 2114847;
srom_1(73836) <= 2510660;
srom_1(73837) <= 2934038;
srom_1(73838) <= 3382993;
srom_1(73839) <= 3855421;
srom_1(73840) <= 4349107;
srom_1(73841) <= 4861736;
srom_1(73842) <= 5390904;
srom_1(73843) <= 5934128;
srom_1(73844) <= 6488863;
srom_1(73845) <= 7052506;
srom_1(73846) <= 7622415;
srom_1(73847) <= 8195916;
srom_1(73848) <= 8770321;
srom_1(73849) <= 9342936;
srom_1(73850) <= 9911076;
srom_1(73851) <= 10472077;
srom_1(73852) <= 11023307;
srom_1(73853) <= 11562183;
srom_1(73854) <= 12086176;
srom_1(73855) <= 12592830;
srom_1(73856) <= 13079769;
srom_1(73857) <= 13544710;
srom_1(73858) <= 13985472;
srom_1(73859) <= 14399988;
srom_1(73860) <= 14786315;
srom_1(73861) <= 15142641;
srom_1(73862) <= 15467295;
srom_1(73863) <= 15758755;
srom_1(73864) <= 16015653;
srom_1(73865) <= 16236785;
srom_1(73866) <= 16421115;
srom_1(73867) <= 16567778;
srom_1(73868) <= 16676085;
srom_1(73869) <= 16745530;
srom_1(73870) <= 16775786;
srom_1(73871) <= 16766712;
srom_1(73872) <= 16718350;
srom_1(73873) <= 16630927;
srom_1(73874) <= 16504853;
srom_1(73875) <= 16340719;
srom_1(73876) <= 16139295;
srom_1(73877) <= 15901525;
srom_1(73878) <= 15628525;
srom_1(73879) <= 15321574;
srom_1(73880) <= 14982112;
srom_1(73881) <= 14611731;
srom_1(73882) <= 14212167;
srom_1(73883) <= 13785295;
srom_1(73884) <= 13333116;
srom_1(73885) <= 12857750;
srom_1(73886) <= 12361427;
srom_1(73887) <= 11846474;
srom_1(73888) <= 11315306;
srom_1(73889) <= 10770414;
srom_1(73890) <= 10214352;
srom_1(73891) <= 9649729;
srom_1(73892) <= 9079193;
srom_1(73893) <= 8505417;
srom_1(73894) <= 7931094;
srom_1(73895) <= 7358917;
srom_1(73896) <= 6791568;
srom_1(73897) <= 6231708;
srom_1(73898) <= 5681962;
srom_1(73899) <= 5144909;
srom_1(73900) <= 4623067;
srom_1(73901) <= 4118883;
srom_1(73902) <= 3634720;
srom_1(73903) <= 3172851;
srom_1(73904) <= 2735440;
srom_1(73905) <= 2324538;
srom_1(73906) <= 1942073;
srom_1(73907) <= 1589838;
srom_1(73908) <= 1269485;
srom_1(73909) <= 982516;
srom_1(73910) <= 730276;
srom_1(73911) <= 513950;
srom_1(73912) <= 334550;
srom_1(73913) <= 192918;
srom_1(73914) <= 89718;
srom_1(73915) <= 25435;
srom_1(73916) <= 370;
srom_1(73917) <= 14640;
srom_1(73918) <= 68179;
srom_1(73919) <= 160735;
srom_1(73920) <= 291874;
srom_1(73921) <= 460981;
srom_1(73922) <= 667264;
srom_1(73923) <= 909755;
srom_1(73924) <= 1187317;
srom_1(73925) <= 1498648;
srom_1(73926) <= 1842289;
srom_1(73927) <= 2216627;
srom_1(73928) <= 2619908;
srom_1(73929) <= 3050240;
srom_1(73930) <= 3505606;
srom_1(73931) <= 3983870;
srom_1(73932) <= 4482789;
srom_1(73933) <= 5000024;
srom_1(73934) <= 5533149;
srom_1(73935) <= 6079665;
srom_1(73936) <= 6637008;
srom_1(73937) <= 7202564;
srom_1(73938) <= 7773683;
srom_1(73939) <= 8347685;
srom_1(73940) <= 8921879;
srom_1(73941) <= 9493572;
srom_1(73942) <= 10060083;
srom_1(73943) <= 10618757;
srom_1(73944) <= 11166972;
srom_1(73945) <= 11702159;
srom_1(73946) <= 12221808;
srom_1(73947) <= 12723481;
srom_1(73948) <= 13204827;
srom_1(73949) <= 13663587;
srom_1(73950) <= 14097612;
srom_1(73951) <= 14504865;
srom_1(73952) <= 14883436;
srom_1(73953) <= 15231552;
srom_1(73954) <= 15547578;
srom_1(73955) <= 15830033;
srom_1(73956) <= 16077593;
srom_1(73957) <= 16289097;
srom_1(73958) <= 16463553;
srom_1(73959) <= 16600142;
srom_1(73960) <= 16698225;
srom_1(73961) <= 16757341;
srom_1(73962) <= 16777213;
srom_1(73963) <= 16757748;
srom_1(73964) <= 16699037;
srom_1(73965) <= 16601356;
srom_1(73966) <= 16465163;
srom_1(73967) <= 16291095;
srom_1(73968) <= 16079971;
srom_1(73969) <= 15832779;
srom_1(73970) <= 15550678;
srom_1(73971) <= 15234992;
srom_1(73972) <= 14887201;
srom_1(73973) <= 14508936;
srom_1(73974) <= 14101971;
srom_1(73975) <= 13668213;
srom_1(73976) <= 13209698;
srom_1(73977) <= 12728575;
srom_1(73978) <= 12227100;
srom_1(73979) <= 11707626;
srom_1(73980) <= 11172587;
srom_1(73981) <= 10624493;
srom_1(73982) <= 10065915;
srom_1(73983) <= 9499471;
srom_1(73984) <= 8927818;
srom_1(73985) <= 8353636;
srom_1(73986) <= 7779618;
srom_1(73987) <= 7208456;
srom_1(73988) <= 6642828;
srom_1(73989) <= 6085387;
srom_1(73990) <= 5538746;
srom_1(73991) <= 5005469;
srom_1(73992) <= 4488057;
srom_1(73993) <= 3988936;
srom_1(73994) <= 3510447;
srom_1(73995) <= 3054832;
srom_1(73996) <= 2624230;
srom_1(73997) <= 2220659;
srom_1(73998) <= 1846012;
srom_1(73999) <= 1502045;
srom_1(74000) <= 1190371;
srom_1(74001) <= 912453;
srom_1(74002) <= 669592;
srom_1(74003) <= 462929;
srom_1(74004) <= 293432;
srom_1(74005) <= 161896;
srom_1(74006) <= 68938;
srom_1(74007) <= 14994;
srom_1(74008) <= 316;
srom_1(74009) <= 24974;
srom_1(74010) <= 88852;
srom_1(74011) <= 191651;
srom_1(74012) <= 332888;
srom_1(74013) <= 511900;
srom_1(74014) <= 727850;
srom_1(74015) <= 979723;
srom_1(74016) <= 1266339;
srom_1(74017) <= 1586354;
srom_1(74018) <= 1938267;
srom_1(74019) <= 2320428;
srom_1(74020) <= 2731044;
srom_1(74021) <= 3168191;
srom_1(74022) <= 3629818;
srom_1(74023) <= 4113761;
srom_1(74024) <= 4617750;
srom_1(74025) <= 5139422;
srom_1(74026) <= 5676330;
srom_1(74027) <= 6225957;
srom_1(74028) <= 6785726;
srom_1(74029) <= 7353011;
srom_1(74030) <= 7925152;
srom_1(74031) <= 8499467;
srom_1(74032) <= 9073261;
srom_1(74033) <= 9643846;
srom_1(74034) <= 10208543;
srom_1(74035) <= 10764707;
srom_1(74036) <= 11309728;
srom_1(74037) <= 11841051;
srom_1(74038) <= 12356185;
srom_1(74039) <= 12852713;
srom_1(74040) <= 13328307;
srom_1(74041) <= 13780737;
srom_1(74042) <= 14207882;
srom_1(74043) <= 14607738;
srom_1(74044) <= 14978431;
srom_1(74045) <= 15318222;
srom_1(74046) <= 15625517;
srom_1(74047) <= 15898876;
srom_1(74048) <= 16137016;
srom_1(74049) <= 16338822;
srom_1(74050) <= 16503347;
srom_1(74051) <= 16629818;
srom_1(74052) <= 16717644;
srom_1(74053) <= 16766412;
srom_1(74054) <= 16775894;
srom_1(74055) <= 16746044;
srom_1(74056) <= 16677004;
srom_1(74057) <= 16569097;
srom_1(74058) <= 16422829;
srom_1(74059) <= 16238885;
srom_1(74060) <= 16018129;
srom_1(74061) <= 15761595;
srom_1(74062) <= 15470487;
srom_1(74063) <= 15146169;
srom_1(74064) <= 14790163;
srom_1(74065) <= 14404138;
srom_1(74066) <= 13989904;
srom_1(74067) <= 13549403;
srom_1(74068) <= 13084702;
srom_1(74069) <= 12597979;
srom_1(74070) <= 12091517;
srom_1(74071) <= 11567691;
srom_1(74072) <= 11028957;
srom_1(74073) <= 10477841;
srom_1(74074) <= 9916928;
srom_1(74075) <= 9348849;
srom_1(74076) <= 8776266;
srom_1(74077) <= 8201866;
srom_1(74078) <= 7628341;
srom_1(74079) <= 7058382;
srom_1(74080) <= 6494660;
srom_1(74081) <= 5939820;
srom_1(74082) <= 5396463;
srom_1(74083) <= 4867137;
srom_1(74084) <= 4354324;
srom_1(74085) <= 3860430;
srom_1(74086) <= 3387770;
srom_1(74087) <= 2938560;
srom_1(74088) <= 2514908;
srom_1(74089) <= 2118799;
srom_1(74090) <= 1752092;
srom_1(74091) <= 1416505;
srom_1(74092) <= 1113614;
srom_1(74093) <= 844837;
srom_1(74094) <= 611435;
srom_1(74095) <= 414503;
srom_1(74096) <= 254965;
srom_1(74097) <= 133568;
srom_1(74098) <= 50882;
srom_1(74099) <= 7294;
srom_1(74100) <= 3009;
srom_1(74101) <= 38047;
srom_1(74102) <= 112243;
srom_1(74103) <= 225251;
srom_1(74104) <= 376539;
srom_1(74105) <= 565398;
srom_1(74106) <= 790943;
srom_1(74107) <= 1052117;
srom_1(74108) <= 1347693;
srom_1(74109) <= 1676287;
srom_1(74110) <= 2036357;
srom_1(74111) <= 2426215;
srom_1(74112) <= 2844033;
srom_1(74113) <= 3287851;
srom_1(74114) <= 3755588;
srom_1(74115) <= 4245052;
srom_1(74116) <= 4753945;
srom_1(74117) <= 5279883;
srom_1(74118) <= 5820399;
srom_1(74119) <= 6372958;
srom_1(74120) <= 6934969;
srom_1(74121) <= 7503797;
srom_1(74122) <= 8076773;
srom_1(74123) <= 8651212;
srom_1(74124) <= 9224420;
srom_1(74125) <= 9793708;
srom_1(74126) <= 10356408;
srom_1(74127) <= 10909879;
srom_1(74128) <= 11451528;
srom_1(74129) <= 11978813;
srom_1(74130) <= 12489263;
srom_1(74131) <= 12980483;
srom_1(74132) <= 13450170;
srom_1(74133) <= 13896122;
srom_1(74134) <= 14316247;
srom_1(74135) <= 14708576;
srom_1(74136) <= 15071268;
srom_1(74137) <= 15402623;
srom_1(74138) <= 15701086;
srom_1(74139) <= 15965259;
srom_1(74140) <= 16193903;
srom_1(74141) <= 16385944;
srom_1(74142) <= 16540484;
srom_1(74143) <= 16656796;
srom_1(74144) <= 16734336;
srom_1(74145) <= 16772740;
srom_1(74146) <= 16771828;
srom_1(74147) <= 16731605;
srom_1(74148) <= 16652258;
srom_1(74149) <= 16534159;
srom_1(74150) <= 16377864;
srom_1(74151) <= 16184104;
srom_1(74152) <= 15953789;
srom_1(74153) <= 15687997;
srom_1(74154) <= 15387977;
srom_1(74155) <= 15055134;
srom_1(74156) <= 14691029;
srom_1(74157) <= 14297370;
srom_1(74158) <= 13876003;
srom_1(74159) <= 13428903;
srom_1(74160) <= 12958168;
srom_1(74161) <= 12466005;
srom_1(74162) <= 11954721;
srom_1(74163) <= 11426715;
srom_1(74164) <= 10884461;
srom_1(74165) <= 10330504;
srom_1(74166) <= 9767441;
srom_1(74167) <= 9197912;
srom_1(74168) <= 8624588;
srom_1(74169) <= 8050157;
srom_1(74170) <= 7477313;
srom_1(74171) <= 6908743;
srom_1(74172) <= 6347112;
srom_1(74173) <= 5795054;
srom_1(74174) <= 5255159;
srom_1(74175) <= 4729957;
srom_1(74176) <= 4221912;
srom_1(74177) <= 3733406;
srom_1(74178) <= 3266730;
srom_1(74179) <= 2824072;
srom_1(74180) <= 2407508;
srom_1(74181) <= 2018992;
srom_1(74182) <= 1660345;
srom_1(74183) <= 1333249;
srom_1(74184) <= 1039238;
srom_1(74185) <= 779691;
srom_1(74186) <= 555824;
srom_1(74187) <= 368688;
srom_1(74188) <= 219161;
srom_1(74189) <= 107942;
srom_1(74190) <= 35555;
srom_1(74191) <= 2338;
srom_1(74192) <= 8447;
srom_1(74193) <= 53853;
srom_1(74194) <= 138344;
srom_1(74195) <= 261523;
srom_1(74196) <= 422813;
srom_1(74197) <= 621457;
srom_1(74198) <= 856524;
srom_1(74199) <= 1126912;
srom_1(74200) <= 1431352;
srom_1(74201) <= 1768417;
srom_1(74202) <= 2136527;
srom_1(74203) <= 2533955;
srom_1(74204) <= 2958837;
srom_1(74205) <= 3409181;
srom_1(74206) <= 3882875;
srom_1(74207) <= 4377699;
srom_1(74208) <= 4891330;
srom_1(74209) <= 5421362;
srom_1(74210) <= 5965308;
srom_1(74211) <= 6520618;
srom_1(74212) <= 7084688;
srom_1(74213) <= 7654872;
srom_1(74214) <= 8228497;
srom_1(74215) <= 8802872;
srom_1(74216) <= 9375305;
srom_1(74217) <= 9943111;
srom_1(74218) <= 10503628;
srom_1(74219) <= 11054226;
srom_1(74220) <= 11592324;
srom_1(74221) <= 12115399;
srom_1(74222) <= 12620998;
srom_1(74223) <= 13106750;
srom_1(74224) <= 13570376;
srom_1(74225) <= 14009704;
srom_1(74226) <= 14422672;
srom_1(74227) <= 14807345;
srom_1(74228) <= 15161917;
srom_1(74229) <= 15484728;
srom_1(74230) <= 15774262;
srom_1(74231) <= 16029162;
srom_1(74232) <= 16248234;
srom_1(74233) <= 16430448;
srom_1(74234) <= 16574952;
srom_1(74235) <= 16681067;
srom_1(74236) <= 16748296;
srom_1(74237) <= 16776324;
srom_1(74238) <= 16765018;
srom_1(74239) <= 16714433;
srom_1(74240) <= 16624805;
srom_1(74241) <= 16496555;
srom_1(74242) <= 16330284;
srom_1(74243) <= 16126771;
srom_1(74244) <= 15886972;
srom_1(74245) <= 15612010;
srom_1(74246) <= 15303175;
srom_1(74247) <= 14961916;
srom_1(74248) <= 14589832;
srom_1(74249) <= 14188668;
srom_1(74250) <= 13760305;
srom_1(74251) <= 13306753;
srom_1(74252) <= 12830139;
srom_1(74253) <= 12332696;
srom_1(74254) <= 11816758;
srom_1(74255) <= 11284744;
srom_1(74256) <= 10739149;
srom_1(74257) <= 10182532;
srom_1(74258) <= 9617503;
srom_1(74259) <= 9046710;
srom_1(74260) <= 8472832;
srom_1(74261) <= 7898559;
srom_1(74262) <= 7326583;
srom_1(74263) <= 6759588;
srom_1(74264) <= 6200232;
srom_1(74265) <= 5651138;
srom_1(74266) <= 5114881;
srom_1(74267) <= 4593975;
srom_1(74268) <= 4090864;
srom_1(74269) <= 3607907;
srom_1(74270) <= 3147367;
srom_1(74271) <= 2711406;
srom_1(74272) <= 2302067;
srom_1(74273) <= 1921270;
srom_1(74274) <= 1570801;
srom_1(74275) <= 1252302;
srom_1(74276) <= 967268;
srom_1(74277) <= 717036;
srom_1(74278) <= 502778;
srom_1(74279) <= 325499;
srom_1(74280) <= 186031;
srom_1(74281) <= 85028;
srom_1(74282) <= 22963;
srom_1(74283) <= 127;
srom_1(74284) <= 16628;
srom_1(74285) <= 72388;
srom_1(74286) <= 167146;
srom_1(74287) <= 300456;
srom_1(74288) <= 471695;
srom_1(74289) <= 680059;
srom_1(74290) <= 924571;
srom_1(74291) <= 1204085;
srom_1(74292) <= 1517289;
srom_1(74293) <= 1862715;
srom_1(74294) <= 2238744;
srom_1(74295) <= 2643611;
srom_1(74296) <= 3075418;
srom_1(74297) <= 3532141;
srom_1(74298) <= 4011637;
srom_1(74299) <= 4511659;
srom_1(74300) <= 5029861;
srom_1(74301) <= 5563813;
srom_1(74302) <= 6111011;
srom_1(74303) <= 6668890;
srom_1(74304) <= 7234834;
srom_1(74305) <= 7806187;
srom_1(74306) <= 8380272;
srom_1(74307) <= 8954396;
srom_1(74308) <= 9525867;
srom_1(74309) <= 10092005;
srom_1(74310) <= 10650155;
srom_1(74311) <= 11197700;
srom_1(74312) <= 11732072;
srom_1(74313) <= 12250765;
srom_1(74314) <= 12751348;
srom_1(74315) <= 13231472;
srom_1(74316) <= 13688886;
srom_1(74317) <= 14121445;
srom_1(74318) <= 14527121;
srom_1(74319) <= 14904012;
srom_1(74320) <= 15250349;
srom_1(74321) <= 15564510;
srom_1(74322) <= 15845020;
srom_1(74323) <= 16090564;
srom_1(74324) <= 16299991;
srom_1(74325) <= 16472320;
srom_1(74326) <= 16606740;
srom_1(74327) <= 16702624;
srom_1(74328) <= 16759519;
srom_1(74329) <= 16777161;
srom_1(74330) <= 16755466;
srom_1(74331) <= 16694536;
srom_1(74332) <= 16594657;
srom_1(74333) <= 16456296;
srom_1(74334) <= 16280104;
srom_1(74335) <= 16066905;
srom_1(74336) <= 15817700;
srom_1(74337) <= 15533658;
srom_1(74338) <= 15216110;
srom_1(74339) <= 14866546;
srom_1(74340) <= 14486604;
srom_1(74341) <= 14078067;
srom_1(74342) <= 13642849;
srom_1(74343) <= 13182993;
srom_1(74344) <= 12700655;
srom_1(74345) <= 12198095;
srom_1(74346) <= 11677672;
srom_1(74347) <= 11141825;
srom_1(74348) <= 10593068;
srom_1(74349) <= 10033973;
srom_1(74350) <= 9467162;
srom_1(74351) <= 8895293;
srom_1(74352) <= 8321049;
srom_1(74353) <= 7747121;
srom_1(74354) <= 7176201;
srom_1(74355) <= 6610967;
srom_1(74356) <= 6054069;
srom_1(74357) <= 5508118;
srom_1(74358) <= 4975675;
srom_1(74359) <= 4459236;
srom_1(74360) <= 3961223;
srom_1(74361) <= 3483972;
srom_1(74362) <= 3029721;
srom_1(74363) <= 2600599;
srom_1(74364) <= 2198619;
srom_1(74365) <= 1825666;
srom_1(74366) <= 1483489;
srom_1(74367) <= 1173692;
srom_1(74368) <= 897729;
srom_1(74369) <= 656892;
srom_1(74370) <= 452313;
srom_1(74371) <= 284949;
srom_1(74372) <= 155587;
srom_1(74373) <= 64832;
srom_1(74374) <= 13110;
srom_1(74375) <= 663;
srom_1(74376) <= 27550;
srom_1(74377) <= 93646;
srom_1(74378) <= 198639;
srom_1(74379) <= 342038;
srom_1(74380) <= 523169;
srom_1(74381) <= 741185;
srom_1(74382) <= 995062;
srom_1(74383) <= 1283610;
srom_1(74384) <= 1605476;
srom_1(74385) <= 1959150;
srom_1(74386) <= 2342974;
srom_1(74387) <= 2755148;
srom_1(74388) <= 3193739;
srom_1(74389) <= 3656691;
srom_1(74390) <= 4141832;
srom_1(74391) <= 4646888;
srom_1(74392) <= 5169490;
srom_1(74393) <= 5707188;
srom_1(74394) <= 6257460;
srom_1(74395) <= 6817725;
srom_1(74396) <= 7385357;
srom_1(74397) <= 7957694;
srom_1(74398) <= 8532051;
srom_1(74399) <= 9105735;
srom_1(74400) <= 9676057;
srom_1(74401) <= 10240341;
srom_1(74402) <= 10795942;
srom_1(74403) <= 11340254;
srom_1(74404) <= 11870725;
srom_1(74405) <= 12384867;
srom_1(74406) <= 12880269;
srom_1(74407) <= 13354608;
srom_1(74408) <= 13805660;
srom_1(74409) <= 14231310;
srom_1(74410) <= 14629561;
srom_1(74411) <= 14998546;
srom_1(74412) <= 15336534;
srom_1(74413) <= 15641942;
srom_1(74414) <= 15913336;
srom_1(74415) <= 16149444;
srom_1(74416) <= 16349159;
srom_1(74417) <= 16511544;
srom_1(74418) <= 16635838;
srom_1(74419) <= 16721458;
srom_1(74420) <= 16768002;
srom_1(74421) <= 16775252;
srom_1(74422) <= 16743175;
srom_1(74423) <= 16671920;
srom_1(74424) <= 16561821;
srom_1(74425) <= 16413396;
srom_1(74426) <= 16227340;
srom_1(74427) <= 16004525;
srom_1(74428) <= 15745996;
srom_1(74429) <= 15452967;
srom_1(74430) <= 15126810;
srom_1(74431) <= 14769055;
srom_1(74432) <= 14381380;
srom_1(74433) <= 13965603;
srom_1(74434) <= 13523673;
srom_1(74435) <= 13057664;
srom_1(74436) <= 12569759;
srom_1(74437) <= 12062248;
srom_1(74438) <= 11537510;
srom_1(74439) <= 10998005;
srom_1(74440) <= 10446264;
srom_1(74441) <= 9884874;
srom_1(74442) <= 9316468;
srom_1(74443) <= 8743710;
srom_1(74444) <= 8169287;
srom_1(74445) <= 7595893;
srom_1(74446) <= 7026216;
srom_1(74447) <= 6462928;
srom_1(74448) <= 5908670;
srom_1(74449) <= 5366041;
srom_1(74450) <= 4837586;
srom_1(74451) <= 4325783;
srom_1(74452) <= 3833032;
srom_1(74453) <= 3361644;
srom_1(74454) <= 2913828;
srom_1(74455) <= 2491686;
srom_1(74456) <= 2097197;
srom_1(74457) <= 1732210;
srom_1(74458) <= 1398437;
srom_1(74459) <= 1097444;
srom_1(74460) <= 830641;
srom_1(74461) <= 599280;
srom_1(74462) <= 404446;
srom_1(74463) <= 247053;
srom_1(74464) <= 127838;
srom_1(74465) <= 47361;
srom_1(74466) <= 5998;
srom_1(74467) <= 3945;
srom_1(74468) <= 41210;
srom_1(74469) <= 117619;
srom_1(74470) <= 232813;
srom_1(74471) <= 386253;
srom_1(74472) <= 577219;
srom_1(74473) <= 804814;
srom_1(74474) <= 1067973;
srom_1(74475) <= 1365461;
srom_1(74476) <= 1695883;
srom_1(74477) <= 2057689;
srom_1(74478) <= 2449183;
srom_1(74479) <= 2868529;
srom_1(74480) <= 3313761;
srom_1(74481) <= 3782790;
srom_1(74482) <= 4273418;
srom_1(74483) <= 4783343;
srom_1(74484) <= 5310174;
srom_1(74485) <= 5851441;
srom_1(74486) <= 6404606;
srom_1(74487) <= 6967075;
srom_1(74488) <= 7536209;
srom_1(74489) <= 8109341;
srom_1(74490) <= 8683782;
srom_1(74491) <= 9256839;
srom_1(74492) <= 9825825;
srom_1(74493) <= 10388071;
srom_1(74494) <= 10940941;
srom_1(74495) <= 11481842;
srom_1(74496) <= 12008238;
srom_1(74497) <= 12517660;
srom_1(74498) <= 13007720;
srom_1(74499) <= 13476119;
srom_1(74500) <= 13920661;
srom_1(74501) <= 14339261;
srom_1(74502) <= 14729957;
srom_1(74503) <= 15090916;
srom_1(74504) <= 15420445;
srom_1(74505) <= 15717000;
srom_1(74506) <= 15979189;
srom_1(74507) <= 16205783;
srom_1(74508) <= 16395721;
srom_1(74509) <= 16548109;
srom_1(74510) <= 16662236;
srom_1(74511) <= 16737564;
srom_1(74512) <= 16773741;
srom_1(74513) <= 16770598;
srom_1(74514) <= 16728148;
srom_1(74515) <= 16646591;
srom_1(74516) <= 16526310;
srom_1(74517) <= 16367869;
srom_1(74518) <= 16172010;
srom_1(74519) <= 15939651;
srom_1(74520) <= 15671884;
srom_1(74521) <= 15369962;
srom_1(74522) <= 15035303;
srom_1(74523) <= 14669475;
srom_1(74524) <= 14274194;
srom_1(74525) <= 13851313;
srom_1(74526) <= 13402816;
srom_1(74527) <= 12930805;
srom_1(74528) <= 12437495;
srom_1(74529) <= 11925198;
srom_1(74530) <= 11396316;
srom_1(74531) <= 10853331;
srom_1(74532) <= 10298787;
srom_1(74533) <= 9735286;
srom_1(74534) <= 9165470;
srom_1(74535) <= 8592011;
srom_1(74536) <= 8017598;
srom_1(74537) <= 7444925;
srom_1(74538) <= 6876677;
srom_1(74539) <= 6315519;
srom_1(74540) <= 5764083;
srom_1(74541) <= 5224954;
srom_1(74542) <= 4700660;
srom_1(74543) <= 4193660;
srom_1(74544) <= 3706332;
srom_1(74545) <= 3240961;
srom_1(74546) <= 2799728;
srom_1(74547) <= 2384704;
srom_1(74548) <= 1997835;
srom_1(74549) <= 1640933;
srom_1(74550) <= 1315674;
srom_1(74551) <= 1023583;
srom_1(74552) <= 766028;
srom_1(74553) <= 544219;
srom_1(74554) <= 359194;
srom_1(74555) <= 211822;
srom_1(74556) <= 102794;
srom_1(74557) <= 32621;
srom_1(74558) <= 1632;
srom_1(74559) <= 9972;
srom_1(74560) <= 57603;
srom_1(74561) <= 144300;
srom_1(74562) <= 269658;
srom_1(74563) <= 433089;
srom_1(74564) <= 633825;
srom_1(74565) <= 870927;
srom_1(74566) <= 1143281;
srom_1(74567) <= 1449612;
srom_1(74568) <= 1788481;
srom_1(74569) <= 2158301;
srom_1(74570) <= 2557337;
srom_1(74571) <= 2983718;
srom_1(74572) <= 3435444;
srom_1(74573) <= 3910397;
srom_1(74574) <= 4406350;
srom_1(74575) <= 4920977;
srom_1(74576) <= 5451866;
srom_1(74577) <= 5996525;
srom_1(74578) <= 6552402;
srom_1(74579) <= 7116889;
srom_1(74580) <= 7687340;
srom_1(74581) <= 8261080;
srom_1(74582) <= 8835417;
srom_1(74583) <= 9407659;
srom_1(74584) <= 9975123;
srom_1(74585) <= 10535147;
srom_1(74586) <= 11085104;
srom_1(74587) <= 11622418;
srom_1(74588) <= 12144566;
srom_1(74589) <= 12649102;
srom_1(74590) <= 13133659;
srom_1(74591) <= 13595964;
srom_1(74592) <= 14033851;
srom_1(74593) <= 14445265;
srom_1(74594) <= 14828277;
srom_1(74595) <= 15181091;
srom_1(74596) <= 15502053;
srom_1(74597) <= 15789658;
srom_1(74598) <= 16042557;
srom_1(74599) <= 16259563;
srom_1(74600) <= 16439660;
srom_1(74601) <= 16582003;
srom_1(74602) <= 16685925;
srom_1(74603) <= 16750937;
srom_1(74604) <= 16776735;
srom_1(74605) <= 16763199;
srom_1(74606) <= 16710391;
srom_1(74607) <= 16618559;
srom_1(74608) <= 16488135;
srom_1(74609) <= 16319729;
srom_1(74610) <= 16114131;
srom_1(74611) <= 15872306;
srom_1(74612) <= 15595387;
srom_1(74613) <= 15284673;
srom_1(74614) <= 14941620;
srom_1(74615) <= 14567839;
srom_1(74616) <= 14165081;
srom_1(74617) <= 13735235;
srom_1(74618) <= 13280317;
srom_1(74619) <= 12802460;
srom_1(74620) <= 12303905;
srom_1(74621) <= 11786990;
srom_1(74622) <= 11254138;
srom_1(74623) <= 10707849;
srom_1(74624) <= 10150685;
srom_1(74625) <= 9585257;
srom_1(74626) <= 9014218;
srom_1(74627) <= 8440245;
srom_1(74628) <= 7866030;
srom_1(74629) <= 7294266;
srom_1(74630) <= 6727633;
srom_1(74631) <= 6168789;
srom_1(74632) <= 5620355;
srom_1(74633) <= 5084902;
srom_1(74634) <= 4564941;
srom_1(74635) <= 4062911;
srom_1(74636) <= 3581165;
srom_1(74637) <= 3121963;
srom_1(74638) <= 2687458;
srom_1(74639) <= 2279688;
srom_1(74640) <= 1900565;
srom_1(74641) <= 1551866;
srom_1(74642) <= 1235227;
srom_1(74643) <= 952133;
srom_1(74644) <= 703911;
srom_1(74645) <= 491725;
srom_1(74646) <= 316570;
srom_1(74647) <= 179268;
srom_1(74648) <= 80462;
srom_1(74649) <= 20616;
srom_1(74650) <= 11;
srom_1(74651) <= 18742;
srom_1(74652) <= 76723;
srom_1(74653) <= 173680;
srom_1(74654) <= 309161;
srom_1(74655) <= 482529;
srom_1(74656) <= 692971;
srom_1(74657) <= 939500;
srom_1(74658) <= 1220961;
srom_1(74659) <= 1536034;
srom_1(74660) <= 1883240;
srom_1(74661) <= 2260953;
srom_1(74662) <= 2667400;
srom_1(74663) <= 3100676;
srom_1(74664) <= 3558749;
srom_1(74665) <= 4039470;
srom_1(74666) <= 4540587;
srom_1(74667) <= 5059747;
srom_1(74668) <= 5594519;
srom_1(74669) <= 6142392;
srom_1(74670) <= 6700799;
srom_1(74671) <= 7267120;
srom_1(74672) <= 7838701;
srom_1(74673) <= 8412860;
srom_1(74674) <= 8986906;
srom_1(74675) <= 9558146;
srom_1(74676) <= 10123901;
srom_1(74677) <= 10681519;
srom_1(74678) <= 11228385;
srom_1(74679) <= 11761934;
srom_1(74680) <= 12279665;
srom_1(74681) <= 12779149;
srom_1(74682) <= 13258044;
srom_1(74683) <= 13714105;
srom_1(74684) <= 14145192;
srom_1(74685) <= 14549285;
srom_1(74686) <= 14924489;
srom_1(74687) <= 15269043;
srom_1(74688) <= 15581333;
srom_1(74689) <= 15859894;
srom_1(74690) <= 16103419;
srom_1(74691) <= 16310767;
srom_1(74692) <= 16480965;
srom_1(74693) <= 16613215;
srom_1(74694) <= 16706897;
srom_1(74695) <= 16761572;
srom_1(74696) <= 16776983;
srom_1(74697) <= 16753058;
srom_1(74698) <= 16689909;
srom_1(74699) <= 16587833;
srom_1(74700) <= 16447308;
srom_1(74701) <= 16268993;
srom_1(74702) <= 16053723;
srom_1(74703) <= 15802510;
srom_1(74704) <= 15516530;
srom_1(74705) <= 15197125;
srom_1(74706) <= 14845792;
srom_1(74707) <= 14464180;
srom_1(74708) <= 14054077;
srom_1(74709) <= 13617406;
srom_1(74710) <= 13156216;
srom_1(74711) <= 12672669;
srom_1(74712) <= 12169033;
srom_1(74713) <= 11647669;
srom_1(74714) <= 11111022;
srom_1(74715) <= 10561609;
srom_1(74716) <= 10002005;
srom_1(74717) <= 9434836;
srom_1(74718) <= 8862761;
srom_1(74719) <= 8288462;
srom_1(74720) <= 7714633;
srom_1(74721) <= 7143965;
srom_1(74722) <= 6579133;
srom_1(74723) <= 6022786;
srom_1(74724) <= 5477533;
srom_1(74725) <= 4945932;
srom_1(74726) <= 4430474;
srom_1(74727) <= 3933577;
srom_1(74728) <= 3457572;
srom_1(74729) <= 3004690;
srom_1(74730) <= 2577055;
srom_1(74731) <= 2176672;
srom_1(74732) <= 1805419;
srom_1(74733) <= 1465037;
srom_1(74734) <= 1157122;
srom_1(74735) <= 883118;
srom_1(74736) <= 644309;
srom_1(74737) <= 441817;
srom_1(74738) <= 276589;
srom_1(74739) <= 149402;
srom_1(74740) <= 60851;
srom_1(74741) <= 11352;
srom_1(74742) <= 1136;
srom_1(74743) <= 30252;
srom_1(74744) <= 98564;
srom_1(74745) <= 205750;
srom_1(74746) <= 351309;
srom_1(74747) <= 534557;
srom_1(74748) <= 754636;
srom_1(74749) <= 1010513;
srom_1(74750) <= 1300988;
srom_1(74751) <= 1624700;
srom_1(74752) <= 1980129;
srom_1(74753) <= 2365611;
srom_1(74754) <= 2779336;
srom_1(74755) <= 3219365;
srom_1(74756) <= 3683635;
srom_1(74757) <= 4169967;
srom_1(74758) <= 4676083;
srom_1(74759) <= 5199607;
srom_1(74760) <= 5738086;
srom_1(74761) <= 6288994;
srom_1(74762) <= 6849748;
srom_1(74763) <= 7417719;
srom_1(74764) <= 7990242;
srom_1(74765) <= 8564633;
srom_1(74766) <= 9138198;
srom_1(74767) <= 9708249;
srom_1(74768) <= 10272111;
srom_1(74769) <= 10827141;
srom_1(74770) <= 11370736;
srom_1(74771) <= 11900346;
srom_1(74772) <= 12413489;
srom_1(74773) <= 12907758;
srom_1(74774) <= 13380835;
srom_1(74775) <= 13830501;
srom_1(74776) <= 14254649;
srom_1(74777) <= 14651289;
srom_1(74778) <= 15018561;
srom_1(74779) <= 15354742;
srom_1(74780) <= 15658258;
srom_1(74781) <= 15927683;
srom_1(74782) <= 16161755;
srom_1(74783) <= 16359376;
srom_1(74784) <= 16519619;
srom_1(74785) <= 16641733;
srom_1(74786) <= 16725146;
srom_1(74787) <= 16769466;
srom_1(74788) <= 16774484;
srom_1(74789) <= 16740179;
srom_1(74790) <= 16666710;
srom_1(74791) <= 16554422;
srom_1(74792) <= 16403842;
srom_1(74793) <= 16215676;
srom_1(74794) <= 15990806;
srom_1(74795) <= 15730287;
srom_1(74796) <= 15435340;
srom_1(74797) <= 15107348;
srom_1(74798) <= 14747850;
srom_1(74799) <= 14358532;
srom_1(74800) <= 13941218;
srom_1(74801) <= 13497866;
srom_1(74802) <= 13030555;
srom_1(74803) <= 12541476;
srom_1(74804) <= 12032924;
srom_1(74805) <= 11507281;
srom_1(74806) <= 10967014;
srom_1(74807) <= 10414657;
srom_1(74808) <= 9852798;
srom_1(74809) <= 9284073;
srom_1(74810) <= 8711149;
srom_1(74811) <= 8136713;
srom_1(74812) <= 7563457;
srom_1(74813) <= 6994071;
srom_1(74814) <= 6431225;
srom_1(74815) <= 5877557;
srom_1(74816) <= 5335665;
srom_1(74817) <= 4808089;
srom_1(74818) <= 4297303;
srom_1(74819) <= 3805703;
srom_1(74820) <= 3335593;
srom_1(74821) <= 2889179;
srom_1(74822) <= 2468554;
srom_1(74823) <= 2075689;
srom_1(74824) <= 1712428;
srom_1(74825) <= 1380474;
srom_1(74826) <= 1081384;
srom_1(74827) <= 816560;
srom_1(74828) <= 587243;
srom_1(74829) <= 394510;
srom_1(74830) <= 239264;
srom_1(74831) <= 122233;
srom_1(74832) <= 43966;
srom_1(74833) <= 4829;
srom_1(74834) <= 5008;
srom_1(74835) <= 44499;
srom_1(74836) <= 123119;
srom_1(74837) <= 240499;
srom_1(74838) <= 396088;
srom_1(74839) <= 589157;
srom_1(74840) <= 818800;
srom_1(74841) <= 1083940;
srom_1(74842) <= 1383335;
srom_1(74843) <= 1715580;
srom_1(74844) <= 2079116;
srom_1(74845) <= 2472241;
srom_1(74846) <= 2893109;
srom_1(74847) <= 3339747;
srom_1(74848) <= 3810061;
srom_1(74849) <= 4301846;
srom_1(74850) <= 4812794;
srom_1(74851) <= 5340511;
srom_1(74852) <= 5882522;
srom_1(74853) <= 6436284;
srom_1(74854) <= 6999202;
srom_1(74855) <= 7568635;
srom_1(74856) <= 8141913;
srom_1(74857) <= 8716348;
srom_1(74858) <= 9289246;
srom_1(74859) <= 9857920;
srom_1(74860) <= 10419705;
srom_1(74861) <= 10971965;
srom_1(74862) <= 11512110;
srom_1(74863) <= 12037609;
srom_1(74864) <= 12545996;
srom_1(74865) <= 13034888;
srom_1(74866) <= 13501991;
srom_1(74867) <= 13945116;
srom_1(74868) <= 14362185;
srom_1(74869) <= 14751242;
srom_1(74870) <= 15110462;
srom_1(74871) <= 15438161;
srom_1(74872) <= 15732802;
srom_1(74873) <= 15993004;
srom_1(74874) <= 16217546;
srom_1(74875) <= 16405376;
srom_1(74876) <= 16555612;
srom_1(74877) <= 16667550;
srom_1(74878) <= 16740666;
srom_1(74879) <= 16774615;
srom_1(74880) <= 16769240;
srom_1(74881) <= 16724566;
srom_1(74882) <= 16640801;
srom_1(74883) <= 16518338;
srom_1(74884) <= 16357753;
srom_1(74885) <= 16159797;
srom_1(74886) <= 15925400;
srom_1(74887) <= 15655660;
srom_1(74888) <= 15351843;
srom_1(74889) <= 15015372;
srom_1(74890) <= 14647826;
srom_1(74891) <= 14250929;
srom_1(74892) <= 13826541;
srom_1(74893) <= 13376653;
srom_1(74894) <= 12903374;
srom_1(74895) <= 12408924;
srom_1(74896) <= 11895621;
srom_1(74897) <= 11365873;
srom_1(74898) <= 10822163;
srom_1(74899) <= 10267041;
srom_1(74900) <= 9703111;
srom_1(74901) <= 9133017;
srom_1(74902) <= 8559431;
srom_1(74903) <= 7985045;
srom_1(74904) <= 7412551;
srom_1(74905) <= 6844634;
srom_1(74906) <= 6283958;
srom_1(74907) <= 5733151;
srom_1(74908) <= 5194796;
srom_1(74909) <= 4671418;
srom_1(74910) <= 4165471;
srom_1(74911) <= 3679328;
srom_1(74912) <= 3215269;
srom_1(74913) <= 2775469;
srom_1(74914) <= 2361991;
srom_1(74915) <= 1976774;
srom_1(74916) <= 1621624;
srom_1(74917) <= 1298206;
srom_1(74918) <= 1008039;
srom_1(74919) <= 752481;
srom_1(74920) <= 532731;
srom_1(74921) <= 349821;
srom_1(74922) <= 204607;
srom_1(74923) <= 97770;
srom_1(74924) <= 29813;
srom_1(74925) <= 1052;
srom_1(74926) <= 11624;
srom_1(74927) <= 61478;
srom_1(74928) <= 150381;
srom_1(74929) <= 277916;
srom_1(74930) <= 443484;
srom_1(74931) <= 646310;
srom_1(74932) <= 885443;
srom_1(74933) <= 1159760;
srom_1(74934) <= 1467976;
srom_1(74935) <= 1808645;
srom_1(74936) <= 2180169;
srom_1(74937) <= 2580807;
srom_1(74938) <= 3008680;
srom_1(74939) <= 3461782;
srom_1(74940) <= 3937987;
srom_1(74941) <= 4435062;
srom_1(74942) <= 4950677;
srom_1(74943) <= 5482413;
srom_1(74944) <= 6027778;
srom_1(74945) <= 6584213;
srom_1(74946) <= 7149110;
srom_1(74947) <= 7719819;
srom_1(74948) <= 8293665;
srom_1(74949) <= 8867955;
srom_1(74950) <= 9439998;
srom_1(74951) <= 10007110;
srom_1(74952) <= 10566633;
srom_1(74953) <= 11115942;
srom_1(74954) <= 11652462;
srom_1(74955) <= 12173677;
srom_1(74956) <= 12677142;
srom_1(74957) <= 13160496;
srom_1(74958) <= 13621474;
srom_1(74959) <= 14057912;
srom_1(74960) <= 14467766;
srom_1(74961) <= 14849112;
srom_1(74962) <= 15200163;
srom_1(74963) <= 15519272;
srom_1(74964) <= 15804943;
srom_1(74965) <= 16055836;
srom_1(74966) <= 16270774;
srom_1(74967) <= 16448751;
srom_1(74968) <= 16588931;
srom_1(74969) <= 16690656;
srom_1(74970) <= 16753451;
srom_1(74971) <= 16777020;
srom_1(74972) <= 16761253;
srom_1(74973) <= 16706223;
srom_1(74974) <= 16612189;
srom_1(74975) <= 16479593;
srom_1(74976) <= 16309054;
srom_1(74977) <= 16101374;
srom_1(74978) <= 15857527;
srom_1(74979) <= 15578654;
srom_1(74980) <= 15266066;
srom_1(74981) <= 14921226;
srom_1(74982) <= 14545753;
srom_1(74983) <= 14141407;
srom_1(74984) <= 13710084;
srom_1(74985) <= 13253807;
srom_1(74986) <= 12774715;
srom_1(74987) <= 12275055;
srom_1(74988) <= 11757170;
srom_1(74989) <= 11223489;
srom_1(74990) <= 10676514;
srom_1(74991) <= 10118811;
srom_1(74992) <= 9552994;
srom_1(74993) <= 8981716;
srom_1(74994) <= 8407658;
srom_1(74995) <= 7833510;
srom_1(74996) <= 7261965;
srom_1(74997) <= 6695703;
srom_1(74998) <= 6137380;
srom_1(74999) <= 5589614;
srom_1(75000) <= 5054973;
srom_1(75001) <= 4535964;
srom_1(75002) <= 4035022;
srom_1(75003) <= 3554496;
srom_1(75004) <= 3096638;
srom_1(75005) <= 2663596;
srom_1(75006) <= 2257401;
srom_1(75007) <= 1879957;
srom_1(75008) <= 1533034;
srom_1(75009) <= 1218260;
srom_1(75010) <= 937109;
srom_1(75011) <= 690902;
srom_1(75012) <= 480791;
srom_1(75013) <= 307763;
srom_1(75014) <= 172629;
srom_1(75015) <= 76022;
srom_1(75016) <= 18396;
srom_1(75017) <= 21;
srom_1(75018) <= 20982;
srom_1(75019) <= 81183;
srom_1(75020) <= 180339;
srom_1(75021) <= 317987;
srom_1(75022) <= 493481;
srom_1(75023) <= 705998;
srom_1(75024) <= 954542;
srom_1(75025) <= 1237946;
srom_1(75026) <= 1554882;
srom_1(75027) <= 1903864;
srom_1(75028) <= 2283255;
srom_1(75029) <= 2691276;
srom_1(75030) <= 3126013;
srom_1(75031) <= 3585429;
srom_1(75032) <= 4067369;
srom_1(75033) <= 4569572;
srom_1(75034) <= 5089685;
srom_1(75035) <= 5625267;
srom_1(75036) <= 6173807;
srom_1(75037) <= 6732733;
srom_1(75038) <= 7299424;
srom_1(75039) <= 7871223;
srom_1(75040) <= 8445448;
srom_1(75041) <= 9019406;
srom_1(75042) <= 9590406;
srom_1(75043) <= 10155771;
srom_1(75044) <= 10712849;
srom_1(75045) <= 11259027;
srom_1(75046) <= 11791745;
srom_1(75047) <= 12308505;
srom_1(75048) <= 12806883;
srom_1(75049) <= 13284542;
srom_1(75050) <= 13739243;
srom_1(75051) <= 14168852;
srom_1(75052) <= 14571356;
srom_1(75053) <= 14944867;
srom_1(75054) <= 15287633;
srom_1(75055) <= 15598048;
srom_1(75056) <= 15874655;
srom_1(75057) <= 16116157;
srom_1(75058) <= 16321422;
srom_1(75059) <= 16489487;
srom_1(75060) <= 16619565;
srom_1(75061) <= 16711045;
srom_1(75062) <= 16763498;
srom_1(75063) <= 16776678;
srom_1(75064) <= 16750524;
srom_1(75065) <= 16685157;
srom_1(75066) <= 16580886;
srom_1(75067) <= 16438198;
srom_1(75068) <= 16257763;
srom_1(75069) <= 16040426;
srom_1(75070) <= 15787208;
srom_1(75071) <= 15499295;
srom_1(75072) <= 15178037;
srom_1(75073) <= 14824942;
srom_1(75074) <= 14441664;
srom_1(75075) <= 14030001;
srom_1(75076) <= 13591884;
srom_1(75077) <= 13129368;
srom_1(75078) <= 12644620;
srom_1(75079) <= 12139914;
srom_1(75080) <= 11617617;
srom_1(75081) <= 11080178;
srom_1(75082) <= 10530117;
srom_1(75083) <= 9970014;
srom_1(75084) <= 9402495;
srom_1(75085) <= 8830222;
srom_1(75086) <= 8255878;
srom_1(75087) <= 7682156;
srom_1(75088) <= 7111747;
srom_1(75089) <= 6547326;
srom_1(75090) <= 5991539;
srom_1(75091) <= 5446993;
srom_1(75092) <= 4916241;
srom_1(75093) <= 4401772;
srom_1(75094) <= 3905999;
srom_1(75095) <= 3431246;
srom_1(75096) <= 2979740;
srom_1(75097) <= 2553598;
srom_1(75098) <= 2154819;
srom_1(75099) <= 1785271;
srom_1(75100) <= 1446690;
srom_1(75101) <= 1140661;
srom_1(75102) <= 868620;
srom_1(75103) <= 631843;
srom_1(75104) <= 431440;
srom_1(75105) <= 268351;
srom_1(75106) <= 143341;
srom_1(75107) <= 56996;
srom_1(75108) <= 9720;
srom_1(75109) <= 1736;
srom_1(75110) <= 33081;
srom_1(75111) <= 103607;
srom_1(75112) <= 212985;
srom_1(75113) <= 360702;
srom_1(75114) <= 546063;
srom_1(75115) <= 768202;
srom_1(75116) <= 1026075;
srom_1(75117) <= 1318473;
srom_1(75118) <= 1644026;
srom_1(75119) <= 2001206;
srom_1(75120) <= 2388339;
srom_1(75121) <= 2803609;
srom_1(75122) <= 3245069;
srom_1(75123) <= 3710650;
srom_1(75124) <= 4198166;
srom_1(75125) <= 4705333;
srom_1(75126) <= 5229773;
srom_1(75127) <= 5769025;
srom_1(75128) <= 6320561;
srom_1(75129) <= 6881795;
srom_1(75130) <= 7450095;
srom_1(75131) <= 8022796;
srom_1(75132) <= 8597212;
srom_1(75133) <= 9170650;
srom_1(75134) <= 9740421;
srom_1(75135) <= 10303853;
srom_1(75136) <= 10858303;
srom_1(75137) <= 11401172;
srom_1(75138) <= 11929915;
srom_1(75139) <= 12442050;
srom_1(75140) <= 12935178;
srom_1(75141) <= 13406986;
srom_1(75142) <= 13855260;
srom_1(75143) <= 14277900;
srom_1(75144) <= 14672922;
srom_1(75145) <= 15038476;
srom_1(75146) <= 15372845;
srom_1(75147) <= 15674464;
srom_1(75148) <= 15941916;
srom_1(75149) <= 16173948;
srom_1(75150) <= 16369472;
srom_1(75151) <= 16527572;
srom_1(75152) <= 16647504;
srom_1(75153) <= 16728708;
srom_1(75154) <= 16770803;
srom_1(75155) <= 16773590;
srom_1(75156) <= 16737057;
srom_1(75157) <= 16661376;
srom_1(75158) <= 16546900;
srom_1(75159) <= 16394168;
srom_1(75160) <= 16203895;
srom_1(75161) <= 15976973;
srom_1(75162) <= 15714467;
srom_1(75163) <= 15417607;
srom_1(75164) <= 15087786;
srom_1(75165) <= 14726550;
srom_1(75166) <= 14335593;
srom_1(75167) <= 13916749;
srom_1(75168) <= 13471982;
srom_1(75169) <= 13003376;
srom_1(75170) <= 12513131;
srom_1(75171) <= 12003544;
srom_1(75172) <= 11477006;
srom_1(75173) <= 10935985;
srom_1(75174) <= 10383018;
srom_1(75175) <= 9820699;
srom_1(75176) <= 9251665;
srom_1(75177) <= 8678583;
srom_1(75178) <= 8104141;
srom_1(75179) <= 7531034;
srom_1(75180) <= 6961948;
srom_1(75181) <= 6399552;
srom_1(75182) <= 5846483;
srom_1(75183) <= 5305335;
srom_1(75184) <= 4778646;
srom_1(75185) <= 4268885;
srom_1(75186) <= 3778443;
srom_1(75187) <= 3309619;
srom_1(75188) <= 2864613;
srom_1(75189) <= 2445510;
srom_1(75190) <= 2054277;
srom_1(75191) <= 1692748;
srom_1(75192) <= 1362617;
srom_1(75193) <= 1065434;
srom_1(75194) <= 802592;
srom_1(75195) <= 575324;
srom_1(75196) <= 384694;
srom_1(75197) <= 231598;
srom_1(75198) <= 116752;
srom_1(75199) <= 40697;
srom_1(75200) <= 3787;
srom_1(75201) <= 6197;
srom_1(75202) <= 47914;
srom_1(75203) <= 128744;
srom_1(75204) <= 248308;
srom_1(75205) <= 406044;
srom_1(75206) <= 601213;
srom_1(75207) <= 832900;
srom_1(75208) <= 1100018;
srom_1(75209) <= 1401315;
srom_1(75210) <= 1735377;
srom_1(75211) <= 2100639;
srom_1(75212) <= 2495387;
srom_1(75213) <= 2917771;
srom_1(75214) <= 3365809;
srom_1(75215) <= 3837401;
srom_1(75216) <= 4330335;
srom_1(75217) <= 4842300;
srom_1(75218) <= 5370895;
srom_1(75219) <= 5913640;
srom_1(75220) <= 6467992;
srom_1(75221) <= 7031350;
srom_1(75222) <= 7601073;
srom_1(75223) <= 8174488;
srom_1(75224) <= 8748908;
srom_1(75225) <= 9321638;
srom_1(75226) <= 9889993;
srom_1(75227) <= 10451307;
srom_1(75228) <= 11002949;
srom_1(75229) <= 11542331;
srom_1(75230) <= 12066924;
srom_1(75231) <= 12574269;
srom_1(75232) <= 13061985;
srom_1(75233) <= 13527786;
srom_1(75234) <= 13969488;
srom_1(75235) <= 14385019;
srom_1(75236) <= 14772431;
srom_1(75237) <= 15129907;
srom_1(75238) <= 15455771;
srom_1(75239) <= 15748494;
srom_1(75240) <= 16006704;
srom_1(75241) <= 16229191;
srom_1(75242) <= 16414910;
srom_1(75243) <= 16562991;
srom_1(75244) <= 16672740;
srom_1(75245) <= 16743641;
srom_1(75246) <= 16775363;
srom_1(75247) <= 16767757;
srom_1(75248) <= 16720857;
srom_1(75249) <= 16634885;
srom_1(75250) <= 16510244;
srom_1(75251) <= 16347517;
srom_1(75252) <= 16147468;
srom_1(75253) <= 15911035;
srom_1(75254) <= 15639327;
srom_1(75255) <= 15333618;
srom_1(75256) <= 14995341;
srom_1(75257) <= 14626083;
srom_1(75258) <= 14227575;
srom_1(75259) <= 13801687;
srom_1(75260) <= 13350414;
srom_1(75261) <= 12875874;
srom_1(75262) <= 12380292;
srom_1(75263) <= 11865991;
srom_1(75264) <= 11335384;
srom_1(75265) <= 10790958;
srom_1(75266) <= 10235267;
srom_1(75267) <= 9670916;
srom_1(75268) <= 9100552;
srom_1(75269) <= 8526849;
srom_1(75270) <= 7952498;
srom_1(75271) <= 7380192;
srom_1(75272) <= 6812615;
srom_1(75273) <= 6252428;
srom_1(75274) <= 5702259;
srom_1(75275) <= 5164687;
srom_1(75276) <= 4642233;
srom_1(75277) <= 4137346;
srom_1(75278) <= 3652396;
srom_1(75279) <= 3189655;
srom_1(75280) <= 2751294;
srom_1(75281) <= 2339368;
srom_1(75282) <= 1955809;
srom_1(75283) <= 1602416;
srom_1(75284) <= 1280846;
srom_1(75285) <= 992606;
srom_1(75286) <= 739048;
srom_1(75287) <= 521362;
srom_1(75288) <= 340569;
srom_1(75289) <= 197515;
srom_1(75290) <= 92872;
srom_1(75291) <= 27131;
srom_1(75292) <= 599;
srom_1(75293) <= 13402;
srom_1(75294) <= 65479;
srom_1(75295) <= 156586;
srom_1(75296) <= 286295;
srom_1(75297) <= 454000;
srom_1(75298) <= 658912;
srom_1(75299) <= 900072;
srom_1(75300) <= 1176347;
srom_1(75301) <= 1486444;
srom_1(75302) <= 1828907;
srom_1(75303) <= 2202131;
srom_1(75304) <= 2604366;
srom_1(75305) <= 3033724;
srom_1(75306) <= 3488194;
srom_1(75307) <= 3965643;
srom_1(75308) <= 4463833;
srom_1(75309) <= 4980428;
srom_1(75310) <= 5513005;
srom_1(75311) <= 6059066;
srom_1(75312) <= 6616052;
srom_1(75313) <= 7181349;
srom_1(75314) <= 7752308;
srom_1(75315) <= 8326251;
srom_1(75316) <= 8900486;
srom_1(75317) <= 9472321;
srom_1(75318) <= 10039074;
srom_1(75319) <= 10598087;
srom_1(75320) <= 11146739;
srom_1(75321) <= 11682457;
srom_1(75322) <= 12202730;
srom_1(75323) <= 12705116;
srom_1(75324) <= 13187262;
srom_1(75325) <= 13646904;
srom_1(75326) <= 14081889;
srom_1(75327) <= 14490175;
srom_1(75328) <= 14869850;
srom_1(75329) <= 15219131;
srom_1(75330) <= 15536382;
srom_1(75331) <= 15820115;
srom_1(75332) <= 16068999;
srom_1(75333) <= 16281866;
srom_1(75334) <= 16457720;
srom_1(75335) <= 16595735;
srom_1(75336) <= 16695263;
srom_1(75337) <= 16755839;
srom_1(75338) <= 16777178;
srom_1(75339) <= 16759180;
srom_1(75340) <= 16701930;
srom_1(75341) <= 16605695;
srom_1(75342) <= 16470928;
srom_1(75343) <= 16298260;
srom_1(75344) <= 16088501;
srom_1(75345) <= 15842635;
srom_1(75346) <= 15561814;
srom_1(75347) <= 15247355;
srom_1(75348) <= 14900733;
srom_1(75349) <= 14523574;
srom_1(75350) <= 14117646;
srom_1(75351) <= 13684852;
srom_1(75352) <= 13227223;
srom_1(75353) <= 12746903;
srom_1(75354) <= 12246146;
srom_1(75355) <= 11727300;
srom_1(75356) <= 11192797;
srom_1(75357) <= 10645145;
srom_1(75358) <= 10086911;
srom_1(75359) <= 9520713;
srom_1(75360) <= 8949206;
srom_1(75361) <= 8375070;
srom_1(75362) <= 7800998;
srom_1(75363) <= 7229681;
srom_1(75364) <= 6663799;
srom_1(75365) <= 6106005;
srom_1(75366) <= 5558915;
srom_1(75367) <= 5025094;
srom_1(75368) <= 4507046;
srom_1(75369) <= 4007200;
srom_1(75370) <= 3527900;
srom_1(75371) <= 3071393;
srom_1(75372) <= 2639821;
srom_1(75373) <= 2235207;
srom_1(75374) <= 1859448;
srom_1(75375) <= 1514306;
srom_1(75376) <= 1201401;
srom_1(75377) <= 922199;
srom_1(75378) <= 678009;
srom_1(75379) <= 469977;
srom_1(75380) <= 299078;
srom_1(75381) <= 166114;
srom_1(75382) <= 71708;
srom_1(75383) <= 16302;
srom_1(75384) <= 157;
srom_1(75385) <= 23349;
srom_1(75386) <= 85768;
srom_1(75387) <= 187122;
srom_1(75388) <= 326936;
srom_1(75389) <= 504553;
srom_1(75390) <= 719142;
srom_1(75391) <= 969695;
srom_1(75392) <= 1255038;
srom_1(75393) <= 1573833;
srom_1(75394) <= 1924585;
srom_1(75395) <= 2305649;
srom_1(75396) <= 2715237;
srom_1(75397) <= 3151430;
srom_1(75398) <= 3612183;
srom_1(75399) <= 4095333;
srom_1(75400) <= 4598616;
srom_1(75401) <= 5119672;
srom_1(75402) <= 5656056;
srom_1(75403) <= 6205255;
srom_1(75404) <= 6764692;
srom_1(75405) <= 7331744;
srom_1(75406) <= 7903752;
srom_1(75407) <= 8478034;
srom_1(75408) <= 9051897;
srom_1(75409) <= 9622649;
srom_1(75410) <= 10187614;
srom_1(75411) <= 10744143;
srom_1(75412) <= 11289626;
srom_1(75413) <= 11821505;
srom_1(75414) <= 12337287;
srom_1(75415) <= 12834551;
srom_1(75416) <= 13310967;
srom_1(75417) <= 13764300;
srom_1(75418) <= 14192425;
srom_1(75419) <= 14593334;
srom_1(75420) <= 14965147;
srom_1(75421) <= 15306120;
srom_1(75422) <= 15614654;
srom_1(75423) <= 15889303;
srom_1(75424) <= 16128778;
srom_1(75425) <= 16331958;
srom_1(75426) <= 16497888;
srom_1(75427) <= 16625791;
srom_1(75428) <= 16715067;
srom_1(75429) <= 16765297;
srom_1(75430) <= 16776246;
srom_1(75431) <= 16747863;
srom_1(75432) <= 16680280;
srom_1(75433) <= 16573815;
srom_1(75434) <= 16428967;
srom_1(75435) <= 16246414;
srom_1(75436) <= 16027013;
srom_1(75437) <= 15771794;
srom_1(75438) <= 15481952;
srom_1(75439) <= 15158847;
srom_1(75440) <= 14803994;
srom_1(75441) <= 14419057;
srom_1(75442) <= 14005841;
srom_1(75443) <= 13566284;
srom_1(75444) <= 13102447;
srom_1(75445) <= 12616505;
srom_1(75446) <= 12110738;
srom_1(75447) <= 11587515;
srom_1(75448) <= 11049293;
srom_1(75449) <= 10498593;
srom_1(75450) <= 9937999;
srom_1(75451) <= 9370139;
srom_1(75452) <= 8797676;
srom_1(75453) <= 8223295;
srom_1(75454) <= 7649689;
srom_1(75455) <= 7079549;
srom_1(75456) <= 6515547;
srom_1(75457) <= 5960328;
srom_1(75458) <= 5416497;
srom_1(75459) <= 4886602;
srom_1(75460) <= 4373130;
srom_1(75461) <= 3878488;
srom_1(75462) <= 3404995;
srom_1(75463) <= 2954872;
srom_1(75464) <= 2530230;
srom_1(75465) <= 2133059;
srom_1(75466) <= 1765224;
srom_1(75467) <= 1428447;
srom_1(75468) <= 1124309;
srom_1(75469) <= 854236;
srom_1(75470) <= 619494;
srom_1(75471) <= 421184;
srom_1(75472) <= 260236;
srom_1(75473) <= 137405;
srom_1(75474) <= 53266;
srom_1(75475) <= 8215;
srom_1(75476) <= 2462;
srom_1(75477) <= 36035;
srom_1(75478) <= 108776;
srom_1(75479) <= 220344;
srom_1(75480) <= 370215;
srom_1(75481) <= 557688;
srom_1(75482) <= 781882;
srom_1(75483) <= 1041748;
srom_1(75484) <= 1336065;
srom_1(75485) <= 1663453;
srom_1(75486) <= 2022379;
srom_1(75487) <= 2411157;
srom_1(75488) <= 2827966;
srom_1(75489) <= 3270851;
srom_1(75490) <= 3737735;
srom_1(75491) <= 4226428;
srom_1(75492) <= 4734640;
srom_1(75493) <= 5259985;
srom_1(75494) <= 5800002;
srom_1(75495) <= 6352158;
srom_1(75496) <= 6913864;
srom_1(75497) <= 7482485;
srom_1(75498) <= 8055355;
srom_1(75499) <= 8629788;
srom_1(75500) <= 9203090;
srom_1(75501) <= 9772573;
srom_1(75502) <= 10335565;
srom_1(75503) <= 10889428;
srom_1(75504) <= 11431563;
srom_1(75505) <= 11959429;
srom_1(75506) <= 12470551;
srom_1(75507) <= 12962530;
srom_1(75508) <= 13433061;
srom_1(75509) <= 13879937;
srom_1(75510) <= 14301062;
srom_1(75511) <= 14694461;
srom_1(75512) <= 15058290;
srom_1(75513) <= 15390843;
srom_1(75514) <= 15690560;
srom_1(75515) <= 15956035;
srom_1(75516) <= 16186024;
srom_1(75517) <= 16379449;
srom_1(75518) <= 16535401;
srom_1(75519) <= 16653151;
srom_1(75520) <= 16732145;
srom_1(75521) <= 16772013;
srom_1(75522) <= 16772569;
srom_1(75523) <= 16733809;
srom_1(75524) <= 16655916;
srom_1(75525) <= 16539255;
srom_1(75526) <= 16384373;
srom_1(75527) <= 16191995;
srom_1(75528) <= 15963025;
srom_1(75529) <= 15698536;
srom_1(75530) <= 15399768;
srom_1(75531) <= 15068122;
srom_1(75532) <= 14705154;
srom_1(75533) <= 14312565;
srom_1(75534) <= 13892197;
srom_1(75535) <= 13446020;
srom_1(75536) <= 12976128;
srom_1(75537) <= 12484723;
srom_1(75538) <= 11974110;
srom_1(75539) <= 11446684;
srom_1(75540) <= 10904917;
srom_1(75541) <= 10351350;
srom_1(75542) <= 9788579;
srom_1(75543) <= 9219243;
srom_1(75544) <= 8646012;
srom_1(75545) <= 8071575;
srom_1(75546) <= 7498623;
srom_1(75547) <= 6929845;
srom_1(75548) <= 6367908;
srom_1(75549) <= 5815447;
srom_1(75550) <= 5275052;
srom_1(75551) <= 4749257;
srom_1(75552) <= 4240529;
srom_1(75553) <= 3751252;
srom_1(75554) <= 3283722;
srom_1(75555) <= 2840130;
srom_1(75556) <= 2422557;
srom_1(75557) <= 2032960;
srom_1(75558) <= 1673168;
srom_1(75559) <= 1344866;
srom_1(75560) <= 1049595;
srom_1(75561) <= 788740;
srom_1(75562) <= 563522;
srom_1(75563) <= 374999;
srom_1(75564) <= 224055;
srom_1(75565) <= 111397;
srom_1(75566) <= 37553;
srom_1(75567) <= 2871;
srom_1(75568) <= 7512;
srom_1(75569) <= 51455;
srom_1(75570) <= 134494;
srom_1(75571) <= 256239;
srom_1(75572) <= 416120;
srom_1(75573) <= 613386;
srom_1(75574) <= 847114;
srom_1(75575) <= 1116205;
srom_1(75576) <= 1419400;
srom_1(75577) <= 1755275;
srom_1(75578) <= 2122257;
srom_1(75579) <= 2518623;
srom_1(75580) <= 2942516;
srom_1(75581) <= 3391948;
srom_1(75582) <= 3864810;
srom_1(75583) <= 4358886;
srom_1(75584) <= 4871859;
srom_1(75585) <= 5401324;
srom_1(75586) <= 5944796;
srom_1(75587) <= 6499728;
srom_1(75588) <= 7063519;
srom_1(75589) <= 7633522;
srom_1(75590) <= 8207067;
srom_1(75591) <= 8781463;
srom_1(75592) <= 9354017;
srom_1(75593) <= 9922043;
srom_1(75594) <= 10482879;
srom_1(75595) <= 11033894;
srom_1(75596) <= 11572504;
srom_1(75597) <= 12096184;
srom_1(75598) <= 12602478;
srom_1(75599) <= 13089012;
srom_1(75600) <= 13553504;
srom_1(75601) <= 13993775;
srom_1(75602) <= 14407763;
srom_1(75603) <= 14793524;
srom_1(75604) <= 15149250;
srom_1(75605) <= 15473274;
srom_1(75606) <= 15764075;
srom_1(75607) <= 16020290;
srom_1(75608) <= 16240717;
srom_1(75609) <= 16424323;
srom_1(75610) <= 16570247;
srom_1(75611) <= 16677804;
srom_1(75612) <= 16746491;
srom_1(75613) <= 16775984;
srom_1(75614) <= 16766146;
srom_1(75615) <= 16717023;
srom_1(75616) <= 16628846;
srom_1(75617) <= 16502027;
srom_1(75618) <= 16337161;
srom_1(75619) <= 16135022;
srom_1(75620) <= 15896557;
srom_1(75621) <= 15622885;
srom_1(75622) <= 15315288;
srom_1(75623) <= 14975210;
srom_1(75624) <= 14604246;
srom_1(75625) <= 14204134;
srom_1(75626) <= 13776751;
srom_1(75627) <= 13324101;
srom_1(75628) <= 12848307;
srom_1(75629) <= 12351600;
srom_1(75630) <= 11836309;
srom_1(75631) <= 11304851;
srom_1(75632) <= 10759717;
srom_1(75633) <= 10203464;
srom_1(75634) <= 9638701;
srom_1(75635) <= 9068076;
srom_1(75636) <= 8494265;
srom_1(75637) <= 7919958;
srom_1(75638) <= 7347848;
srom_1(75639) <= 6780620;
srom_1(75640) <= 6220931;
srom_1(75641) <= 5671408;
srom_1(75642) <= 5134626;
srom_1(75643) <= 4613104;
srom_1(75644) <= 4109286;
srom_1(75645) <= 3625535;
srom_1(75646) <= 3164120;
srom_1(75647) <= 2727204;
srom_1(75648) <= 2316837;
srom_1(75649) <= 1934942;
srom_1(75650) <= 1583311;
srom_1(75651) <= 1263592;
srom_1(75652) <= 977285;
srom_1(75653) <= 725732;
srom_1(75654) <= 510112;
srom_1(75655) <= 331438;
srom_1(75656) <= 190547;
srom_1(75657) <= 88099;
srom_1(75658) <= 24575;
srom_1(75659) <= 273;
srom_1(75660) <= 15306;
srom_1(75661) <= 69605;
srom_1(75662) <= 162915;
srom_1(75663) <= 294798;
srom_1(75664) <= 464635;
srom_1(75665) <= 671630;
srom_1(75666) <= 914814;
srom_1(75667) <= 1193044;
srom_1(75668) <= 1505017;
srom_1(75669) <= 1849269;
srom_1(75670) <= 2224186;
srom_1(75671) <= 2628011;
srom_1(75672) <= 3058849;
srom_1(75673) <= 3514680;
srom_1(75674) <= 3993366;
srom_1(75675) <= 4492664;
srom_1(75676) <= 5010231;
srom_1(75677) <= 5543640;
srom_1(75678) <= 6090390;
srom_1(75679) <= 6647917;
srom_1(75680) <= 7213607;
srom_1(75681) <= 7784807;
srom_1(75682) <= 8358838;
srom_1(75683) <= 8933009;
srom_1(75684) <= 9504627;
srom_1(75685) <= 10071012;
srom_1(75686) <= 10629507;
srom_1(75687) <= 11177494;
srom_1(75688) <= 11712403;
srom_1(75689) <= 12231726;
srom_1(75690) <= 12733026;
srom_1(75691) <= 13213955;
srom_1(75692) <= 13672255;
srom_1(75693) <= 14105779;
srom_1(75694) <= 14512493;
srom_1(75695) <= 14890490;
srom_1(75696) <= 15237997;
srom_1(75697) <= 15553385;
srom_1(75698) <= 15835175;
srom_1(75699) <= 16082046;
srom_1(75700) <= 16292839;
srom_1(75701) <= 16466567;
srom_1(75702) <= 16602414;
srom_1(75703) <= 16699744;
srom_1(75704) <= 16758101;
srom_1(75705) <= 16777210;
srom_1(75706) <= 16756981;
srom_1(75707) <= 16697511;
srom_1(75708) <= 16599077;
srom_1(75709) <= 16462142;
srom_1(75710) <= 16287347;
srom_1(75711) <= 16075512;
srom_1(75712) <= 15827630;
srom_1(75713) <= 15544865;
srom_1(75714) <= 15228541;
srom_1(75715) <= 14880142;
srom_1(75716) <= 14501303;
srom_1(75717) <= 14093799;
srom_1(75718) <= 13659541;
srom_1(75719) <= 13200566;
srom_1(75720) <= 12719026;
srom_1(75721) <= 12217179;
srom_1(75722) <= 11697379;
srom_1(75723) <= 11162063;
srom_1(75724) <= 10613741;
srom_1(75725) <= 10054985;
srom_1(75726) <= 9488414;
srom_1(75727) <= 8916687;
srom_1(75728) <= 8342482;
srom_1(75729) <= 7768494;
srom_1(75730) <= 7197414;
srom_1(75731) <= 6631920;
srom_1(75732) <= 6074664;
srom_1(75733) <= 5528258;
srom_1(75734) <= 4995266;
srom_1(75735) <= 4478186;
srom_1(75736) <= 3979443;
srom_1(75737) <= 3501377;
srom_1(75738) <= 3046228;
srom_1(75739) <= 2616132;
srom_1(75740) <= 2213105;
srom_1(75741) <= 1839037;
srom_1(75742) <= 1495682;
srom_1(75743) <= 1184650;
srom_1(75744) <= 907400;
srom_1(75745) <= 665232;
srom_1(75746) <= 459282;
srom_1(75747) <= 290515;
srom_1(75748) <= 159723;
srom_1(75749) <= 67519;
srom_1(75750) <= 14335;
srom_1(75751) <= 421;
srom_1(75752) <= 25842;
srom_1(75753) <= 90479;
srom_1(75754) <= 194029;
srom_1(75755) <= 336006;
srom_1(75756) <= 515744;
srom_1(75757) <= 732401;
srom_1(75758) <= 984961;
srom_1(75759) <= 1272238;
srom_1(75760) <= 1592887;
srom_1(75761) <= 1945403;
srom_1(75762) <= 2328134;
srom_1(75763) <= 2739285;
srom_1(75764) <= 3176927;
srom_1(75765) <= 3639008;
srom_1(75766) <= 4123362;
srom_1(75767) <= 4627717;
srom_1(75768) <= 5149708;
srom_1(75769) <= 5686887;
srom_1(75770) <= 6236736;
srom_1(75771) <= 6796676;
srom_1(75772) <= 7364080;
srom_1(75773) <= 7936289;
srom_1(75774) <= 8510619;
srom_1(75775) <= 9084377;
srom_1(75776) <= 9654873;
srom_1(75777) <= 10219430;
srom_1(75778) <= 10775402;
srom_1(75779) <= 11320181;
srom_1(75780) <= 11851214;
srom_1(75781) <= 12366008;
srom_1(75782) <= 12862152;
srom_1(75783) <= 13337317;
srom_1(75784) <= 13789277;
srom_1(75785) <= 14215910;
srom_1(75786) <= 14615218;
srom_1(75787) <= 14985327;
srom_1(75788) <= 15324501;
srom_1(75789) <= 15631151;
srom_1(75790) <= 15903838;
srom_1(75791) <= 16141283;
srom_1(75792) <= 16342374;
srom_1(75793) <= 16506166;
srom_1(75794) <= 16631893;
srom_1(75795) <= 16718963;
srom_1(75796) <= 16766970;
srom_1(75797) <= 16775688;
srom_1(75798) <= 16745076;
srom_1(75799) <= 16675278;
srom_1(75800) <= 16566621;
srom_1(75801) <= 16419614;
srom_1(75802) <= 16234947;
srom_1(75803) <= 16013485;
srom_1(75804) <= 15756269;
srom_1(75805) <= 15464502;
srom_1(75806) <= 15139554;
srom_1(75807) <= 14782949;
srom_1(75808) <= 14396359;
srom_1(75809) <= 13981596;
srom_1(75810) <= 13540605;
srom_1(75811) <= 13075456;
srom_1(75812) <= 12588327;
srom_1(75813) <= 12081505;
srom_1(75814) <= 11557366;
srom_1(75815) <= 11018367;
srom_1(75816) <= 10467037;
srom_1(75817) <= 9905960;
srom_1(75818) <= 9337767;
srom_1(75819) <= 8765124;
srom_1(75820) <= 8190715;
srom_1(75821) <= 7617234;
srom_1(75822) <= 7047370;
srom_1(75823) <= 6483796;
srom_1(75824) <= 5929154;
srom_1(75825) <= 5386045;
srom_1(75826) <= 4857017;
srom_1(75827) <= 4344549;
srom_1(75828) <= 3851045;
srom_1(75829) <= 3378819;
srom_1(75830) <= 2930086;
srom_1(75831) <= 2506950;
srom_1(75832) <= 2111395;
srom_1(75833) <= 1745276;
srom_1(75834) <= 1410309;
srom_1(75835) <= 1108067;
srom_1(75836) <= 839965;
srom_1(75837) <= 607262;
srom_1(75838) <= 411048;
srom_1(75839) <= 252243;
srom_1(75840) <= 131593;
srom_1(75841) <= 49662;
srom_1(75842) <= 6836;
srom_1(75843) <= 3315;
srom_1(75844) <= 39115;
srom_1(75845) <= 114069;
srom_1(75846) <= 227825;
srom_1(75847) <= 379850;
srom_1(75848) <= 569431;
srom_1(75849) <= 795678;
srom_1(75850) <= 1057531;
srom_1(75851) <= 1353763;
srom_1(75852) <= 1682983;
srom_1(75853) <= 2043648;
srom_1(75854) <= 2434066;
srom_1(75855) <= 2852408;
srom_1(75856) <= 3296710;
srom_1(75857) <= 3764891;
srom_1(75858) <= 4254753;
srom_1(75859) <= 4764001;
srom_1(75860) <= 5290245;
srom_1(75861) <= 5831019;
srom_1(75862) <= 6383787;
srom_1(75863) <= 6945955;
srom_1(75864) <= 7514889;
srom_1(75865) <= 8087920;
srom_1(75866) <= 8662360;
srom_1(75867) <= 9235518;
srom_1(75868) <= 9804703;
srom_1(75869) <= 10367248;
srom_1(75870) <= 10920515;
srom_1(75871) <= 11461909;
srom_1(75872) <= 11988890;
srom_1(75873) <= 12498989;
srom_1(75874) <= 12989813;
srom_1(75875) <= 13459060;
srom_1(75876) <= 13904530;
srom_1(75877) <= 14324134;
srom_1(75878) <= 14715905;
srom_1(75879) <= 15078004;
srom_1(75880) <= 15408735;
srom_1(75881) <= 15706545;
srom_1(75882) <= 15970040;
srom_1(75883) <= 16197982;
srom_1(75884) <= 16389304;
srom_1(75885) <= 16543108;
srom_1(75886) <= 16658672;
srom_1(75887) <= 16735455;
srom_1(75888) <= 16773097;
srom_1(75889) <= 16771421;
srom_1(75890) <= 16730436;
srom_1(75891) <= 16650332;
srom_1(75892) <= 16531487;
srom_1(75893) <= 16374456;
srom_1(75894) <= 16179978;
srom_1(75895) <= 15948963;
srom_1(75896) <= 15682495;
srom_1(75897) <= 15381823;
srom_1(75898) <= 15048358;
srom_1(75899) <= 14683662;
srom_1(75900) <= 14289448;
srom_1(75901) <= 13867562;
srom_1(75902) <= 13419983;
srom_1(75903) <= 12948811;
srom_1(75904) <= 12456254;
srom_1(75905) <= 11944622;
srom_1(75906) <= 11416315;
srom_1(75907) <= 10873811;
srom_1(75908) <= 10319652;
srom_1(75909) <= 9756438;
srom_1(75910) <= 9186810;
srom_1(75911) <= 8613438;
srom_1(75912) <= 8039012;
srom_1(75913) <= 7466226;
srom_1(75914) <= 6897765;
srom_1(75915) <= 6336295;
srom_1(75916) <= 5784449;
srom_1(75917) <= 5244815;
srom_1(75918) <= 4719923;
srom_1(75919) <= 4212235;
srom_1(75920) <= 3724132;
srom_1(75921) <= 3257901;
srom_1(75922) <= 2815731;
srom_1(75923) <= 2399693;
srom_1(75924) <= 2011740;
srom_1(75925) <= 1653690;
srom_1(75926) <= 1327222;
srom_1(75927) <= 1033867;
srom_1(75928) <= 775002;
srom_1(75929) <= 551839;
srom_1(75930) <= 365425;
srom_1(75931) <= 216635;
srom_1(75932) <= 106166;
srom_1(75933) <= 34536;
srom_1(75934) <= 2082;
srom_1(75935) <= 8954;
srom_1(75936) <= 55122;
srom_1(75937) <= 140369;
srom_1(75938) <= 264294;
srom_1(75939) <= 426317;
srom_1(75940) <= 625677;
srom_1(75941) <= 861441;
srom_1(75942) <= 1132502;
srom_1(75943) <= 1437590;
srom_1(75944) <= 1775273;
srom_1(75945) <= 2143969;
srom_1(75946) <= 2541948;
srom_1(75947) <= 2967343;
srom_1(75948) <= 3418161;
srom_1(75949) <= 3892287;
srom_1(75950) <= 4387498;
srom_1(75951) <= 4901472;
srom_1(75952) <= 5431797;
srom_1(75953) <= 5975989;
srom_1(75954) <= 6531494;
srom_1(75955) <= 7095707;
srom_1(75956) <= 7665983;
srom_1(75957) <= 8239648;
srom_1(75958) <= 8814012;
srom_1(75959) <= 9386381;
srom_1(75960) <= 9954070;
srom_1(75961) <= 10514419;
srom_1(75962) <= 11064799;
srom_1(75963) <= 11602630;
srom_1(75964) <= 12125388;
srom_1(75965) <= 12630624;
srom_1(75966) <= 13115968;
srom_1(75967) <= 13579143;
srom_1(75968) <= 14017978;
srom_1(75969) <= 14430415;
srom_1(75970) <= 14814520;
srom_1(75971) <= 15168491;
srom_1(75972) <= 15490670;
srom_1(75973) <= 15779544;
srom_1(75974) <= 16033760;
srom_1(75975) <= 16252125;
srom_1(75976) <= 16433615;
srom_1(75977) <= 16577379;
srom_1(75978) <= 16682744;
srom_1(75979) <= 16749214;
srom_1(75980) <= 16776479;
srom_1(75981) <= 16764410;
srom_1(75982) <= 16713064;
srom_1(75983) <= 16622682;
srom_1(75984) <= 16493687;
srom_1(75985) <= 16326685;
srom_1(75986) <= 16122458;
srom_1(75987) <= 15881965;
srom_1(75988) <= 15606333;
srom_1(75989) <= 15296854;
srom_1(75990) <= 14954980;
srom_1(75991) <= 14582315;
srom_1(75992) <= 14180605;
srom_1(75993) <= 13751734;
srom_1(75994) <= 13297713;
srom_1(75995) <= 12820673;
srom_1(75996) <= 12322848;
srom_1(75997) <= 11806575;
srom_1(75998) <= 11274274;
srom_1(75999) <= 10728440;
srom_1(76000) <= 10171635;
srom_1(76001) <= 9606468;
srom_1(76002) <= 9035590;
srom_1(76003) <= 8461679;
srom_1(76004) <= 7887424;
srom_1(76005) <= 7315520;
srom_1(76006) <= 6748648;
srom_1(76007) <= 6189467;
srom_1(76008) <= 5640597;
srom_1(76009) <= 5104615;
srom_1(76010) <= 4584031;
srom_1(76011) <= 4081289;
srom_1(76012) <= 3598746;
srom_1(76013) <= 3138663;
srom_1(76014) <= 2703200;
srom_1(76015) <= 2294397;
srom_1(76016) <= 1914172;
srom_1(76017) <= 1564308;
srom_1(76018) <= 1246446;
srom_1(76019) <= 962075;
srom_1(76020) <= 712530;
srom_1(76021) <= 498981;
srom_1(76022) <= 322429;
srom_1(76023) <= 183702;
srom_1(76024) <= 83451;
srom_1(76025) <= 22145;
srom_1(76026) <= 73;
srom_1(76027) <= 17337;
srom_1(76028) <= 73857;
srom_1(76029) <= 169368;
srom_1(76030) <= 303422;
srom_1(76031) <= 475390;
srom_1(76032) <= 684465;
srom_1(76033) <= 929668;
srom_1(76034) <= 1209849;
srom_1(76035) <= 1523693;
srom_1(76036) <= 1869729;
srom_1(76037) <= 2246335;
srom_1(76038) <= 2651743;
srom_1(76039) <= 3084054;
srom_1(76040) <= 3541240;
srom_1(76041) <= 4021156;
srom_1(76042) <= 4521553;
srom_1(76043) <= 5040084;
srom_1(76044) <= 5574318;
srom_1(76045) <= 6121748;
srom_1(76046) <= 6679809;
srom_1(76047) <= 7245882;
srom_1(76048) <= 7817315;
srom_1(76049) <= 8391426;
srom_1(76050) <= 8965524;
srom_1(76051) <= 9536917;
srom_1(76052) <= 10102925;
srom_1(76053) <= 10660894;
srom_1(76054) <= 11208207;
srom_1(76055) <= 11742298;
srom_1(76056) <= 12260663;
srom_1(76057) <= 12760870;
srom_1(76058) <= 13240575;
srom_1(76059) <= 13697526;
srom_1(76060) <= 14129583;
srom_1(76061) <= 14534718;
srom_1(76062) <= 14911031;
srom_1(76063) <= 15256759;
srom_1(76064) <= 15570280;
srom_1(76065) <= 15850123;
srom_1(76066) <= 16094977;
srom_1(76067) <= 16303693;
srom_1(76068) <= 16475292;
srom_1(76069) <= 16608970;
srom_1(76070) <= 16704100;
srom_1(76071) <= 16760236;
srom_1(76072) <= 16777114;
srom_1(76073) <= 16754656;
srom_1(76074) <= 16692967;
srom_1(76075) <= 16592335;
srom_1(76076) <= 16453233;
srom_1(76077) <= 16276314;
srom_1(76078) <= 16062406;
srom_1(76079) <= 15812514;
srom_1(76080) <= 15527808;
srom_1(76081) <= 15209624;
srom_1(76082) <= 14859453;
srom_1(76083) <= 14478939;
srom_1(76084) <= 14069865;
srom_1(76085) <= 13634150;
srom_1(76086) <= 13173837;
srom_1(76087) <= 12691084;
srom_1(76088) <= 12188155;
srom_1(76089) <= 11667409;
srom_1(76090) <= 11131287;
srom_1(76091) <= 10582304;
srom_1(76092) <= 10023034;
srom_1(76093) <= 9456100;
srom_1(76094) <= 8884159;
srom_1(76095) <= 8309895;
srom_1(76096) <= 7736000;
srom_1(76097) <= 7165166;
srom_1(76098) <= 6600068;
srom_1(76099) <= 6043358;
srom_1(76100) <= 5497645;
srom_1(76101) <= 4965489;
srom_1(76102) <= 4449385;
srom_1(76103) <= 3951754;
srom_1(76104) <= 3474928;
srom_1(76105) <= 3021144;
srom_1(76106) <= 2592531;
srom_1(76107) <= 2191097;
srom_1(76108) <= 1818725;
srom_1(76109) <= 1477161;
srom_1(76110) <= 1168008;
srom_1(76111) <= 892715;
srom_1(76112) <= 652572;
srom_1(76113) <= 448707;
srom_1(76114) <= 282074;
srom_1(76115) <= 153456;
srom_1(76116) <= 63455;
srom_1(76117) <= 12494;
srom_1(76118) <= 811;
srom_1(76119) <= 28461;
srom_1(76120) <= 95315;
srom_1(76121) <= 201059;
srom_1(76122) <= 345197;
srom_1(76123) <= 527054;
srom_1(76124) <= 745776;
srom_1(76125) <= 1000338;
srom_1(76126) <= 1289546;
srom_1(76127) <= 1612044;
srom_1(76128) <= 1966319;
srom_1(76129) <= 2350711;
srom_1(76130) <= 2763417;
srom_1(76131) <= 3202501;
srom_1(76132) <= 3665905;
srom_1(76133) <= 4151455;
srom_1(76134) <= 4656874;
srom_1(76135) <= 5179793;
srom_1(76136) <= 5717759;
srom_1(76137) <= 6268249;
srom_1(76138) <= 6828683;
srom_1(76139) <= 7396432;
srom_1(76140) <= 7968833;
srom_1(76141) <= 8543203;
srom_1(76142) <= 9116848;
srom_1(76143) <= 9687077;
srom_1(76144) <= 10251218;
srom_1(76145) <= 10806625;
srom_1(76146) <= 11350692;
srom_1(76147) <= 11880869;
srom_1(76148) <= 12394670;
srom_1(76149) <= 12889685;
srom_1(76150) <= 13363593;
srom_1(76151) <= 13814172;
srom_1(76152) <= 14239308;
srom_1(76153) <= 14637008;
srom_1(76154) <= 15005407;
srom_1(76155) <= 15342778;
srom_1(76156) <= 15647539;
srom_1(76157) <= 15918259;
srom_1(76158) <= 16153671;
srom_1(76159) <= 16352670;
srom_1(76160) <= 16514322;
srom_1(76161) <= 16637870;
srom_1(76162) <= 16722734;
srom_1(76163) <= 16768517;
srom_1(76164) <= 16775004;
srom_1(76165) <= 16742164;
srom_1(76166) <= 16670151;
srom_1(76167) <= 16559303;
srom_1(76168) <= 16410140;
srom_1(76169) <= 16223361;
srom_1(76170) <= 15999842;
srom_1(76171) <= 15740632;
srom_1(76172) <= 15446946;
srom_1(76173) <= 15120160;
srom_1(76174) <= 14761808;
srom_1(76175) <= 14373570;
srom_1(76176) <= 13957266;
srom_1(76177) <= 13514849;
srom_1(76178) <= 13048393;
srom_1(76179) <= 12560086;
srom_1(76180) <= 12052217;
srom_1(76181) <= 11527169;
srom_1(76182) <= 10987402;
srom_1(76183) <= 10435449;
srom_1(76184) <= 9873898;
srom_1(76185) <= 9305382;
srom_1(76186) <= 8732566;
srom_1(76187) <= 8158138;
srom_1(76188) <= 7584790;
srom_1(76189) <= 7015212;
srom_1(76190) <= 6452074;
srom_1(76191) <= 5898017;
srom_1(76192) <= 5355639;
srom_1(76193) <= 4827484;
srom_1(76194) <= 4316028;
srom_1(76195) <= 3823670;
srom_1(76196) <= 3352719;
srom_1(76197) <= 2905382;
srom_1(76198) <= 2483759;
srom_1(76199) <= 2089825;
srom_1(76200) <= 1725428;
srom_1(76201) <= 1392277;
srom_1(76202) <= 1091935;
srom_1(76203) <= 825809;
srom_1(76204) <= 595147;
srom_1(76205) <= 401032;
srom_1(76206) <= 244373;
srom_1(76207) <= 125906;
srom_1(76208) <= 46185;
srom_1(76209) <= 5584;
srom_1(76210) <= 4294;
srom_1(76211) <= 42322;
srom_1(76212) <= 119488;
srom_1(76213) <= 235430;
srom_1(76214) <= 389606;
srom_1(76215) <= 581291;
srom_1(76216) <= 809588;
srom_1(76217) <= 1073426;
srom_1(76218) <= 1371567;
srom_1(76219) <= 1702613;
srom_1(76220) <= 2065012;
srom_1(76221) <= 2457065;
srom_1(76222) <= 2876933;
srom_1(76223) <= 3322646;
srom_1(76224) <= 3792116;
srom_1(76225) <= 4283141;
srom_1(76226) <= 4793417;
srom_1(76227) <= 5320552;
srom_1(76228) <= 5862075;
srom_1(76229) <= 6415445;
srom_1(76230) <= 6978068;
srom_1(76231) <= 7547306;
srom_1(76232) <= 8120489;
srom_1(76233) <= 8694929;
srom_1(76234) <= 9267932;
srom_1(76235) <= 9836813;
srom_1(76236) <= 10398902;
srom_1(76237) <= 10951564;
srom_1(76238) <= 11492207;
srom_1(76239) <= 12018297;
srom_1(76240) <= 12527366;
srom_1(76241) <= 13017026;
srom_1(76242) <= 13484983;
srom_1(76243) <= 13929041;
srom_1(76244) <= 14347118;
srom_1(76245) <= 14737253;
srom_1(76246) <= 15097617;
srom_1(76247) <= 15426521;
srom_1(76248) <= 15722421;
srom_1(76249) <= 15983930;
srom_1(76250) <= 16209823;
srom_1(76251) <= 16399039;
srom_1(76252) <= 16550691;
srom_1(76253) <= 16664069;
srom_1(76254) <= 16738640;
srom_1(76255) <= 16774055;
srom_1(76256) <= 16770147;
srom_1(76257) <= 16726936;
srom_1(76258) <= 16644623;
srom_1(76259) <= 16523596;
srom_1(76260) <= 16364420;
srom_1(76261) <= 16167843;
srom_1(76262) <= 15934786;
srom_1(76263) <= 15666343;
srom_1(76264) <= 15363772;
srom_1(76265) <= 15028493;
srom_1(76266) <= 14662076;
srom_1(76267) <= 14266241;
srom_1(76268) <= 13842844;
srom_1(76269) <= 13393870;
srom_1(76270) <= 12921424;
srom_1(76271) <= 12427723;
srom_1(76272) <= 11915081;
srom_1(76273) <= 11385902;
srom_1(76274) <= 10842667;
srom_1(76275) <= 10287925;
srom_1(76276) <= 9724276;
srom_1(76277) <= 9154364;
srom_1(76278) <= 8580860;
srom_1(76279) <= 8006456;
srom_1(76280) <= 7433843;
srom_1(76281) <= 6865707;
srom_1(76282) <= 6304713;
srom_1(76283) <= 5753491;
srom_1(76284) <= 5214626;
srom_1(76285) <= 4690645;
srom_1(76286) <= 4184005;
srom_1(76287) <= 3697082;
srom_1(76288) <= 3232158;
srom_1(76289) <= 2791416;
srom_1(76290) <= 2376920;
srom_1(76291) <= 1990615;
srom_1(76292) <= 1634313;
srom_1(76293) <= 1309684;
srom_1(76294) <= 1018250;
srom_1(76295) <= 761378;
srom_1(76296) <= 540273;
srom_1(76297) <= 355972;
srom_1(76298) <= 209339;
srom_1(76299) <= 101060;
srom_1(76300) <= 31645;
srom_1(76301) <= 1419;
srom_1(76302) <= 10523;
srom_1(76303) <= 58915;
srom_1(76304) <= 146367;
srom_1(76305) <= 272471;
srom_1(76306) <= 436633;
srom_1(76307) <= 638085;
srom_1(76308) <= 875882;
srom_1(76309) <= 1148909;
srom_1(76310) <= 1455885;
srom_1(76311) <= 1795371;
srom_1(76312) <= 2165775;
srom_1(76313) <= 2565360;
srom_1(76314) <= 2992252;
srom_1(76315) <= 3444450;
srom_1(76316) <= 3919832;
srom_1(76317) <= 4416170;
srom_1(76318) <= 4931137;
srom_1(76319) <= 5462316;
srom_1(76320) <= 6007218;
srom_1(76321) <= 6563287;
srom_1(76322) <= 7127915;
srom_1(76323) <= 7698456;
srom_1(76324) <= 8272232;
srom_1(76325) <= 8846555;
srom_1(76326) <= 9418730;
srom_1(76327) <= 9986074;
srom_1(76328) <= 10545927;
srom_1(76329) <= 11095664;
srom_1(76330) <= 11632706;
srom_1(76331) <= 12154536;
srom_1(76332) <= 12658706;
srom_1(76333) <= 13142852;
srom_1(76334) <= 13604704;
srom_1(76335) <= 14042096;
srom_1(76336) <= 14452976;
srom_1(76337) <= 14835419;
srom_1(76338) <= 15187630;
srom_1(76339) <= 15507959;
srom_1(76340) <= 15794902;
srom_1(76341) <= 16047115;
srom_1(76342) <= 16263414;
srom_1(76343) <= 16442786;
srom_1(76344) <= 16584388;
srom_1(76345) <= 16687558;
srom_1(76346) <= 16751811;
srom_1(76347) <= 16776847;
srom_1(76348) <= 16762547;
srom_1(76349) <= 16708979;
srom_1(76350) <= 16616393;
srom_1(76351) <= 16485225;
srom_1(76352) <= 16316089;
srom_1(76353) <= 16109778;
srom_1(76354) <= 15867260;
srom_1(76355) <= 15589672;
srom_1(76356) <= 15278316;
srom_1(76357) <= 14934651;
srom_1(76358) <= 14560290;
srom_1(76359) <= 14156988;
srom_1(76360) <= 13726636;
srom_1(76361) <= 13271252;
srom_1(76362) <= 12792971;
srom_1(76363) <= 12294037;
srom_1(76364) <= 11776789;
srom_1(76365) <= 11243653;
srom_1(76366) <= 10697128;
srom_1(76367) <= 10139778;
srom_1(76368) <= 9574216;
srom_1(76369) <= 9003095;
srom_1(76370) <= 8429092;
srom_1(76371) <= 7854899;
srom_1(76372) <= 7283208;
srom_1(76373) <= 6716702;
srom_1(76374) <= 6158035;
srom_1(76375) <= 5609829;
srom_1(76376) <= 5074653;
srom_1(76377) <= 4555017;
srom_1(76378) <= 4053358;
srom_1(76379) <= 3572029;
srom_1(76380) <= 3113286;
srom_1(76381) <= 2679281;
srom_1(76382) <= 2272050;
srom_1(76383) <= 1893500;
srom_1(76384) <= 1545409;
srom_1(76385) <= 1229408;
srom_1(76386) <= 946978;
srom_1(76387) <= 699445;
srom_1(76388) <= 487969;
srom_1(76389) <= 313542;
srom_1(76390) <= 176982;
srom_1(76391) <= 78928;
srom_1(76392) <= 19842;
srom_1(76393) <= 0;
srom_1(76394) <= 19495;
srom_1(76395) <= 78235;
srom_1(76396) <= 175946;
srom_1(76397) <= 312168;
srom_1(76398) <= 486264;
srom_1(76399) <= 697417;
srom_1(76400) <= 944636;
srom_1(76401) <= 1226762;
srom_1(76402) <= 1542473;
srom_1(76403) <= 1890288;
srom_1(76404) <= 2268576;
srom_1(76405) <= 2675562;
srom_1(76406) <= 3109339;
srom_1(76407) <= 3567872;
srom_1(76408) <= 4049012;
srom_1(76409) <= 4550501;
srom_1(76410) <= 5069988;
srom_1(76411) <= 5605038;
srom_1(76412) <= 6153140;
srom_1(76413) <= 6711726;
srom_1(76414) <= 7278175;
srom_1(76415) <= 7849831;
srom_1(76416) <= 8424014;
srom_1(76417) <= 8998030;
srom_1(76418) <= 9569189;
srom_1(76419) <= 10134812;
srom_1(76420) <= 10692246;
srom_1(76421) <= 11238878;
srom_1(76422) <= 11772143;
srom_1(76423) <= 12289542;
srom_1(76424) <= 12788649;
srom_1(76425) <= 13267122;
srom_1(76426) <= 13722718;
srom_1(76427) <= 14153300;
srom_1(76428) <= 14556850;
srom_1(76429) <= 14931475;
srom_1(76430) <= 15275418;
srom_1(76431) <= 15587066;
srom_1(76432) <= 15864959;
srom_1(76433) <= 16107792;
srom_1(76434) <= 16314427;
srom_1(76435) <= 16483895;
srom_1(76436) <= 16615402;
srom_1(76437) <= 16708331;
srom_1(76438) <= 16762245;
srom_1(76439) <= 16776893;
srom_1(76440) <= 16752205;
srom_1(76441) <= 16688297;
srom_1(76442) <= 16585469;
srom_1(76443) <= 16444204;
srom_1(76444) <= 16265162;
srom_1(76445) <= 16049185;
srom_1(76446) <= 15797285;
srom_1(76447) <= 15510643;
srom_1(76448) <= 15190603;
srom_1(76449) <= 14838667;
srom_1(76450) <= 14456484;
srom_1(76451) <= 14045846;
srom_1(76452) <= 13608680;
srom_1(76453) <= 13147035;
srom_1(76454) <= 12663076;
srom_1(76455) <= 12159073;
srom_1(76456) <= 11637389;
srom_1(76457) <= 11100470;
srom_1(76458) <= 10550834;
srom_1(76459) <= 9991058;
srom_1(76460) <= 9423769;
srom_1(76461) <= 8851625;
srom_1(76462) <= 8277310;
srom_1(76463) <= 7703516;
srom_1(76464) <= 7132936;
srom_1(76465) <= 6568243;
srom_1(76466) <= 6012087;
srom_1(76467) <= 5467075;
srom_1(76468) <= 4935764;
srom_1(76469) <= 4420644;
srom_1(76470) <= 3924131;
srom_1(76471) <= 3448553;
srom_1(76472) <= 2996141;
srom_1(76473) <= 2569016;
srom_1(76474) <= 2169182;
srom_1(76475) <= 1798512;
srom_1(76476) <= 1458745;
srom_1(76477) <= 1151475;
srom_1(76478) <= 878143;
srom_1(76479) <= 640029;
srom_1(76480) <= 438252;
srom_1(76481) <= 273756;
srom_1(76482) <= 147313;
srom_1(76483) <= 59517;
srom_1(76484) <= 10779;
srom_1(76485) <= 1327;
srom_1(76486) <= 31206;
srom_1(76487) <= 100276;
srom_1(76488) <= 208213;
srom_1(76489) <= 354510;
srom_1(76490) <= 538482;
srom_1(76491) <= 759266;
srom_1(76492) <= 1015826;
srom_1(76493) <= 1306960;
srom_1(76494) <= 1631303;
srom_1(76495) <= 1987332;
srom_1(76496) <= 2373380;
srom_1(76497) <= 2787634;
srom_1(76498) <= 3228154;
srom_1(76499) <= 3692873;
srom_1(76500) <= 4179612;
srom_1(76501) <= 4686088;
srom_1(76502) <= 5209926;
srom_1(76503) <= 5748671;
srom_1(76504) <= 6299795;
srom_1(76505) <= 6860714;
srom_1(76506) <= 7428798;
srom_1(76507) <= 8001383;
srom_1(76508) <= 8575784;
srom_1(76509) <= 9149307;
srom_1(76510) <= 9719263;
srom_1(76511) <= 10282978;
srom_1(76512) <= 10837811;
srom_1(76513) <= 11381158;
srom_1(76514) <= 11910473;
srom_1(76515) <= 12423272;
srom_1(76516) <= 12917151;
srom_1(76517) <= 13389794;
srom_1(76518) <= 13838985;
srom_1(76519) <= 14262617;
srom_1(76520) <= 14658704;
srom_1(76521) <= 15025388;
srom_1(76522) <= 15360950;
srom_1(76523) <= 15663817;
srom_1(76524) <= 15932567;
srom_1(76525) <= 16165942;
srom_1(76526) <= 16362845;
srom_1(76527) <= 16522355;
srom_1(76528) <= 16643723;
srom_1(76529) <= 16726379;
srom_1(76530) <= 16769937;
srom_1(76531) <= 16774192;
srom_1(76532) <= 16739125;
srom_1(76533) <= 16664898;
srom_1(76534) <= 16551862;
srom_1(76535) <= 16400545;
srom_1(76536) <= 16211657;
srom_1(76537) <= 15986084;
srom_1(76538) <= 15724885;
srom_1(76539) <= 15429282;
srom_1(76540) <= 15100664;
srom_1(76541) <= 14740571;
srom_1(76542) <= 14350691;
srom_1(76543) <= 13932852;
srom_1(76544) <= 13489015;
srom_1(76545) <= 13021261;
srom_1(76546) <= 12531782;
srom_1(76547) <= 12022874;
srom_1(76548) <= 11496924;
srom_1(76549) <= 10956398;
srom_1(76550) <= 10403831;
srom_1(76551) <= 9841814;
srom_1(76552) <= 9272982;
srom_1(76553) <= 8700003;
srom_1(76554) <= 8125564;
srom_1(76555) <= 7552358;
srom_1(76556) <= 6983074;
srom_1(76557) <= 6420381;
srom_1(76558) <= 5866917;
srom_1(76559) <= 5325279;
srom_1(76560) <= 4798005;
srom_1(76561) <= 4287569;
srom_1(76562) <= 3796365;
srom_1(76563) <= 3326695;
srom_1(76564) <= 2880762;
srom_1(76565) <= 2460657;
srom_1(76566) <= 2068350;
srom_1(76567) <= 1705681;
srom_1(76568) <= 1374351;
srom_1(76569) <= 1075913;
srom_1(76570) <= 811766;
srom_1(76571) <= 583150;
srom_1(76572) <= 391137;
srom_1(76573) <= 236626;
srom_1(76574) <= 120343;
srom_1(76575) <= 42833;
srom_1(76576) <= 4458;
srom_1(76577) <= 5400;
srom_1(76578) <= 45654;
srom_1(76579) <= 125031;
srom_1(76580) <= 243158;
srom_1(76581) <= 399482;
srom_1(76582) <= 593270;
srom_1(76583) <= 823613;
srom_1(76584) <= 1089431;
srom_1(76585) <= 1389477;
srom_1(76586) <= 1722344;
srom_1(76587) <= 2086472;
srom_1(76588) <= 2480153;
srom_1(76589) <= 2901540;
srom_1(76590) <= 3348659;
srom_1(76591) <= 3819411;
srom_1(76592) <= 4311590;
srom_1(76593) <= 4822887;
srom_1(76594) <= 5350905;
srom_1(76595) <= 5893168;
srom_1(76596) <= 6447133;
srom_1(76597) <= 7010203;
srom_1(76598) <= 7579736;
srom_1(76599) <= 8153062;
srom_1(76600) <= 8727493;
srom_1(76601) <= 9300334;
srom_1(76602) <= 9868900;
srom_1(76603) <= 10430525;
srom_1(76604) <= 10982574;
srom_1(76605) <= 11522459;
srom_1(76606) <= 12047649;
srom_1(76607) <= 12555680;
srom_1(76608) <= 13044170;
srom_1(76609) <= 13510829;
srom_1(76610) <= 13953467;
srom_1(76611) <= 14370011;
srom_1(76612) <= 14758505;
srom_1(76613) <= 15117129;
srom_1(76614) <= 15444200;
srom_1(76615) <= 15738186;
srom_1(76616) <= 15997706;
srom_1(76617) <= 16221545;
srom_1(76618) <= 16408653;
srom_1(76619) <= 16558151;
srom_1(76620) <= 16669340;
srom_1(76621) <= 16741698;
srom_1(76622) <= 16774886;
srom_1(76623) <= 16768747;
srom_1(76624) <= 16723311;
srom_1(76625) <= 16638790;
srom_1(76626) <= 16515582;
srom_1(76627) <= 16354263;
srom_1(76628) <= 16155591;
srom_1(76629) <= 15920496;
srom_1(76630) <= 15650082;
srom_1(76631) <= 15345617;
srom_1(76632) <= 15008527;
srom_1(76633) <= 14640395;
srom_1(76634) <= 14242946;
srom_1(76635) <= 13818043;
srom_1(76636) <= 13367681;
srom_1(76637) <= 12893969;
srom_1(76638) <= 12399131;
srom_1(76639) <= 11885486;
srom_1(76640) <= 11355442;
srom_1(76641) <= 10811487;
srom_1(76642) <= 10256169;
srom_1(76643) <= 9692094;
srom_1(76644) <= 9121906;
srom_1(76645) <= 8548280;
srom_1(76646) <= 7973905;
srom_1(76647) <= 7401474;
srom_1(76648) <= 6833673;
srom_1(76649) <= 6273163;
srom_1(76650) <= 5722573;
srom_1(76651) <= 5184485;
srom_1(76652) <= 4661423;
srom_1(76653) <= 4155838;
srom_1(76654) <= 3670102;
srom_1(76655) <= 3206493;
srom_1(76656) <= 2767185;
srom_1(76657) <= 2354238;
srom_1(76658) <= 1969587;
srom_1(76659) <= 1615038;
srom_1(76660) <= 1292252;
srom_1(76661) <= 1002744;
srom_1(76662) <= 747870;
srom_1(76663) <= 528827;
srom_1(76664) <= 346640;
srom_1(76665) <= 202166;
srom_1(76666) <= 96080;
srom_1(76667) <= 28880;
srom_1(76668) <= 883;
srom_1(76669) <= 12218;
srom_1(76670) <= 62833;
srom_1(76671) <= 152491;
srom_1(76672) <= 280770;
srom_1(76673) <= 447070;
srom_1(76674) <= 650610;
srom_1(76675) <= 890437;
srom_1(76676) <= 1165425;
srom_1(76677) <= 1474285;
srom_1(76678) <= 1815569;
srom_1(76679) <= 2187676;
srom_1(76680) <= 2588861;
srom_1(76681) <= 3017243;
srom_1(76682) <= 3470813;
srom_1(76683) <= 3947445;
srom_1(76684) <= 4444903;
srom_1(76685) <= 4960854;
srom_1(76686) <= 5492879;
srom_1(76687) <= 6038483;
srom_1(76688) <= 6595107;
srom_1(76689) <= 7160142;
srom_1(76690) <= 7730938;
srom_1(76691) <= 8304818;
srom_1(76692) <= 8879090;
srom_1(76693) <= 9451063;
srom_1(76694) <= 10018053;
srom_1(76695) <= 10577402;
srom_1(76696) <= 11126488;
srom_1(76697) <= 11662734;
srom_1(76698) <= 12183627;
srom_1(76699) <= 12686724;
srom_1(76700) <= 13169665;
srom_1(76701) <= 13630186;
srom_1(76702) <= 14066128;
srom_1(76703) <= 14475446;
srom_1(76704) <= 14856221;
srom_1(76705) <= 15206667;
srom_1(76706) <= 15525140;
srom_1(76707) <= 15810148;
srom_1(76708) <= 16060354;
srom_1(76709) <= 16274584;
srom_1(76710) <= 16451834;
srom_1(76711) <= 16591273;
srom_1(76712) <= 16692247;
srom_1(76713) <= 16754283;
srom_1(76714) <= 16777088;
srom_1(76715) <= 16760557;
srom_1(76716) <= 16704768;
srom_1(76717) <= 16609981;
srom_1(76718) <= 16476641;
srom_1(76719) <= 16305373;
srom_1(76720) <= 16096981;
srom_1(76721) <= 15852442;
srom_1(76722) <= 15572903;
srom_1(76723) <= 15259673;
srom_1(76724) <= 14914223;
srom_1(76725) <= 14538172;
srom_1(76726) <= 14133284;
srom_1(76727) <= 13701457;
srom_1(76728) <= 13244716;
srom_1(76729) <= 12765203;
srom_1(76730) <= 12265167;
srom_1(76731) <= 11746952;
srom_1(76732) <= 11212989;
srom_1(76733) <= 10665781;
srom_1(76734) <= 10107895;
srom_1(76735) <= 9541947;
srom_1(76736) <= 8970590;
srom_1(76737) <= 8396504;
srom_1(76738) <= 7822381;
srom_1(76739) <= 7250913;
srom_1(76740) <= 6684780;
srom_1(76741) <= 6126637;
srom_1(76742) <= 5579102;
srom_1(76743) <= 5044741;
srom_1(76744) <= 4526060;
srom_1(76745) <= 4025492;
srom_1(76746) <= 3545385;
srom_1(76747) <= 3087989;
srom_1(76748) <= 2655449;
srom_1(76749) <= 2249794;
srom_1(76750) <= 1872926;
srom_1(76751) <= 1526613;
srom_1(76752) <= 1212477;
srom_1(76753) <= 931993;
srom_1(76754) <= 686476;
srom_1(76755) <= 477076;
srom_1(76756) <= 304777;
srom_1(76757) <= 170385;
srom_1(76758) <= 74531;
srom_1(76759) <= 17665;
srom_1(76760) <= 53;
srom_1(76761) <= 21778;
srom_1(76762) <= 82738;
srom_1(76763) <= 182647;
srom_1(76764) <= 321036;
srom_1(76765) <= 497258;
srom_1(76766) <= 710484;
srom_1(76767) <= 959716;
srom_1(76768) <= 1243784;
srom_1(76769) <= 1561357;
srom_1(76770) <= 1910945;
srom_1(76771) <= 2290909;
srom_1(76772) <= 2699467;
srom_1(76773) <= 3134704;
srom_1(76774) <= 3594578;
srom_1(76775) <= 4076933;
srom_1(76776) <= 4579507;
srom_1(76777) <= 5099943;
srom_1(76778) <= 5635800;
srom_1(76779) <= 6184567;
srom_1(76780) <= 6743669;
srom_1(76781) <= 7310484;
srom_1(76782) <= 7882356;
srom_1(76783) <= 8456601;
srom_1(76784) <= 9030527;
srom_1(76785) <= 9601444;
srom_1(76786) <= 10166673;
srom_1(76787) <= 10723564;
srom_1(76788) <= 11269505;
srom_1(76789) <= 11801937;
srom_1(76790) <= 12318363;
srom_1(76791) <= 12816361;
srom_1(76792) <= 13293595;
srom_1(76793) <= 13747828;
srom_1(76794) <= 14176930;
srom_1(76795) <= 14578889;
srom_1(76796) <= 14951819;
srom_1(76797) <= 15293972;
srom_1(76798) <= 15603744;
srom_1(76799) <= 15879681;
srom_1(76800) <= 16120490;
srom_1(76801) <= 16325042;
srom_1(76802) <= 16492376;
srom_1(76803) <= 16621710;
srom_1(76804) <= 16712436;
srom_1(76805) <= 16764128;
srom_1(76806) <= 16776545;
srom_1(76807) <= 16749627;
srom_1(76808) <= 16683502;
srom_1(76809) <= 16578480;
srom_1(76810) <= 16435052;
srom_1(76811) <= 16253892;
srom_1(76812) <= 16035848;
srom_1(76813) <= 15781945;
srom_1(76814) <= 15493371;
srom_1(76815) <= 15171480;
srom_1(76816) <= 14817783;
srom_1(76817) <= 14433937;
srom_1(76818) <= 14021742;
srom_1(76819) <= 13583131;
srom_1(76820) <= 13120162;
srom_1(76821) <= 12635004;
srom_1(76822) <= 12129934;
srom_1(76823) <= 11607319;
srom_1(76824) <= 11069611;
srom_1(76825) <= 10519331;
srom_1(76826) <= 9959059;
srom_1(76827) <= 9391422;
srom_1(76828) <= 8819083;
srom_1(76829) <= 8244726;
srom_1(76830) <= 7671043;
srom_1(76831) <= 7100725;
srom_1(76832) <= 6536446;
srom_1(76833) <= 5980853;
srom_1(76834) <= 5436550;
srom_1(76835) <= 4906091;
srom_1(76836) <= 4391962;
srom_1(76837) <= 3896575;
srom_1(76838) <= 3422253;
srom_1(76839) <= 2971219;
srom_1(76840) <= 2545590;
srom_1(76841) <= 2147361;
srom_1(76842) <= 1778398;
srom_1(76843) <= 1440434;
srom_1(76844) <= 1135052;
srom_1(76845) <= 863684;
srom_1(76846) <= 627603;
srom_1(76847) <= 427916;
srom_1(76848) <= 265560;
srom_1(76849) <= 141295;
srom_1(76850) <= 55705;
srom_1(76851) <= 9191;
srom_1(76852) <= 1970;
srom_1(76853) <= 34078;
srom_1(76854) <= 105362;
srom_1(76855) <= 215490;
srom_1(76856) <= 363944;
srom_1(76857) <= 550029;
srom_1(76858) <= 772871;
srom_1(76859) <= 1031426;
srom_1(76860) <= 1324482;
srom_1(76861) <= 1650664;
srom_1(76862) <= 2008442;
srom_1(76863) <= 2396139;
srom_1(76864) <= 2811936;
srom_1(76865) <= 3253885;
srom_1(76866) <= 3719912;
srom_1(76867) <= 4207832;
srom_1(76868) <= 4715358;
srom_1(76869) <= 5240108;
srom_1(76870) <= 5779623;
srom_1(76871) <= 6331372;
srom_1(76872) <= 6892768;
srom_1(76873) <= 7461179;
srom_1(76874) <= 8033939;
srom_1(76875) <= 8608362;
srom_1(76876) <= 9181755;
srom_1(76877) <= 9751428;
srom_1(76878) <= 10314710;
srom_1(76879) <= 10868960;
srom_1(76880) <= 11411579;
srom_1(76881) <= 11940023;
srom_1(76882) <= 12451812;
srom_1(76883) <= 12944548;
srom_1(76884) <= 13415919;
srom_1(76885) <= 13863716;
srom_1(76886) <= 14285837;
srom_1(76887) <= 14680305;
srom_1(76888) <= 15045269;
srom_1(76889) <= 15379017;
srom_1(76890) <= 15679985;
srom_1(76891) <= 15946761;
srom_1(76892) <= 16178095;
srom_1(76893) <= 16372900;
srom_1(76894) <= 16530265;
srom_1(76895) <= 16649451;
srom_1(76896) <= 16729899;
srom_1(76897) <= 16771231;
srom_1(76898) <= 16773255;
srom_1(76899) <= 16735960;
srom_1(76900) <= 16659521;
srom_1(76901) <= 16544297;
srom_1(76902) <= 16390829;
srom_1(76903) <= 16199835;
srom_1(76904) <= 15972212;
srom_1(76905) <= 15709026;
srom_1(76906) <= 15411513;
srom_1(76907) <= 15081067;
srom_1(76908) <= 14719237;
srom_1(76909) <= 14327722;
srom_1(76910) <= 13908355;
srom_1(76911) <= 13463105;
srom_1(76912) <= 12994058;
srom_1(76913) <= 12503415;
srom_1(76914) <= 11993476;
srom_1(76915) <= 11466633;
srom_1(76916) <= 10925356;
srom_1(76917) <= 10372183;
srom_1(76918) <= 9809708;
srom_1(76919) <= 9240569;
srom_1(76920) <= 8667436;
srom_1(76921) <= 8092994;
srom_1(76922) <= 7519939;
srom_1(76923) <= 6950958;
srom_1(76924) <= 6388718;
srom_1(76925) <= 5835856;
srom_1(76926) <= 5294965;
srom_1(76927) <= 4768581;
srom_1(76928) <= 4259173;
srom_1(76929) <= 3769128;
srom_1(76930) <= 3300747;
srom_1(76931) <= 2856224;
srom_1(76932) <= 2437644;
srom_1(76933) <= 2046970;
srom_1(76934) <= 1686035;
srom_1(76935) <= 1356530;
srom_1(76936) <= 1060001;
srom_1(76937) <= 797838;
srom_1(76938) <= 571271;
srom_1(76939) <= 381362;
srom_1(76940) <= 229002;
srom_1(76941) <= 114905;
srom_1(76942) <= 39607;
srom_1(76943) <= 3459;
srom_1(76944) <= 6633;
srom_1(76945) <= 49112;
srom_1(76946) <= 130698;
srom_1(76947) <= 251009;
srom_1(76948) <= 409479;
srom_1(76949) <= 605366;
srom_1(76950) <= 837752;
srom_1(76951) <= 1105546;
srom_1(76952) <= 1407493;
srom_1(76953) <= 1742176;
srom_1(76954) <= 2108027;
srom_1(76955) <= 2503330;
srom_1(76956) <= 2926231;
srom_1(76957) <= 3374747;
srom_1(76958) <= 3846775;
srom_1(76959) <= 4340101;
srom_1(76960) <= 4852411;
srom_1(76961) <= 5381304;
srom_1(76962) <= 5924300;
srom_1(76963) <= 6478851;
srom_1(76964) <= 7042358;
srom_1(76965) <= 7612178;
srom_1(76966) <= 8185639;
srom_1(76967) <= 8760051;
srom_1(76968) <= 9332722;
srom_1(76969) <= 9900965;
srom_1(76970) <= 10462117;
srom_1(76971) <= 11013545;
srom_1(76972) <= 11552664;
srom_1(76973) <= 12076945;
srom_1(76974) <= 12583931;
srom_1(76975) <= 13071243;
srom_1(76976) <= 13536597;
srom_1(76977) <= 13977810;
srom_1(76978) <= 14392814;
srom_1(76979) <= 14779661;
srom_1(76980) <= 15136539;
srom_1(76981) <= 15461773;
srom_1(76982) <= 15753839;
srom_1(76983) <= 16011367;
srom_1(76984) <= 16233149;
srom_1(76985) <= 16418145;
srom_1(76986) <= 16565489;
srom_1(76987) <= 16674487;
srom_1(76988) <= 16744631;
srom_1(76989) <= 16775590;
srom_1(76990) <= 16767220;
srom_1(76991) <= 16719559;
srom_1(76992) <= 16632832;
srom_1(76993) <= 16507445;
srom_1(76994) <= 16343986;
srom_1(76995) <= 16143221;
srom_1(76996) <= 15906092;
srom_1(76997) <= 15633712;
srom_1(76998) <= 15327356;
srom_1(76999) <= 14988462;
srom_1(77000) <= 14618620;
srom_1(77001) <= 14219562;
srom_1(77002) <= 13793161;
srom_1(77003) <= 13341417;
srom_1(77004) <= 12866447;
srom_1(77005) <= 12370479;
srom_1(77006) <= 11855838;
srom_1(77007) <= 11324938;
srom_1(77008) <= 10780269;
srom_1(77009) <= 10224385;
srom_1(77010) <= 9659892;
srom_1(77011) <= 9089438;
srom_1(77012) <= 8515697;
srom_1(77013) <= 7941360;
srom_1(77014) <= 7369120;
srom_1(77015) <= 6801661;
srom_1(77016) <= 6241644;
srom_1(77017) <= 5691695;
srom_1(77018) <= 5154392;
srom_1(77019) <= 4632256;
srom_1(77020) <= 4127735;
srom_1(77021) <= 3643194;
srom_1(77022) <= 3180906;
srom_1(77023) <= 2743039;
srom_1(77024) <= 2331646;
srom_1(77025) <= 1948656;
srom_1(77026) <= 1595865;
srom_1(77027) <= 1274928;
srom_1(77028) <= 987349;
srom_1(77029) <= 734478;
srom_1(77030) <= 517499;
srom_1(77031) <= 337430;
srom_1(77032) <= 195116;
srom_1(77033) <= 91224;
srom_1(77034) <= 26242;
srom_1(77035) <= 473;
srom_1(77036) <= 14040;
srom_1(77037) <= 66877;
srom_1(77038) <= 158738;
srom_1(77039) <= 289192;
srom_1(77040) <= 457626;
srom_1(77041) <= 663252;
srom_1(77042) <= 905105;
srom_1(77043) <= 1182050;
srom_1(77044) <= 1492789;
srom_1(77045) <= 1835865;
srom_1(77046) <= 2209669;
srom_1(77047) <= 2612449;
srom_1(77048) <= 3042314;
srom_1(77049) <= 3497251;
srom_1(77050) <= 3975124;
srom_1(77051) <= 4473694;
srom_1(77052) <= 4990623;
srom_1(77053) <= 5523485;
srom_1(77054) <= 6069783;
srom_1(77055) <= 6626955;
srom_1(77056) <= 7192388;
srom_1(77057) <= 7763430;
srom_1(77058) <= 8337404;
srom_1(77059) <= 8911619;
srom_1(77060) <= 9483380;
srom_1(77061) <= 10050008;
srom_1(77062) <= 10608845;
srom_1(77063) <= 11157270;
srom_1(77064) <= 11692712;
srom_1(77065) <= 12212661;
srom_1(77066) <= 12714676;
srom_1(77067) <= 13196406;
srom_1(77068) <= 13655590;
srom_1(77069) <= 14090075;
srom_1(77070) <= 14497824;
srom_1(77071) <= 14876925;
srom_1(77072) <= 15225600;
srom_1(77073) <= 15542214;
srom_1(77074) <= 15825282;
srom_1(77075) <= 16073477;
srom_1(77076) <= 16285635;
srom_1(77077) <= 16460762;
srom_1(77078) <= 16598035;
srom_1(77079) <= 16696811;
srom_1(77080) <= 16756627;
srom_1(77081) <= 16777203;
srom_1(77082) <= 16758442;
srom_1(77083) <= 16700431;
srom_1(77084) <= 16603444;
srom_1(77085) <= 16467935;
srom_1(77086) <= 16294538;
srom_1(77087) <= 16084068;
srom_1(77088) <= 15837512;
srom_1(77089) <= 15556025;
srom_1(77090) <= 15240927;
srom_1(77091) <= 14893697;
srom_1(77092) <= 14515962;
srom_1(77093) <= 14109494;
srom_1(77094) <= 13676198;
srom_1(77095) <= 13218107;
srom_1(77096) <= 12737369;
srom_1(77097) <= 12236238;
srom_1(77098) <= 11717065;
srom_1(77099) <= 11182283;
srom_1(77100) <= 10634400;
srom_1(77101) <= 10075986;
srom_1(77102) <= 9509660;
srom_1(77103) <= 8938076;
srom_1(77104) <= 8363916;
srom_1(77105) <= 7789872;
srom_1(77106) <= 7218635;
srom_1(77107) <= 6652885;
srom_1(77108) <= 6095274;
srom_1(77109) <= 5548417;
srom_1(77110) <= 5014879;
srom_1(77111) <= 4497162;
srom_1(77112) <= 3997692;
srom_1(77113) <= 3518814;
srom_1(77114) <= 3062771;
srom_1(77115) <= 2631703;
srom_1(77116) <= 2227631;
srom_1(77117) <= 1852451;
srom_1(77118) <= 1507920;
srom_1(77119) <= 1195655;
srom_1(77120) <= 917121;
srom_1(77121) <= 673623;
srom_1(77122) <= 466303;
srom_1(77123) <= 296133;
srom_1(77124) <= 163912;
srom_1(77125) <= 70260;
srom_1(77126) <= 15615;
srom_1(77127) <= 233;
srom_1(77128) <= 24188;
srom_1(77129) <= 87366;
srom_1(77130) <= 189472;
srom_1(77131) <= 330026;
srom_1(77132) <= 508370;
srom_1(77133) <= 723667;
srom_1(77134) <= 974907;
srom_1(77135) <= 1260913;
srom_1(77136) <= 1580343;
srom_1(77137) <= 1931699;
srom_1(77138) <= 2313334;
srom_1(77139) <= 2723458;
srom_1(77140) <= 3160148;
srom_1(77141) <= 3621356;
srom_1(77142) <= 4104919;
srom_1(77143) <= 4608570;
srom_1(77144) <= 5129946;
srom_1(77145) <= 5666604;
srom_1(77146) <= 6216026;
srom_1(77147) <= 6775636;
srom_1(77148) <= 7342810;
srom_1(77149) <= 7914888;
srom_1(77150) <= 8489187;
srom_1(77151) <= 9063015;
srom_1(77152) <= 9633680;
srom_1(77153) <= 10198507;
srom_1(77154) <= 10754846;
srom_1(77155) <= 11300089;
srom_1(77156) <= 11831679;
srom_1(77157) <= 12347124;
srom_1(77158) <= 12844006;
srom_1(77159) <= 13319994;
srom_1(77160) <= 13772858;
srom_1(77161) <= 14200473;
srom_1(77162) <= 14600835;
srom_1(77163) <= 14972065;
srom_1(77164) <= 15312423;
srom_1(77165) <= 15620313;
srom_1(77166) <= 15894290;
srom_1(77167) <= 16133072;
srom_1(77168) <= 16335536;
srom_1(77169) <= 16500735;
srom_1(77170) <= 16627893;
srom_1(77171) <= 16716415;
srom_1(77172) <= 16765884;
srom_1(77173) <= 16776070;
srom_1(77174) <= 16746924;
srom_1(77175) <= 16678582;
srom_1(77176) <= 16571367;
srom_1(77177) <= 16425779;
srom_1(77178) <= 16242502;
srom_1(77179) <= 16022396;
srom_1(77180) <= 15766493;
srom_1(77181) <= 15475991;
srom_1(77182) <= 15152255;
srom_1(77183) <= 14796802;
srom_1(77184) <= 14411298;
srom_1(77185) <= 13997552;
srom_1(77186) <= 13557504;
srom_1(77187) <= 13093217;
srom_1(77188) <= 12606868;
srom_1(77189) <= 12100739;
srom_1(77190) <= 11577202;
srom_1(77191) <= 11038712;
srom_1(77192) <= 10487796;
srom_1(77193) <= 9927035;
srom_1(77194) <= 9359061;
srom_1(77195) <= 8786535;
srom_1(77196) <= 8212144;
srom_1(77197) <= 7638580;
srom_1(77198) <= 7068533;
srom_1(77199) <= 6504676;
srom_1(77200) <= 5949654;
srom_1(77201) <= 5406069;
srom_1(77202) <= 4876470;
srom_1(77203) <= 4363341;
srom_1(77204) <= 3869087;
srom_1(77205) <= 3396027;
srom_1(77206) <= 2946379;
srom_1(77207) <= 2522252;
srom_1(77208) <= 2125634;
srom_1(77209) <= 1758385;
srom_1(77210) <= 1422227;
srom_1(77211) <= 1118737;
srom_1(77212) <= 849339;
srom_1(77213) <= 615294;
srom_1(77214) <= 417701;
srom_1(77215) <= 257486;
srom_1(77216) <= 135401;
srom_1(77217) <= 52018;
srom_1(77218) <= 7729;
srom_1(77219) <= 2740;
srom_1(77220) <= 37075;
srom_1(77221) <= 110574;
srom_1(77222) <= 222891;
srom_1(77223) <= 373499;
srom_1(77224) <= 561694;
srom_1(77225) <= 786591;
srom_1(77226) <= 1047137;
srom_1(77227) <= 1342110;
srom_1(77228) <= 1670126;
srom_1(77229) <= 2029647;
srom_1(77230) <= 2418988;
srom_1(77231) <= 2836322;
srom_1(77232) <= 3279693;
srom_1(77233) <= 3747022;
srom_1(77234) <= 4236116;
srom_1(77235) <= 4744683;
srom_1(77236) <= 5270337;
srom_1(77237) <= 5810614;
srom_1(77238) <= 6362980;
srom_1(77239) <= 6924845;
srom_1(77240) <= 7493574;
srom_1(77241) <= 8066500;
srom_1(77242) <= 8640937;
srom_1(77243) <= 9214190;
srom_1(77244) <= 9783572;
srom_1(77245) <= 10346413;
srom_1(77246) <= 10900072;
srom_1(77247) <= 11441955;
srom_1(77248) <= 11969519;
srom_1(77249) <= 12480291;
srom_1(77250) <= 12971876;
srom_1(77251) <= 13441968;
srom_1(77252) <= 13888364;
srom_1(77253) <= 14308969;
srom_1(77254) <= 14701811;
srom_1(77255) <= 15065049;
srom_1(77256) <= 15396979;
srom_1(77257) <= 15696043;
srom_1(77258) <= 15960841;
srom_1(77259) <= 16190130;
srom_1(77260) <= 16382835;
srom_1(77261) <= 16538053;
srom_1(77262) <= 16655054;
srom_1(77263) <= 16733292;
srom_1(77264) <= 16772398;
srom_1(77265) <= 16772190;
srom_1(77266) <= 16732669;
srom_1(77267) <= 16654019;
srom_1(77268) <= 16536610;
srom_1(77269) <= 16380992;
srom_1(77270) <= 16187895;
srom_1(77271) <= 15958225;
srom_1(77272) <= 15693058;
srom_1(77273) <= 15393638;
srom_1(77274) <= 15061369;
srom_1(77275) <= 14697809;
srom_1(77276) <= 14304663;
srom_1(77277) <= 13883774;
srom_1(77278) <= 13437117;
srom_1(77279) <= 12966786;
srom_1(77280) <= 12474986;
srom_1(77281) <= 11964024;
srom_1(77282) <= 11436295;
srom_1(77283) <= 10894274;
srom_1(77284) <= 10340504;
srom_1(77285) <= 9777581;
srom_1(77286) <= 9208144;
srom_1(77287) <= 8634864;
srom_1(77288) <= 8060429;
srom_1(77289) <= 7487533;
srom_1(77290) <= 6918863;
srom_1(77291) <= 6357085;
srom_1(77292) <= 5804833;
srom_1(77293) <= 5264697;
srom_1(77294) <= 4739211;
srom_1(77295) <= 4230838;
srom_1(77296) <= 3741962;
srom_1(77297) <= 3274876;
srom_1(77298) <= 2831769;
srom_1(77299) <= 2414721;
srom_1(77300) <= 2025686;
srom_1(77301) <= 1666490;
srom_1(77302) <= 1338815;
srom_1(77303) <= 1044200;
srom_1(77304) <= 784025;
srom_1(77305) <= 559510;
srom_1(77306) <= 371709;
srom_1(77307) <= 221501;
srom_1(77308) <= 109592;
srom_1(77309) <= 36507;
srom_1(77310) <= 2587;
srom_1(77311) <= 7992;
srom_1(77312) <= 52696;
srom_1(77313) <= 136491;
srom_1(77314) <= 258982;
srom_1(77315) <= 419596;
srom_1(77316) <= 617580;
srom_1(77317) <= 852005;
srom_1(77318) <= 1121771;
srom_1(77319) <= 1425614;
srom_1(77320) <= 1762109;
srom_1(77321) <= 2129677;
srom_1(77322) <= 2526596;
srom_1(77323) <= 2951004;
srom_1(77324) <= 3400911;
srom_1(77325) <= 3874207;
srom_1(77326) <= 4368672;
srom_1(77327) <= 4881989;
srom_1(77328) <= 5411749;
srom_1(77329) <= 5955468;
srom_1(77330) <= 6510597;
srom_1(77331) <= 7074533;
srom_1(77332) <= 7644631;
srom_1(77333) <= 8218218;
srom_1(77334) <= 8792604;
srom_1(77335) <= 9365095;
srom_1(77336) <= 9933008;
srom_1(77337) <= 10493678;
srom_1(77338) <= 11044476;
srom_1(77339) <= 11582821;
srom_1(77340) <= 12106186;
srom_1(77341) <= 12612119;
srom_1(77342) <= 13098246;
srom_1(77343) <= 13562288;
srom_1(77344) <= 14002069;
srom_1(77345) <= 14415526;
srom_1(77346) <= 14800721;
srom_1(77347) <= 15155847;
srom_1(77348) <= 15479240;
srom_1(77349) <= 15769382;
srom_1(77350) <= 16024913;
srom_1(77351) <= 16244635;
srom_1(77352) <= 16427517;
srom_1(77353) <= 16572702;
srom_1(77354) <= 16679509;
srom_1(77355) <= 16747437;
srom_1(77356) <= 16776168;
srom_1(77357) <= 16765566;
srom_1(77358) <= 16715682;
srom_1(77359) <= 16626750;
srom_1(77360) <= 16499186;
srom_1(77361) <= 16333589;
srom_1(77362) <= 16130735;
srom_1(77363) <= 15891575;
srom_1(77364) <= 15617232;
srom_1(77365) <= 15308991;
srom_1(77366) <= 14968298;
srom_1(77367) <= 14596750;
srom_1(77368) <= 14196090;
srom_1(77369) <= 13768198;
srom_1(77370) <= 13315078;
srom_1(77371) <= 12838856;
srom_1(77372) <= 12341766;
srom_1(77373) <= 11826138;
srom_1(77374) <= 11294390;
srom_1(77375) <= 10749016;
srom_1(77376) <= 10192573;
srom_1(77377) <= 9627671;
srom_1(77378) <= 9056958;
srom_1(77379) <= 8483112;
srom_1(77380) <= 7908822;
srom_1(77381) <= 7336782;
srom_1(77382) <= 6769674;
srom_1(77383) <= 6210158;
srom_1(77384) <= 5660858;
srom_1(77385) <= 5124349;
srom_1(77386) <= 4603147;
srom_1(77387) <= 4099696;
srom_1(77388) <= 3616358;
srom_1(77389) <= 3155398;
srom_1(77390) <= 2718979;
srom_1(77391) <= 2309146;
srom_1(77392) <= 1927822;
srom_1(77393) <= 1576795;
srom_1(77394) <= 1257711;
srom_1(77395) <= 972066;
srom_1(77396) <= 721200;
srom_1(77397) <= 506289;
srom_1(77398) <= 328341;
srom_1(77399) <= 188190;
srom_1(77400) <= 86494;
srom_1(77401) <= 23729;
srom_1(77402) <= 190;
srom_1(77403) <= 15987;
srom_1(77404) <= 71047;
srom_1(77405) <= 165110;
srom_1(77406) <= 297736;
srom_1(77407) <= 468303;
srom_1(77408) <= 676010;
srom_1(77409) <= 919885;
srom_1(77410) <= 1198783;
srom_1(77411) <= 1511397;
srom_1(77412) <= 1856261;
srom_1(77413) <= 2231757;
srom_1(77414) <= 2636124;
srom_1(77415) <= 3067467;
srom_1(77416) <= 3523762;
srom_1(77417) <= 4002870;
srom_1(77418) <= 4502545;
srom_1(77419) <= 5020443;
srom_1(77420) <= 5554135;
srom_1(77421) <= 6101119;
srom_1(77422) <= 6658830;
srom_1(77423) <= 7224652;
srom_1(77424) <= 7795932;
srom_1(77425) <= 8369992;
srom_1(77426) <= 8944139;
srom_1(77427) <= 9515681;
srom_1(77428) <= 10081938;
srom_1(77429) <= 10640254;
srom_1(77430) <= 11188011;
srom_1(77431) <= 11722641;
srom_1(77432) <= 12241636;
srom_1(77433) <= 12742564;
srom_1(77434) <= 13223074;
srom_1(77435) <= 13680914;
srom_1(77436) <= 14113936;
srom_1(77437) <= 14520110;
srom_1(77438) <= 14897531;
srom_1(77439) <= 15244430;
srom_1(77440) <= 15559180;
srom_1(77441) <= 15840304;
srom_1(77442) <= 16086485;
srom_1(77443) <= 16296568;
srom_1(77444) <= 16469567;
srom_1(77445) <= 16604672;
srom_1(77446) <= 16701249;
srom_1(77447) <= 16758846;
srom_1(77448) <= 16777191;
srom_1(77449) <= 16756200;
srom_1(77450) <= 16695970;
srom_1(77451) <= 16596784;
srom_1(77452) <= 16459106;
srom_1(77453) <= 16283584;
srom_1(77454) <= 16071039;
srom_1(77455) <= 15822469;
srom_1(77456) <= 15539039;
srom_1(77457) <= 15222078;
srom_1(77458) <= 14873072;
srom_1(77459) <= 14493659;
srom_1(77460) <= 14085617;
srom_1(77461) <= 13650859;
srom_1(77462) <= 13191426;
srom_1(77463) <= 12709470;
srom_1(77464) <= 12207252;
srom_1(77465) <= 11687127;
srom_1(77466) <= 11151534;
srom_1(77467) <= 10602985;
srom_1(77468) <= 10044052;
srom_1(77469) <= 9477356;
srom_1(77470) <= 8905554;
srom_1(77471) <= 8331329;
srom_1(77472) <= 7757372;
srom_1(77473) <= 7186375;
srom_1(77474) <= 6621015;
srom_1(77475) <= 6063945;
srom_1(77476) <= 5517775;
srom_1(77477) <= 4985068;
srom_1(77478) <= 4468322;
srom_1(77479) <= 3969959;
srom_1(77480) <= 3492316;
srom_1(77481) <= 3037634;
srom_1(77482) <= 2608044;
srom_1(77483) <= 2205562;
srom_1(77484) <= 1832074;
srom_1(77485) <= 1489331;
srom_1(77486) <= 1178942;
srom_1(77487) <= 902361;
srom_1(77488) <= 660886;
srom_1(77489) <= 455649;
srom_1(77490) <= 287612;
srom_1(77491) <= 157564;
srom_1(77492) <= 66114;
srom_1(77493) <= 13690;
srom_1(77494) <= 540;
srom_1(77495) <= 26724;
srom_1(77496) <= 92120;
srom_1(77497) <= 196421;
srom_1(77498) <= 339138;
srom_1(77499) <= 519602;
srom_1(77500) <= 736966;
srom_1(77501) <= 990211;
srom_1(77502) <= 1278150;
srom_1(77503) <= 1599432;
srom_1(77504) <= 1952551;
srom_1(77505) <= 2335851;
srom_1(77506) <= 2747535;
srom_1(77507) <= 3185671;
srom_1(77508) <= 3648206;
srom_1(77509) <= 4132970;
srom_1(77510) <= 4637690;
srom_1(77511) <= 5159999;
srom_1(77512) <= 5697449;
srom_1(77513) <= 6247518;
srom_1(77514) <= 6807628;
srom_1(77515) <= 7375151;
srom_1(77516) <= 7947427;
srom_1(77517) <= 8521772;
srom_1(77518) <= 9095492;
srom_1(77519) <= 9665897;
srom_1(77520) <= 10230313;
srom_1(77521) <= 10786092;
srom_1(77522) <= 11330629;
srom_1(77523) <= 11861370;
srom_1(77524) <= 12375825;
srom_1(77525) <= 12871583;
srom_1(77526) <= 13346319;
srom_1(77527) <= 13797807;
srom_1(77528) <= 14223929;
srom_1(77529) <= 14622687;
srom_1(77530) <= 14992211;
srom_1(77531) <= 15330769;
srom_1(77532) <= 15636772;
srom_1(77533) <= 15908787;
srom_1(77534) <= 16145536;
srom_1(77535) <= 16345911;
srom_1(77536) <= 16508971;
srom_1(77537) <= 16633952;
srom_1(77538) <= 16720268;
srom_1(77539) <= 16767514;
srom_1(77540) <= 16775468;
srom_1(77541) <= 16744094;
srom_1(77542) <= 16673537;
srom_1(77543) <= 16564130;
srom_1(77544) <= 16416385;
srom_1(77545) <= 16230995;
srom_1(77546) <= 16008829;
srom_1(77547) <= 15750929;
srom_1(77548) <= 15458505;
srom_1(77549) <= 15132928;
srom_1(77550) <= 14775724;
srom_1(77551) <= 14388569;
srom_1(77552) <= 13973278;
srom_1(77553) <= 13531799;
srom_1(77554) <= 13066201;
srom_1(77555) <= 12578668;
srom_1(77556) <= 12071487;
srom_1(77557) <= 11547036;
srom_1(77558) <= 11007774;
srom_1(77559) <= 10456229;
srom_1(77560) <= 9894989;
srom_1(77561) <= 9326684;
srom_1(77562) <= 8753981;
srom_1(77563) <= 8179565;
srom_1(77564) <= 7606128;
srom_1(77565) <= 7036361;
srom_1(77566) <= 6472935;
srom_1(77567) <= 5918493;
srom_1(77568) <= 5375633;
srom_1(77569) <= 4846903;
srom_1(77570) <= 4334780;
srom_1(77571) <= 3841668;
srom_1(77572) <= 3369877;
srom_1(77573) <= 2921622;
srom_1(77574) <= 2499002;
srom_1(77575) <= 2104001;
srom_1(77576) <= 1738471;
srom_1(77577) <= 1404126;
srom_1(77578) <= 1102533;
srom_1(77579) <= 835107;
srom_1(77580) <= 603102;
srom_1(77581) <= 407606;
srom_1(77582) <= 249536;
srom_1(77583) <= 129632;
srom_1(77584) <= 48458;
srom_1(77585) <= 6393;
srom_1(77586) <= 3636;
srom_1(77587) <= 40199;
srom_1(77588) <= 115910;
srom_1(77589) <= 230414;
srom_1(77590) <= 383176;
srom_1(77591) <= 573477;
srom_1(77592) <= 800426;
srom_1(77593) <= 1062959;
srom_1(77594) <= 1359844;
srom_1(77595) <= 1689690;
srom_1(77596) <= 2050949;
srom_1(77597) <= 2441928;
srom_1(77598) <= 2860792;
srom_1(77599) <= 3305579;
srom_1(77600) <= 3774201;
srom_1(77601) <= 4264462;
srom_1(77602) <= 4774063;
srom_1(77603) <= 5300613;
srom_1(77604) <= 5841644;
srom_1(77605) <= 6394619;
srom_1(77606) <= 6956944;
srom_1(77607) <= 7525983;
srom_1(77608) <= 8099066;
srom_1(77609) <= 8673508;
srom_1(77610) <= 9246614;
srom_1(77611) <= 9815696;
srom_1(77612) <= 10378086;
srom_1(77613) <= 10931146;
srom_1(77614) <= 11472284;
srom_1(77615) <= 11998961;
srom_1(77616) <= 12508709;
srom_1(77617) <= 12999135;
srom_1(77618) <= 13467941;
srom_1(77619) <= 13912929;
srom_1(77620) <= 14332011;
srom_1(77621) <= 14723222;
srom_1(77622) <= 15084728;
srom_1(77623) <= 15414834;
srom_1(77624) <= 15711992;
srom_1(77625) <= 15974807;
srom_1(77626) <= 16202048;
srom_1(77627) <= 16392650;
srom_1(77628) <= 16545717;
srom_1(77629) <= 16660533;
srom_1(77630) <= 16736559;
srom_1(77631) <= 16773439;
srom_1(77632) <= 16771000;
srom_1(77633) <= 16729252;
srom_1(77634) <= 16648392;
srom_1(77635) <= 16528800;
srom_1(77636) <= 16371035;
srom_1(77637) <= 16175838;
srom_1(77638) <= 15944124;
srom_1(77639) <= 15676979;
srom_1(77640) <= 15375657;
srom_1(77641) <= 15041570;
srom_1(77642) <= 14676285;
srom_1(77643) <= 14281515;
srom_1(77644) <= 13859111;
srom_1(77645) <= 13411054;
srom_1(77646) <= 12939445;
srom_1(77647) <= 12446495;
srom_1(77648) <= 11934517;
srom_1(77649) <= 11405911;
srom_1(77650) <= 10863155;
srom_1(77651) <= 10308796;
srom_1(77652) <= 9745432;
srom_1(77653) <= 9175706;
srom_1(77654) <= 8602288;
srom_1(77655) <= 8027869;
srom_1(77656) <= 7455141;
srom_1(77657) <= 6886790;
srom_1(77658) <= 6325482;
srom_1(77659) <= 5773849;
srom_1(77660) <= 5234477;
srom_1(77661) <= 4709896;
srom_1(77662) <= 4202566;
srom_1(77663) <= 3714865;
srom_1(77664) <= 3249082;
srom_1(77665) <= 2807399;
srom_1(77666) <= 2391889;
srom_1(77667) <= 2004499;
srom_1(77668) <= 1647046;
srom_1(77669) <= 1321207;
srom_1(77670) <= 1028509;
srom_1(77671) <= 770326;
srom_1(77672) <= 547867;
srom_1(77673) <= 362176;
srom_1(77674) <= 214124;
srom_1(77675) <= 104404;
srom_1(77676) <= 33533;
srom_1(77677) <= 1841;
srom_1(77678) <= 9477;
srom_1(77679) <= 56406;
srom_1(77680) <= 142408;
srom_1(77681) <= 267079;
srom_1(77682) <= 429834;
srom_1(77683) <= 629911;
srom_1(77684) <= 866371;
srom_1(77685) <= 1138105;
srom_1(77686) <= 1443840;
srom_1(77687) <= 1782141;
srom_1(77688) <= 2151422;
srom_1(77689) <= 2549951;
srom_1(77690) <= 2975860;
srom_1(77691) <= 3427151;
srom_1(77692) <= 3901708;
srom_1(77693) <= 4397305;
srom_1(77694) <= 4911619;
srom_1(77695) <= 5442238;
srom_1(77696) <= 5986673;
srom_1(77697) <= 6542372;
srom_1(77698) <= 7106729;
srom_1(77699) <= 7677096;
srom_1(77700) <= 8250801;
srom_1(77701) <= 8825151;
srom_1(77702) <= 9397454;
srom_1(77703) <= 9965027;
srom_1(77704) <= 10525207;
srom_1(77705) <= 11075368;
srom_1(77706) <= 11612929;
srom_1(77707) <= 12135371;
srom_1(77708) <= 12640243;
srom_1(77709) <= 13125177;
srom_1(77710) <= 13587901;
srom_1(77711) <= 14026242;
srom_1(77712) <= 14438147;
srom_1(77713) <= 14821684;
srom_1(77714) <= 15175054;
srom_1(77715) <= 15496599;
srom_1(77716) <= 15784813;
srom_1(77717) <= 16038344;
srom_1(77718) <= 16256002;
srom_1(77719) <= 16436767;
srom_1(77720) <= 16579792;
srom_1(77721) <= 16684406;
srom_1(77722) <= 16750117;
srom_1(77723) <= 16776619;
srom_1(77724) <= 16763786;
srom_1(77725) <= 16711680;
srom_1(77726) <= 16620543;
srom_1(77727) <= 16490804;
srom_1(77728) <= 16323072;
srom_1(77729) <= 16118131;
srom_1(77730) <= 15876945;
srom_1(77731) <= 15600643;
srom_1(77732) <= 15290521;
srom_1(77733) <= 14948034;
srom_1(77734) <= 14574787;
srom_1(77735) <= 14172531;
srom_1(77736) <= 13743153;
srom_1(77737) <= 13288665;
srom_1(77738) <= 12811199;
srom_1(77739) <= 12312994;
srom_1(77740) <= 11796386;
srom_1(77741) <= 11263798;
srom_1(77742) <= 10717727;
srom_1(77743) <= 10160734;
srom_1(77744) <= 9595431;
srom_1(77745) <= 9024469;
srom_1(77746) <= 8450525;
srom_1(77747) <= 7876291;
srom_1(77748) <= 7304459;
srom_1(77749) <= 6737711;
srom_1(77750) <= 6178705;
srom_1(77751) <= 5630062;
srom_1(77752) <= 5094354;
srom_1(77753) <= 4574094;
srom_1(77754) <= 4071722;
srom_1(77755) <= 3589593;
srom_1(77756) <= 3129969;
srom_1(77757) <= 2695004;
srom_1(77758) <= 2286738;
srom_1(77759) <= 1907086;
srom_1(77760) <= 1557828;
srom_1(77761) <= 1240602;
srom_1(77762) <= 956895;
srom_1(77763) <= 708039;
srom_1(77764) <= 495199;
srom_1(77765) <= 319374;
srom_1(77766) <= 181388;
srom_1(77767) <= 81889;
srom_1(77768) <= 21343;
srom_1(77769) <= 34;
srom_1(77770) <= 18062;
srom_1(77771) <= 75342;
srom_1(77772) <= 171606;
srom_1(77773) <= 306402;
srom_1(77774) <= 479098;
srom_1(77775) <= 688885;
srom_1(77776) <= 934779;
srom_1(77777) <= 1215626;
srom_1(77778) <= 1530109;
srom_1(77779) <= 1876755;
srom_1(77780) <= 2253937;
srom_1(77781) <= 2659886;
srom_1(77782) <= 3092699;
srom_1(77783) <= 3550347;
srom_1(77784) <= 4030683;
srom_1(77785) <= 4531454;
srom_1(77786) <= 5050314;
srom_1(77787) <= 5584827;
srom_1(77788) <= 6132489;
srom_1(77789) <= 6690730;
srom_1(77790) <= 7256933;
srom_1(77791) <= 7828443;
srom_1(77792) <= 8402580;
srom_1(77793) <= 8976651;
srom_1(77794) <= 9547965;
srom_1(77795) <= 10113842;
srom_1(77796) <= 10671629;
srom_1(77797) <= 11218709;
srom_1(77798) <= 11752519;
srom_1(77799) <= 12270554;
srom_1(77800) <= 12770385;
srom_1(77801) <= 13249669;
srom_1(77802) <= 13706158;
srom_1(77803) <= 14137710;
srom_1(77804) <= 14542303;
srom_1(77805) <= 14918040;
srom_1(77806) <= 15263157;
srom_1(77807) <= 15576037;
srom_1(77808) <= 15855214;
srom_1(77809) <= 16099376;
srom_1(77810) <= 16307380;
srom_1(77811) <= 16478251;
srom_1(77812) <= 16611186;
srom_1(77813) <= 16705562;
srom_1(77814) <= 16760938;
srom_1(77815) <= 16777053;
srom_1(77816) <= 16753831;
srom_1(77817) <= 16691383;
srom_1(77818) <= 16589999;
srom_1(77819) <= 16450157;
srom_1(77820) <= 16272511;
srom_1(77821) <= 16057894;
srom_1(77822) <= 15807314;
srom_1(77823) <= 15521945;
srom_1(77824) <= 15203125;
srom_1(77825) <= 14852350;
srom_1(77826) <= 14471264;
srom_1(77827) <= 14061654;
srom_1(77828) <= 13625441;
srom_1(77829) <= 13164671;
srom_1(77830) <= 12681505;
srom_1(77831) <= 12178207;
srom_1(77832) <= 11657139;
srom_1(77833) <= 11120744;
srom_1(77834) <= 10571537;
srom_1(77835) <= 10012093;
srom_1(77836) <= 9445036;
srom_1(77837) <= 8873025;
srom_1(77838) <= 8298742;
srom_1(77839) <= 7724881;
srom_1(77840) <= 7154132;
srom_1(77841) <= 6589173;
srom_1(77842) <= 6032651;
srom_1(77843) <= 5487177;
srom_1(77844) <= 4955309;
srom_1(77845) <= 4439541;
srom_1(77846) <= 3942292;
srom_1(77847) <= 3465892;
srom_1(77848) <= 3012577;
srom_1(77849) <= 2584473;
srom_1(77850) <= 2183585;
srom_1(77851) <= 1811795;
srom_1(77852) <= 1470846;
srom_1(77853) <= 1162337;
srom_1(77854) <= 887715;
srom_1(77855) <= 648266;
srom_1(77856) <= 445115;
srom_1(77857) <= 279213;
srom_1(77858) <= 151339;
srom_1(77859) <= 62093;
srom_1(77860) <= 11892;
srom_1(77861) <= 973;
srom_1(77862) <= 29386;
srom_1(77863) <= 96999;
srom_1(77864) <= 203494;
srom_1(77865) <= 348371;
srom_1(77866) <= 530952;
srom_1(77867) <= 750380;
srom_1(77868) <= 1005626;
srom_1(77869) <= 1295494;
srom_1(77870) <= 1618624;
srom_1(77871) <= 1973501;
srom_1(77872) <= 2358460;
srom_1(77873) <= 2771696;
srom_1(77874) <= 3211273;
srom_1(77875) <= 3675127;
srom_1(77876) <= 4161085;
srom_1(77877) <= 4666867;
srom_1(77878) <= 5190101;
srom_1(77879) <= 5728335;
srom_1(77880) <= 6279043;
srom_1(77881) <= 6839644;
srom_1(77882) <= 7407508;
srom_1(77883) <= 7979973;
srom_1(77884) <= 8554354;
srom_1(77885) <= 9127959;
srom_1(77886) <= 9698096;
srom_1(77887) <= 10262092;
srom_1(77888) <= 10817303;
srom_1(77889) <= 11361125;
srom_1(77890) <= 11891008;
srom_1(77891) <= 12404466;
srom_1(77892) <= 12899093;
srom_1(77893) <= 13372569;
srom_1(77894) <= 13822674;
srom_1(77895) <= 14247296;
srom_1(77896) <= 14644444;
srom_1(77897) <= 15012257;
srom_1(77898) <= 15349010;
srom_1(77899) <= 15653122;
srom_1(77900) <= 15923169;
srom_1(77901) <= 16157884;
srom_1(77902) <= 16356166;
srom_1(77903) <= 16517085;
srom_1(77904) <= 16639887;
srom_1(77905) <= 16723996;
srom_1(77906) <= 16769017;
srom_1(77907) <= 16774740;
srom_1(77908) <= 16741138;
srom_1(77909) <= 16668367;
srom_1(77910) <= 16556770;
srom_1(77911) <= 16406869;
srom_1(77912) <= 16219368;
srom_1(77913) <= 15995146;
srom_1(77914) <= 15735255;
srom_1(77915) <= 15440912;
srom_1(77916) <= 15113499;
srom_1(77917) <= 14754550;
srom_1(77918) <= 14365749;
srom_1(77919) <= 13948920;
srom_1(77920) <= 13506016;
srom_1(77921) <= 13039115;
srom_1(77922) <= 12550406;
srom_1(77923) <= 12042180;
srom_1(77924) <= 11516822;
srom_1(77925) <= 10976795;
srom_1(77926) <= 10424631;
srom_1(77927) <= 9862919;
srom_1(77928) <= 9294294;
srom_1(77929) <= 8721422;
srom_1(77930) <= 8146988;
srom_1(77931) <= 7573688;
srom_1(77932) <= 7004210;
srom_1(77933) <= 6441223;
srom_1(77934) <= 5887368;
srom_1(77935) <= 5345243;
srom_1(77936) <= 4817388;
srom_1(77937) <= 4306281;
srom_1(77938) <= 3814317;
srom_1(77939) <= 3343803;
srom_1(77940) <= 2896946;
srom_1(77941) <= 2475842;
srom_1(77942) <= 2082464;
srom_1(77943) <= 1718658;
srom_1(77944) <= 1386130;
srom_1(77945) <= 1086438;
srom_1(77946) <= 820990;
srom_1(77947) <= 591028;
srom_1(77948) <= 397632;
srom_1(77949) <= 241708;
srom_1(77950) <= 123988;
srom_1(77951) <= 45023;
srom_1(77952) <= 5185;
srom_1(77953) <= 4659;
srom_1(77954) <= 43448;
srom_1(77955) <= 121371;
srom_1(77956) <= 238061;
srom_1(77957) <= 392973;
srom_1(77958) <= 585378;
srom_1(77959) <= 814376;
srom_1(77960) <= 1078891;
srom_1(77961) <= 1377685;
srom_1(77962) <= 1709355;
srom_1(77963) <= 2072347;
srom_1(77964) <= 2464957;
srom_1(77965) <= 2885346;
srom_1(77966) <= 3331541;
srom_1(77967) <= 3801450;
srom_1(77968) <= 4292871;
srom_1(77969) <= 4803497;
srom_1(77970) <= 5330936;
srom_1(77971) <= 5872713;
srom_1(77972) <= 6426288;
srom_1(77973) <= 6989064;
srom_1(77974) <= 7558404;
srom_1(77975) <= 8131637;
srom_1(77976) <= 8706075;
srom_1(77977) <= 9279024;
srom_1(77978) <= 9847798;
srom_1(77979) <= 10409729;
srom_1(77980) <= 10962182;
srom_1(77981) <= 11502567;
srom_1(77982) <= 12028349;
srom_1(77983) <= 12537064;
srom_1(77984) <= 13026325;
srom_1(77985) <= 13493838;
srom_1(77986) <= 13937411;
srom_1(77987) <= 14354963;
srom_1(77988) <= 14744538;
srom_1(77989) <= 15104307;
srom_1(77990) <= 15432584;
srom_1(77991) <= 15727829;
srom_1(77992) <= 15988658;
srom_1(77993) <= 16213848;
srom_1(77994) <= 16402343;
srom_1(77995) <= 16553258;
srom_1(77996) <= 16665887;
srom_1(77997) <= 16739701;
srom_1(77998) <= 16774353;
srom_1(77999) <= 16769682;
srom_1(78000) <= 16725709;
srom_1(78001) <= 16642641;
srom_1(78002) <= 16520866;
srom_1(78003) <= 16360957;
srom_1(78004) <= 16163663;
srom_1(78005) <= 15929908;
srom_1(78006) <= 15660790;
srom_1(78007) <= 15357570;
srom_1(78008) <= 15021670;
srom_1(78009) <= 14654666;
srom_1(78010) <= 14258278;
srom_1(78011) <= 13834365;
srom_1(78012) <= 13384915;
srom_1(78013) <= 12912035;
srom_1(78014) <= 12417944;
srom_1(78015) <= 11904957;
srom_1(78016) <= 11375481;
srom_1(78017) <= 10831999;
srom_1(78018) <= 10277059;
srom_1(78019) <= 9713263;
srom_1(78020) <= 9143256;
srom_1(78021) <= 8569709;
srom_1(78022) <= 7995314;
srom_1(78023) <= 7422763;
srom_1(78024) <= 6854740;
srom_1(78025) <= 6293911;
srom_1(78026) <= 5742905;
srom_1(78027) <= 5204305;
srom_1(78028) <= 4680637;
srom_1(78029) <= 4174357;
srom_1(78030) <= 3687840;
srom_1(78031) <= 3223365;
srom_1(78032) <= 2783113;
srom_1(78033) <= 2369146;
srom_1(78034) <= 1983407;
srom_1(78035) <= 1627704;
srom_1(78036) <= 1303705;
srom_1(78037) <= 1012930;
srom_1(78038) <= 756742;
srom_1(78039) <= 536342;
srom_1(78040) <= 352765;
srom_1(78041) <= 206870;
srom_1(78042) <= 99342;
srom_1(78043) <= 30685;
srom_1(78044) <= 1221;
srom_1(78045) <= 11089;
srom_1(78046) <= 60242;
srom_1(78047) <= 148449;
srom_1(78048) <= 275297;
srom_1(78049) <= 440192;
srom_1(78050) <= 642359;
srom_1(78051) <= 880851;
srom_1(78052) <= 1154550;
srom_1(78053) <= 1462171;
srom_1(78054) <= 1802273;
srom_1(78055) <= 2173260;
srom_1(78056) <= 2573394;
srom_1(78057) <= 3000797;
srom_1(78058) <= 3453465;
srom_1(78059) <= 3929276;
srom_1(78060) <= 4425998;
srom_1(78061) <= 4941302;
srom_1(78062) <= 5472772;
srom_1(78063) <= 6017915;
srom_1(78064) <= 6574175;
srom_1(78065) <= 7138943;
srom_1(78066) <= 7709572;
srom_1(78067) <= 8283385;
srom_1(78068) <= 8857691;
srom_1(78069) <= 9429798;
srom_1(78070) <= 9997022;
srom_1(78071) <= 10556704;
srom_1(78072) <= 11106218;
srom_1(78073) <= 11642989;
srom_1(78074) <= 12164499;
srom_1(78075) <= 12668303;
srom_1(78076) <= 13152038;
srom_1(78077) <= 13613435;
srom_1(78078) <= 14050331;
srom_1(78079) <= 14460677;
srom_1(78080) <= 14842550;
srom_1(78081) <= 15194157;
srom_1(78082) <= 15513852;
srom_1(78083) <= 15800133;
srom_1(78084) <= 16051659;
srom_1(78085) <= 16267251;
srom_1(78086) <= 16445896;
srom_1(78087) <= 16586759;
srom_1(78088) <= 16689177;
srom_1(78089) <= 16752671;
srom_1(78090) <= 16776944;
srom_1(78091) <= 16761880;
srom_1(78092) <= 16707551;
srom_1(78093) <= 16614212;
srom_1(78094) <= 16482301;
srom_1(78095) <= 16312435;
srom_1(78096) <= 16105411;
srom_1(78097) <= 15862201;
srom_1(78098) <= 15583945;
srom_1(78099) <= 15271947;
srom_1(78100) <= 14927671;
srom_1(78101) <= 14552730;
srom_1(78102) <= 14148885;
srom_1(78103) <= 13718027;
srom_1(78104) <= 13262178;
srom_1(78105) <= 12783475;
srom_1(78106) <= 12284162;
srom_1(78107) <= 11766583;
srom_1(78108) <= 11233163;
srom_1(78109) <= 10686403;
srom_1(78110) <= 10128869;
srom_1(78111) <= 9563174;
srom_1(78112) <= 8991971;
srom_1(78113) <= 8417938;
srom_1(78114) <= 7843768;
srom_1(78115) <= 7272153;
srom_1(78116) <= 6705773;
srom_1(78117) <= 6147285;
srom_1(78118) <= 5599307;
srom_1(78119) <= 5064409;
srom_1(78120) <= 4545099;
srom_1(78121) <= 4043813;
srom_1(78122) <= 3562901;
srom_1(78123) <= 3104619;
srom_1(78124) <= 2671115;
srom_1(78125) <= 2264422;
srom_1(78126) <= 1886447;
srom_1(78127) <= 1538964;
srom_1(78128) <= 1223601;
srom_1(78129) <= 941837;
srom_1(78130) <= 694993;
srom_1(78131) <= 484228;
srom_1(78132) <= 310528;
srom_1(78133) <= 174710;
srom_1(78134) <= 77409;
srom_1(78135) <= 19083;
srom_1(78136) <= 4;
srom_1(78137) <= 20262;
srom_1(78138) <= 79762;
srom_1(78139) <= 178225;
srom_1(78140) <= 315190;
srom_1(78141) <= 490013;
srom_1(78142) <= 701876;
srom_1(78143) <= 949784;
srom_1(78144) <= 1232576;
srom_1(78145) <= 1548925;
srom_1(78146) <= 1897347;
srom_1(78147) <= 2276209;
srom_1(78148) <= 2683734;
srom_1(78149) <= 3118012;
srom_1(78150) <= 3577005;
srom_1(78151) <= 4058561;
srom_1(78152) <= 4560422;
srom_1(78153) <= 5080235;
srom_1(78154) <= 5615562;
srom_1(78155) <= 6163893;
srom_1(78156) <= 6722656;
srom_1(78157) <= 7289232;
srom_1(78158) <= 7860962;
srom_1(78159) <= 8435167;
srom_1(78160) <= 9009154;
srom_1(78161) <= 9580231;
srom_1(78162) <= 10145720;
srom_1(78163) <= 10702969;
srom_1(78164) <= 11249365;
srom_1(78165) <= 11782347;
srom_1(78166) <= 12299413;
srom_1(78167) <= 12798141;
srom_1(78168) <= 13276191;
srom_1(78169) <= 13731321;
srom_1(78170) <= 14161398;
srom_1(78171) <= 14564404;
srom_1(78172) <= 14938449;
srom_1(78173) <= 15281780;
srom_1(78174) <= 15592787;
srom_1(78175) <= 15870010;
srom_1(78176) <= 16112151;
srom_1(78177) <= 16318073;
srom_1(78178) <= 16486812;
srom_1(78179) <= 16617575;
srom_1(78180) <= 16709750;
srom_1(78181) <= 16762904;
srom_1(78182) <= 16776788;
srom_1(78183) <= 16751337;
srom_1(78184) <= 16686670;
srom_1(78185) <= 16583091;
srom_1(78186) <= 16441085;
srom_1(78187) <= 16261318;
srom_1(78188) <= 16044634;
srom_1(78189) <= 15792047;
srom_1(78190) <= 15504743;
srom_1(78191) <= 15184070;
srom_1(78192) <= 14831530;
srom_1(78193) <= 14448777;
srom_1(78194) <= 14037606;
srom_1(78195) <= 13599944;
srom_1(78196) <= 13137845;
srom_1(78197) <= 12653475;
srom_1(78198) <= 12149106;
srom_1(78199) <= 11627102;
srom_1(78200) <= 11089912;
srom_1(78201) <= 10540055;
srom_1(78202) <= 9980109;
srom_1(78203) <= 9412699;
srom_1(78204) <= 8840488;
srom_1(78205) <= 8266157;
srom_1(78206) <= 7692401;
srom_1(78207) <= 7121909;
srom_1(78208) <= 6557357;
srom_1(78209) <= 6001393;
srom_1(78210) <= 5456623;
srom_1(78211) <= 4925602;
srom_1(78212) <= 4410820;
srom_1(78213) <= 3914692;
srom_1(78214) <= 3439543;
srom_1(78215) <= 2987602;
srom_1(78216) <= 2560988;
srom_1(78217) <= 2161702;
srom_1(78218) <= 1791617;
srom_1(78219) <= 1452466;
srom_1(78220) <= 1145842;
srom_1(78221) <= 873181;
srom_1(78222) <= 635763;
srom_1(78223) <= 434701;
srom_1(78224) <= 270937;
srom_1(78225) <= 145239;
srom_1(78226) <= 58198;
srom_1(78227) <= 10221;
srom_1(78228) <= 1533;
srom_1(78229) <= 32175;
srom_1(78230) <= 102003;
srom_1(78231) <= 210690;
srom_1(78232) <= 357725;
srom_1(78233) <= 542421;
srom_1(78234) <= 763910;
srom_1(78235) <= 1021153;
srom_1(78236) <= 1312945;
srom_1(78237) <= 1637918;
srom_1(78238) <= 1994546;
srom_1(78239) <= 2381159;
srom_1(78240) <= 2795943;
srom_1(78241) <= 3236952;
srom_1(78242) <= 3702120;
srom_1(78243) <= 4189264;
srom_1(78244) <= 4696100;
srom_1(78245) <= 5220251;
srom_1(78246) <= 5759260;
srom_1(78247) <= 6310599;
srom_1(78248) <= 6871683;
srom_1(78249) <= 7439880;
srom_1(78250) <= 8012525;
srom_1(78251) <= 8586935;
srom_1(78252) <= 9160414;
srom_1(78253) <= 9730274;
srom_1(78254) <= 10293842;
srom_1(78255) <= 10848477;
srom_1(78256) <= 11391576;
srom_1(78257) <= 11920593;
srom_1(78258) <= 12433047;
srom_1(78259) <= 12926535;
srom_1(78260) <= 13398744;
srom_1(78261) <= 13847459;
srom_1(78262) <= 14270574;
srom_1(78263) <= 14666108;
srom_1(78264) <= 15032204;
srom_1(78265) <= 15367146;
srom_1(78266) <= 15669363;
srom_1(78267) <= 15937438;
srom_1(78268) <= 16170114;
srom_1(78269) <= 16366300;
srom_1(78270) <= 16525076;
srom_1(78271) <= 16645697;
srom_1(78272) <= 16727598;
srom_1(78273) <= 16770394;
srom_1(78274) <= 16773886;
srom_1(78275) <= 16738056;
srom_1(78276) <= 16663072;
srom_1(78277) <= 16549287;
srom_1(78278) <= 16397233;
srom_1(78279) <= 16207624;
srom_1(78280) <= 15981349;
srom_1(78281) <= 15719469;
srom_1(78282) <= 15423213;
srom_1(78283) <= 15093968;
srom_1(78284) <= 14733280;
srom_1(78285) <= 14342839;
srom_1(78286) <= 13924477;
srom_1(78287) <= 13480156;
srom_1(78288) <= 13011958;
srom_1(78289) <= 12522080;
srom_1(78290) <= 12012818;
srom_1(78291) <= 11486562;
srom_1(78292) <= 10945778;
srom_1(78293) <= 10393002;
srom_1(78294) <= 9830828;
srom_1(78295) <= 9261890;
srom_1(78296) <= 8688857;
srom_1(78297) <= 8114416;
srom_1(78298) <= 7541261;
srom_1(78299) <= 6972079;
srom_1(78300) <= 6409540;
srom_1(78301) <= 5856282;
srom_1(78302) <= 5314898;
srom_1(78303) <= 4787928;
srom_1(78304) <= 4277843;
srom_1(78305) <= 3787035;
srom_1(78306) <= 3317805;
srom_1(78307) <= 2872354;
srom_1(78308) <= 2452770;
srom_1(78309) <= 2061022;
srom_1(78310) <= 1698945;
srom_1(78311) <= 1368239;
srom_1(78312) <= 1070454;
srom_1(78313) <= 806986;
srom_1(78314) <= 579071;
srom_1(78315) <= 387778;
srom_1(78316) <= 234003;
srom_1(78317) <= 118468;
srom_1(78318) <= 41714;
srom_1(78319) <= 4102;
srom_1(78320) <= 5808;
srom_1(78321) <= 46823;
srom_1(78322) <= 126956;
srom_1(78323) <= 245831;
srom_1(78324) <= 402890;
srom_1(78325) <= 597397;
srom_1(78326) <= 828439;
srom_1(78327) <= 1094934;
srom_1(78328) <= 1395631;
srom_1(78329) <= 1729121;
srom_1(78330) <= 2093839;
srom_1(78331) <= 2488076;
srom_1(78332) <= 2909982;
srom_1(78333) <= 3357579;
srom_1(78334) <= 3828769;
srom_1(78335) <= 4321341;
srom_1(78336) <= 4832986;
srom_1(78337) <= 5361305;
srom_1(78338) <= 5903819;
srom_1(78339) <= 6457986;
srom_1(78340) <= 7021206;
srom_1(78341) <= 7590838;
srom_1(78342) <= 8164211;
srom_1(78343) <= 8738637;
srom_1(78344) <= 9311421;
srom_1(78345) <= 9879878;
srom_1(78346) <= 10441341;
srom_1(78347) <= 10993179;
srom_1(78348) <= 11532803;
srom_1(78349) <= 12057682;
srom_1(78350) <= 12565356;
srom_1(78351) <= 13053444;
srom_1(78352) <= 13519657;
srom_1(78353) <= 13961809;
srom_1(78354) <= 14377826;
srom_1(78355) <= 14765757;
srom_1(78356) <= 15123784;
srom_1(78357) <= 15450227;
srom_1(78358) <= 15743556;
srom_1(78359) <= 16002395;
srom_1(78360) <= 16225530;
srom_1(78361) <= 16411915;
srom_1(78362) <= 16560677;
srom_1(78363) <= 16671116;
srom_1(78364) <= 16742716;
srom_1(78365) <= 16775141;
srom_1(78366) <= 16768238;
srom_1(78367) <= 16722041;
srom_1(78368) <= 16636765;
srom_1(78369) <= 16512811;
srom_1(78370) <= 16350759;
srom_1(78371) <= 16151370;
srom_1(78372) <= 15915579;
srom_1(78373) <= 15644492;
srom_1(78374) <= 15339379;
srom_1(78375) <= 15001671;
srom_1(78376) <= 14632953;
srom_1(78377) <= 14234952;
srom_1(78378) <= 13809536;
srom_1(78379) <= 13358700;
srom_1(78380) <= 12884557;
srom_1(78381) <= 12389331;
srom_1(78382) <= 11875344;
srom_1(78383) <= 11345007;
srom_1(78384) <= 10800806;
srom_1(78385) <= 10245294;
srom_1(78386) <= 9681074;
srom_1(78387) <= 9110794;
srom_1(78388) <= 8537128;
srom_1(78389) <= 7962765;
srom_1(78390) <= 7390399;
srom_1(78391) <= 6822714;
srom_1(78392) <= 6262371;
srom_1(78393) <= 5712000;
srom_1(78394) <= 5174180;
srom_1(78395) <= 4651434;
srom_1(78396) <= 4146212;
srom_1(78397) <= 3660885;
srom_1(78398) <= 3197727;
srom_1(78399) <= 2758911;
srom_1(78400) <= 2346495;
srom_1(78401) <= 1962412;
srom_1(78402) <= 1608464;
srom_1(78403) <= 1286311;
srom_1(78404) <= 997462;
srom_1(78405) <= 743273;
srom_1(78406) <= 524936;
srom_1(78407) <= 343474;
srom_1(78408) <= 199739;
srom_1(78409) <= 94404;
srom_1(78410) <= 27963;
srom_1(78411) <= 728;
srom_1(78412) <= 12827;
srom_1(78413) <= 64203;
srom_1(78414) <= 154615;
srom_1(78415) <= 283639;
srom_1(78416) <= 450669;
srom_1(78417) <= 654924;
srom_1(78418) <= 895444;
srom_1(78419) <= 1171103;
srom_1(78420) <= 1480607;
srom_1(78421) <= 1822504;
srom_1(78422) <= 2195193;
srom_1(78423) <= 2596924;
srom_1(78424) <= 3025815;
srom_1(78425) <= 3479854;
srom_1(78426) <= 3956911;
srom_1(78427) <= 4454750;
srom_1(78428) <= 4971037;
srom_1(78429) <= 5503349;
srom_1(78430) <= 6049192;
srom_1(78431) <= 6606005;
srom_1(78432) <= 7171177;
srom_1(78433) <= 7742058;
srom_1(78434) <= 8315971;
srom_1(78435) <= 8890224;
srom_1(78436) <= 9462126;
srom_1(78437) <= 10028993;
srom_1(78438) <= 10588168;
srom_1(78439) <= 11137028;
srom_1(78440) <= 11673000;
srom_1(78441) <= 12193571;
srom_1(78442) <= 12696298;
srom_1(78443) <= 13178826;
srom_1(78444) <= 13638890;
srom_1(78445) <= 14074334;
srom_1(78446) <= 14483116;
srom_1(78447) <= 14863318;
srom_1(78448) <= 15213159;
srom_1(78449) <= 15530996;
srom_1(78450) <= 15815341;
srom_1(78451) <= 16064859;
srom_1(78452) <= 16278380;
srom_1(78453) <= 16454904;
srom_1(78454) <= 16593602;
srom_1(78455) <= 16693823;
srom_1(78456) <= 16755099;
srom_1(78457) <= 16777142;
srom_1(78458) <= 16759848;
srom_1(78459) <= 16703298;
srom_1(78460) <= 16607757;
srom_1(78461) <= 16473675;
srom_1(78462) <= 16301678;
srom_1(78463) <= 16092575;
srom_1(78464) <= 15847345;
srom_1(78465) <= 15567138;
srom_1(78466) <= 15253269;
srom_1(78467) <= 14907209;
srom_1(78468) <= 14530581;
srom_1(78469) <= 14125151;
srom_1(78470) <= 13692821;
srom_1(78471) <= 13235617;
srom_1(78472) <= 12755684;
srom_1(78473) <= 12255272;
srom_1(78474) <= 11736728;
srom_1(78475) <= 11202484;
srom_1(78476) <= 10655045;
srom_1(78477) <= 10096977;
srom_1(78478) <= 9530898;
srom_1(78479) <= 8959463;
srom_1(78480) <= 8385350;
srom_1(78481) <= 7811253;
srom_1(78482) <= 7239863;
srom_1(78483) <= 6673861;
srom_1(78484) <= 6115899;
srom_1(78485) <= 5568595;
srom_1(78486) <= 5034514;
srom_1(78487) <= 4516162;
srom_1(78488) <= 4015970;
srom_1(78489) <= 3536282;
srom_1(78490) <= 3079349;
srom_1(78491) <= 2647312;
srom_1(78492) <= 2242198;
srom_1(78493) <= 1865907;
srom_1(78494) <= 1520203;
srom_1(78495) <= 1206708;
srom_1(78496) <= 926890;
srom_1(78497) <= 682064;
srom_1(78498) <= 473376;
srom_1(78499) <= 301805;
srom_1(78500) <= 168156;
srom_1(78501) <= 73055;
srom_1(78502) <= 16949;
srom_1(78503) <= 101;
srom_1(78504) <= 22589;
srom_1(78505) <= 84308;
srom_1(78506) <= 184969;
srom_1(78507) <= 324100;
srom_1(78508) <= 501048;
srom_1(78509) <= 714983;
srom_1(78510) <= 964903;
srom_1(78511) <= 1249634;
srom_1(78512) <= 1567843;
srom_1(78513) <= 1918037;
srom_1(78514) <= 2298574;
srom_1(78515) <= 2707669;
srom_1(78516) <= 3143404;
srom_1(78517) <= 3603735;
srom_1(78518) <= 4086504;
srom_1(78519) <= 4589447;
srom_1(78520) <= 5110206;
srom_1(78521) <= 5646339;
srom_1(78522) <= 6195330;
srom_1(78523) <= 6754607;
srom_1(78524) <= 7321546;
srom_1(78525) <= 7893489;
srom_1(78526) <= 8467754;
srom_1(78527) <= 9041648;
srom_1(78528) <= 9612479;
srom_1(78529) <= 10177571;
srom_1(78530) <= 10734274;
srom_1(78531) <= 11279978;
srom_1(78532) <= 11812123;
srom_1(78533) <= 12328213;
srom_1(78534) <= 12825830;
srom_1(78535) <= 13302639;
srom_1(78536) <= 13756404;
srom_1(78537) <= 14184998;
srom_1(78538) <= 14586411;
srom_1(78539) <= 14958760;
srom_1(78540) <= 15300299;
srom_1(78541) <= 15609427;
srom_1(78542) <= 15884694;
srom_1(78543) <= 16124809;
srom_1(78544) <= 16328647;
srom_1(78545) <= 16495251;
srom_1(78546) <= 16623840;
srom_1(78547) <= 16713812;
srom_1(78548) <= 16764743;
srom_1(78549) <= 16776396;
srom_1(78550) <= 16748716;
srom_1(78551) <= 16681832;
srom_1(78552) <= 16576059;
srom_1(78553) <= 16431892;
srom_1(78554) <= 16250007;
srom_1(78555) <= 16031257;
srom_1(78556) <= 15776668;
srom_1(78557) <= 15487435;
srom_1(78558) <= 15164912;
srom_1(78559) <= 14810613;
srom_1(78560) <= 14426199;
srom_1(78561) <= 14013472;
srom_1(78562) <= 13574369;
srom_1(78563) <= 13110947;
srom_1(78564) <= 12625381;
srom_1(78565) <= 12119948;
srom_1(78566) <= 11597017;
srom_1(78567) <= 11059040;
srom_1(78568) <= 10508541;
srom_1(78569) <= 9948101;
srom_1(78570) <= 9380348;
srom_1(78571) <= 8807944;
srom_1(78572) <= 8233574;
srom_1(78573) <= 7659930;
srom_1(78574) <= 7089704;
srom_1(78575) <= 6525569;
srom_1(78576) <= 5970170;
srom_1(78577) <= 5426112;
srom_1(78578) <= 4895947;
srom_1(78579) <= 4382159;
srom_1(78580) <= 3887159;
srom_1(78581) <= 3413268;
srom_1(78582) <= 2962708;
srom_1(78583) <= 2537592;
srom_1(78584) <= 2139914;
srom_1(78585) <= 1771537;
srom_1(78586) <= 1434191;
srom_1(78587) <= 1129456;
srom_1(78588) <= 858761;
srom_1(78589) <= 623377;
srom_1(78590) <= 424406;
srom_1(78591) <= 262783;
srom_1(78592) <= 139264;
srom_1(78593) <= 54429;
srom_1(78594) <= 8676;
srom_1(78595) <= 2219;
srom_1(78596) <= 35089;
srom_1(78597) <= 107132;
srom_1(78598) <= 218009;
srom_1(78599) <= 367201;
srom_1(78600) <= 554008;
srom_1(78601) <= 777554;
srom_1(78602) <= 1036791;
srom_1(78603) <= 1330503;
srom_1(78604) <= 1657313;
srom_1(78605) <= 2015689;
srom_1(78606) <= 2403949;
srom_1(78607) <= 2820273;
srom_1(78608) <= 3262710;
srom_1(78609) <= 3729183;
srom_1(78610) <= 4217506;
srom_1(78611) <= 4725388;
srom_1(78612) <= 5250449;
srom_1(78613) <= 5790226;
srom_1(78614) <= 6342187;
srom_1(78615) <= 6903745;
srom_1(78616) <= 7472265;
srom_1(78617) <= 8045083;
srom_1(78618) <= 8619512;
srom_1(78619) <= 9192858;
srom_1(78620) <= 9762432;
srom_1(78621) <= 10325564;
srom_1(78622) <= 10879613;
srom_1(78623) <= 11421981;
srom_1(78624) <= 11950124;
srom_1(78625) <= 12461566;
srom_1(78626) <= 12953909;
srom_1(78627) <= 13424843;
srom_1(78628) <= 13872161;
srom_1(78629) <= 14293764;
srom_1(78630) <= 14687677;
srom_1(78631) <= 15052050;
srom_1(78632) <= 15385177;
srom_1(78633) <= 15685494;
srom_1(78634) <= 15951593;
srom_1(78635) <= 16182227;
srom_1(78636) <= 16376314;
srom_1(78637) <= 16532944;
srom_1(78638) <= 16651383;
srom_1(78639) <= 16731074;
srom_1(78640) <= 16771645;
srom_1(78641) <= 16772905;
srom_1(78642) <= 16734848;
srom_1(78643) <= 16657652;
srom_1(78644) <= 16541680;
srom_1(78645) <= 16387476;
srom_1(78646) <= 16195762;
srom_1(78647) <= 15967437;
srom_1(78648) <= 15703573;
srom_1(78649) <= 15405407;
srom_1(78650) <= 15074336;
srom_1(78651) <= 14711914;
srom_1(78652) <= 14319839;
srom_1(78653) <= 13899951;
srom_1(78654) <= 13454219;
srom_1(78655) <= 12984732;
srom_1(78656) <= 12493692;
srom_1(78657) <= 11983402;
srom_1(78658) <= 11456254;
srom_1(78659) <= 10914722;
srom_1(78660) <= 10361343;
srom_1(78661) <= 9798714;
srom_1(78662) <= 9229473;
srom_1(78663) <= 8656288;
srom_1(78664) <= 8081848;
srom_1(78665) <= 7508846;
srom_1(78666) <= 6939970;
srom_1(78667) <= 6377887;
srom_1(78668) <= 5825233;
srom_1(78669) <= 5284600;
srom_1(78670) <= 4758522;
srom_1(78671) <= 4249467;
srom_1(78672) <= 3759822;
srom_1(78673) <= 3291883;
srom_1(78674) <= 2847844;
srom_1(78675) <= 2429788;
srom_1(78676) <= 2039675;
srom_1(78677) <= 1679334;
srom_1(78678) <= 1350455;
srom_1(78679) <= 1054580;
srom_1(78680) <= 793097;
srom_1(78681) <= 567232;
srom_1(78682) <= 378045;
srom_1(78683) <= 226421;
srom_1(78684) <= 113073;
srom_1(78685) <= 38531;
srom_1(78686) <= 3146;
srom_1(78687) <= 7084;
srom_1(78688) <= 50325;
srom_1(78689) <= 132667;
srom_1(78690) <= 253724;
srom_1(78691) <= 412928;
srom_1(78692) <= 609533;
srom_1(78693) <= 842617;
srom_1(78694) <= 1111087;
srom_1(78695) <= 1413683;
srom_1(78696) <= 1748987;
srom_1(78697) <= 2115427;
srom_1(78698) <= 2511284;
srom_1(78699) <= 2934701;
srom_1(78700) <= 3383694;
srom_1(78701) <= 3856156;
srom_1(78702) <= 4349873;
srom_1(78703) <= 4862529;
srom_1(78704) <= 5391719;
srom_1(78705) <= 5934963;
srom_1(78706) <= 6489714;
srom_1(78707) <= 7053368;
srom_1(78708) <= 7623284;
srom_1(78709) <= 8196789;
srom_1(78710) <= 8771194;
srom_1(78711) <= 9343804;
srom_1(78712) <= 9911935;
srom_1(78713) <= 10472923;
srom_1(78714) <= 11024136;
srom_1(78715) <= 11562991;
srom_1(78716) <= 12086960;
srom_1(78717) <= 12593586;
srom_1(78718) <= 13080493;
srom_1(78719) <= 13545399;
srom_1(78720) <= 13986123;
srom_1(78721) <= 14400598;
srom_1(78722) <= 14786880;
srom_1(78723) <= 15143159;
srom_1(78724) <= 15467764;
srom_1(78725) <= 15759172;
srom_1(78726) <= 16016016;
srom_1(78727) <= 16237094;
srom_1(78728) <= 16421367;
srom_1(78729) <= 16567971;
srom_1(78730) <= 16676220;
srom_1(78731) <= 16745606;
srom_1(78732) <= 16775802;
srom_1(78733) <= 16766668;
srom_1(78734) <= 16718247;
srom_1(78735) <= 16630764;
srom_1(78736) <= 16504632;
srom_1(78737) <= 16340441;
srom_1(78738) <= 16138961;
srom_1(78739) <= 15901136;
srom_1(78740) <= 15628083;
srom_1(78741) <= 15321082;
srom_1(78742) <= 14981572;
srom_1(78743) <= 14611145;
srom_1(78744) <= 14211538;
srom_1(78745) <= 13784626;
srom_1(78746) <= 13332410;
srom_1(78747) <= 12857011;
srom_1(78748) <= 12360658;
srom_1(78749) <= 11845679;
srom_1(78750) <= 11314488;
srom_1(78751) <= 10769576;
srom_1(78752) <= 10213500;
srom_1(78753) <= 9648866;
srom_1(78754) <= 9078322;
srom_1(78755) <= 8504544;
srom_1(78756) <= 7930222;
srom_1(78757) <= 7358050;
srom_1(78758) <= 6790711;
srom_1(78759) <= 6230864;
srom_1(78760) <= 5681136;
srom_1(78761) <= 5144104;
srom_1(78762) <= 4622287;
srom_1(78763) <= 4118131;
srom_1(78764) <= 3634001;
srom_1(78765) <= 3172167;
srom_1(78766) <= 2734795;
srom_1(78767) <= 2323935;
srom_1(78768) <= 1941515;
srom_1(78769) <= 1589327;
srom_1(78770) <= 1269023;
srom_1(78771) <= 982106;
srom_1(78772) <= 729920;
srom_1(78773) <= 513649;
srom_1(78774) <= 334305;
srom_1(78775) <= 192732;
srom_1(78776) <= 89591;
srom_1(78777) <= 25368;
srom_1(78778) <= 362;
srom_1(78779) <= 14692;
srom_1(78780) <= 68290;
srom_1(78781) <= 160905;
srom_1(78782) <= 292102;
srom_1(78783) <= 461267;
srom_1(78784) <= 667606;
srom_1(78785) <= 910151;
srom_1(78786) <= 1187765;
srom_1(78787) <= 1499146;
srom_1(78788) <= 1842835;
srom_1(78789) <= 2217219;
srom_1(78790) <= 2620542;
srom_1(78791) <= 3050914;
srom_1(78792) <= 3506316;
srom_1(78793) <= 3984613;
srom_1(78794) <= 4483562;
srom_1(78795) <= 5000823;
srom_1(78796) <= 5533971;
srom_1(78797) <= 6080504;
srom_1(78798) <= 6637862;
srom_1(78799) <= 7203429;
srom_1(78800) <= 7774554;
srom_1(78801) <= 8348558;
srom_1(78802) <= 8922750;
srom_1(78803) <= 9494437;
srom_1(78804) <= 10060939;
srom_1(78805) <= 10619599;
srom_1(78806) <= 11167796;
srom_1(78807) <= 11702962;
srom_1(78808) <= 12222585;
srom_1(78809) <= 12724229;
srom_1(78810) <= 13205542;
srom_1(78811) <= 13664266;
srom_1(78812) <= 14098251;
srom_1(78813) <= 14505462;
srom_1(78814) <= 14883989;
srom_1(78815) <= 15232057;
srom_1(78816) <= 15548033;
srom_1(78817) <= 15830436;
srom_1(78818) <= 16077942;
srom_1(78819) <= 16289391;
srom_1(78820) <= 16463789;
srom_1(78821) <= 16600320;
srom_1(78822) <= 16698344;
srom_1(78823) <= 16757401;
srom_1(78824) <= 16777213;
srom_1(78825) <= 16757689;
srom_1(78826) <= 16698918;
srom_1(78827) <= 16601178;
srom_1(78828) <= 16464927;
srom_1(78829) <= 16290802;
srom_1(78830) <= 16079622;
srom_1(78831) <= 15832376;
srom_1(78832) <= 15550223;
srom_1(78833) <= 15234487;
srom_1(78834) <= 14886649;
srom_1(78835) <= 14508339;
srom_1(78836) <= 14101331;
srom_1(78837) <= 13667535;
srom_1(78838) <= 13208983;
srom_1(78839) <= 12727828;
srom_1(78840) <= 12226324;
srom_1(78841) <= 11706824;
srom_1(78842) <= 11171763;
srom_1(78843) <= 10623652;
srom_1(78844) <= 10065059;
srom_1(78845) <= 9498605;
srom_1(78846) <= 8926946;
srom_1(78847) <= 8352763;
srom_1(78848) <= 7778747;
srom_1(78849) <= 7207591;
srom_1(78850) <= 6641974;
srom_1(78851) <= 6084547;
srom_1(78852) <= 5537925;
srom_1(78853) <= 5004670;
srom_1(78854) <= 4487284;
srom_1(78855) <= 3988193;
srom_1(78856) <= 3509736;
srom_1(78857) <= 3054158;
srom_1(78858) <= 2623596;
srom_1(78859) <= 2220067;
srom_1(78860) <= 1845465;
srom_1(78861) <= 1501546;
srom_1(78862) <= 1189923;
srom_1(78863) <= 912056;
srom_1(78864) <= 669250;
srom_1(78865) <= 462643;
srom_1(78866) <= 293203;
srom_1(78867) <= 161725;
srom_1(78868) <= 68826;
srom_1(78869) <= 14942;
srom_1(78870) <= 324;
srom_1(78871) <= 25042;
srom_1(78872) <= 88979;
srom_1(78873) <= 191837;
srom_1(78874) <= 333131;
srom_1(78875) <= 512201;
srom_1(78876) <= 728206;
srom_1(78877) <= 980133;
srom_1(78878) <= 1266801;
srom_1(78879) <= 1586865;
srom_1(78880) <= 1938825;
srom_1(78881) <= 2321031;
srom_1(78882) <= 2731689;
srom_1(78883) <= 3168875;
srom_1(78884) <= 3630538;
srom_1(78885) <= 4114513;
srom_1(78886) <= 4618530;
srom_1(78887) <= 5140227;
srom_1(78888) <= 5677157;
srom_1(78889) <= 6226801;
srom_1(78890) <= 6786583;
srom_1(78891) <= 7353878;
srom_1(78892) <= 7926024;
srom_1(78893) <= 8500340;
srom_1(78894) <= 9074132;
srom_1(78895) <= 9644709;
srom_1(78896) <= 10209396;
srom_1(78897) <= 10765545;
srom_1(78898) <= 11310547;
srom_1(78899) <= 11841847;
srom_1(78900) <= 12356954;
srom_1(78901) <= 12853452;
srom_1(78902) <= 13329013;
srom_1(78903) <= 13781406;
srom_1(78904) <= 14208511;
srom_1(78905) <= 14608324;
srom_1(78906) <= 14978971;
srom_1(78907) <= 15318714;
srom_1(78908) <= 15625958;
srom_1(78909) <= 15899265;
srom_1(78910) <= 16137351;
srom_1(78911) <= 16339101;
srom_1(78912) <= 16503568;
srom_1(78913) <= 16629981;
srom_1(78914) <= 16717748;
srom_1(78915) <= 16766456;
srom_1(78916) <= 16775878;
srom_1(78917) <= 16745969;
srom_1(78918) <= 16676870;
srom_1(78919) <= 16568904;
srom_1(78920) <= 16422577;
srom_1(78921) <= 16238577;
srom_1(78922) <= 16017766;
srom_1(78923) <= 15761178;
srom_1(78924) <= 15470019;
srom_1(78925) <= 15145652;
srom_1(78926) <= 14789599;
srom_1(78927) <= 14403529;
srom_1(78928) <= 13989253;
srom_1(78929) <= 13548715;
srom_1(78930) <= 13083978;
srom_1(78931) <= 12597224;
srom_1(78932) <= 12090733;
srom_1(78933) <= 11566882;
srom_1(78934) <= 11028128;
srom_1(78935) <= 10476995;
srom_1(78936) <= 9916069;
srom_1(78937) <= 9347981;
srom_1(78938) <= 8775394;
srom_1(78939) <= 8200993;
srom_1(78940) <= 7627471;
srom_1(78941) <= 7057519;
srom_1(78942) <= 6493809;
srom_1(78943) <= 5938984;
srom_1(78944) <= 5395647;
srom_1(78945) <= 4866344;
srom_1(78946) <= 4353559;
srom_1(78947) <= 3859695;
srom_1(78948) <= 3387069;
srom_1(78949) <= 2937896;
srom_1(78950) <= 2514284;
srom_1(78951) <= 2118219;
srom_1(78952) <= 1751558;
srom_1(78953) <= 1416020;
srom_1(78954) <= 1113179;
srom_1(78955) <= 844455;
srom_1(78956) <= 611108;
srom_1(78957) <= 414232;
srom_1(78958) <= 254751;
srom_1(78959) <= 133413;
srom_1(78960) <= 50786;
srom_1(78961) <= 7257;
srom_1(78962) <= 3032;
srom_1(78963) <= 38130;
srom_1(78964) <= 112386;
srom_1(78965) <= 225452;
srom_1(78966) <= 376798;
srom_1(78967) <= 565714;
srom_1(78968) <= 791314;
srom_1(78969) <= 1052540;
srom_1(78970) <= 1348168;
srom_1(78971) <= 1676811;
srom_1(78972) <= 2036928;
srom_1(78973) <= 2426829;
srom_1(78974) <= 2844688;
srom_1(78975) <= 3288544;
srom_1(78976) <= 3756316;
srom_1(78977) <= 4245811;
srom_1(78978) <= 4754732;
srom_1(78979) <= 5280694;
srom_1(78980) <= 5821230;
srom_1(78981) <= 6373806;
srom_1(78982) <= 6935829;
srom_1(78983) <= 7504665;
srom_1(78984) <= 8077646;
srom_1(78985) <= 8652085;
srom_1(78986) <= 9225289;
srom_1(78987) <= 9794569;
srom_1(78988) <= 10357257;
srom_1(78989) <= 10910712;
srom_1(78990) <= 11452341;
srom_1(78991) <= 11979602;
srom_1(78992) <= 12490024;
srom_1(78993) <= 12981214;
srom_1(78994) <= 13450867;
srom_1(78995) <= 13896781;
srom_1(78996) <= 14316865;
srom_1(78997) <= 14709150;
srom_1(78998) <= 15071796;
srom_1(78999) <= 15403102;
srom_1(79000) <= 15701514;
srom_1(79001) <= 15965634;
srom_1(79002) <= 16194223;
srom_1(79003) <= 16386208;
srom_1(79004) <= 16540690;
srom_1(79005) <= 16656944;
srom_1(79006) <= 16734424;
srom_1(79007) <= 16772769;
srom_1(79008) <= 16771797;
srom_1(79009) <= 16731514;
srom_1(79010) <= 16652107;
srom_1(79011) <= 16533951;
srom_1(79012) <= 16377598;
srom_1(79013) <= 16183782;
srom_1(79014) <= 15953411;
srom_1(79015) <= 15687567;
srom_1(79016) <= 15387495;
srom_1(79017) <= 15054604;
srom_1(79018) <= 14690453;
srom_1(79019) <= 14296750;
srom_1(79020) <= 13875342;
srom_1(79021) <= 13428205;
srom_1(79022) <= 12957436;
srom_1(79023) <= 12465242;
srom_1(79024) <= 11953931;
srom_1(79025) <= 11425901;
srom_1(79026) <= 10883628;
srom_1(79027) <= 10329655;
srom_1(79028) <= 9766580;
srom_1(79029) <= 9197043;
srom_1(79030) <= 8623715;
srom_1(79031) <= 8049284;
srom_1(79032) <= 7476445;
srom_1(79033) <= 6907883;
srom_1(79034) <= 6346265;
srom_1(79035) <= 5794224;
srom_1(79036) <= 5254349;
srom_1(79037) <= 4729171;
srom_1(79038) <= 4221154;
srom_1(79039) <= 3732680;
srom_1(79040) <= 3266039;
srom_1(79041) <= 2823419;
srom_1(79042) <= 2406896;
srom_1(79043) <= 2018424;
srom_1(79044) <= 1659823;
srom_1(79045) <= 1332777;
srom_1(79046) <= 1038817;
srom_1(79047) <= 779323;
srom_1(79048) <= 555512;
srom_1(79049) <= 368432;
srom_1(79050) <= 218962;
srom_1(79051) <= 107803;
srom_1(79052) <= 35475;
srom_1(79053) <= 2317;
srom_1(79054) <= 8486;
srom_1(79055) <= 53952;
srom_1(79056) <= 138502;
srom_1(79057) <= 261740;
srom_1(79058) <= 423087;
srom_1(79059) <= 621787;
srom_1(79060) <= 856909;
srom_1(79061) <= 1127349;
srom_1(79062) <= 1431840;
srom_1(79063) <= 1768954;
srom_1(79064) <= 2137109;
srom_1(79065) <= 2534580;
srom_1(79066) <= 2959502;
srom_1(79067) <= 3409884;
srom_1(79068) <= 3883612;
srom_1(79069) <= 4378466;
srom_1(79070) <= 4892124;
srom_1(79071) <= 5422179;
srom_1(79072) <= 5966145;
srom_1(79073) <= 6521470;
srom_1(79074) <= 7085551;
srom_1(79075) <= 7655742;
srom_1(79076) <= 8229370;
srom_1(79077) <= 8803745;
srom_1(79078) <= 9376172;
srom_1(79079) <= 9943969;
srom_1(79080) <= 10504473;
srom_1(79081) <= 11055054;
srom_1(79082) <= 11593131;
srom_1(79083) <= 12116182;
srom_1(79084) <= 12621752;
srom_1(79085) <= 13107472;
srom_1(79086) <= 13571063;
srom_1(79087) <= 14010352;
srom_1(79088) <= 14423279;
srom_1(79089) <= 14807907;
srom_1(79090) <= 15162433;
srom_1(79091) <= 15485194;
srom_1(79092) <= 15774676;
srom_1(79093) <= 16029523;
srom_1(79094) <= 16248539;
srom_1(79095) <= 16430697;
srom_1(79096) <= 16575143;
srom_1(79097) <= 16681199;
srom_1(79098) <= 16748369;
srom_1(79099) <= 16776337;
srom_1(79100) <= 16764971;
srom_1(79101) <= 16714327;
srom_1(79102) <= 16624640;
srom_1(79103) <= 16496331;
srom_1(79104) <= 16330003;
srom_1(79105) <= 16126434;
srom_1(79106) <= 15886580;
srom_1(79107) <= 15611566;
srom_1(79108) <= 15302681;
srom_1(79109) <= 14961373;
srom_1(79110) <= 14589243;
srom_1(79111) <= 14188037;
srom_1(79112) <= 13759635;
srom_1(79113) <= 13306046;
srom_1(79114) <= 12829398;
srom_1(79115) <= 12331925;
srom_1(79116) <= 11815961;
srom_1(79117) <= 11283924;
srom_1(79118) <= 10738311;
srom_1(79119) <= 10181679;
srom_1(79120) <= 9616639;
srom_1(79121) <= 9045840;
srom_1(79122) <= 8471959;
srom_1(79123) <= 7897687;
srom_1(79124) <= 7325717;
srom_1(79125) <= 6758731;
srom_1(79126) <= 6199389;
srom_1(79127) <= 5650313;
srom_1(79128) <= 5114077;
srom_1(79129) <= 4593197;
srom_1(79130) <= 4090114;
srom_1(79131) <= 3607189;
srom_1(79132) <= 3146686;
srom_1(79133) <= 2710763;
srom_1(79134) <= 2301466;
srom_1(79135) <= 1920714;
srom_1(79136) <= 1570292;
srom_1(79137) <= 1251843;
srom_1(79138) <= 966861;
srom_1(79139) <= 716682;
srom_1(79140) <= 502480;
srom_1(79141) <= 325258;
srom_1(79142) <= 185848;
srom_1(79143) <= 84904;
srom_1(79144) <= 22898;
srom_1(79145) <= 122;
srom_1(79146) <= 16683;
srom_1(79147) <= 72503;
srom_1(79148) <= 167319;
srom_1(79149) <= 300688;
srom_1(79150) <= 471984;
srom_1(79151) <= 680404;
srom_1(79152) <= 924970;
srom_1(79153) <= 1204536;
srom_1(79154) <= 1517790;
srom_1(79155) <= 1863264;
srom_1(79156) <= 2239338;
srom_1(79157) <= 2644247;
srom_1(79158) <= 3076094;
srom_1(79159) <= 3532853;
srom_1(79160) <= 4012382;
srom_1(79161) <= 4512433;
srom_1(79162) <= 5030661;
srom_1(79163) <= 5564635;
srom_1(79164) <= 6111852;
srom_1(79165) <= 6669745;
srom_1(79166) <= 7235699;
srom_1(79167) <= 7807059;
srom_1(79168) <= 8381146;
srom_1(79169) <= 8955268;
srom_1(79170) <= 9526732;
srom_1(79171) <= 10092860;
srom_1(79172) <= 10650996;
srom_1(79173) <= 11198523;
srom_1(79174) <= 11732873;
srom_1(79175) <= 12251541;
srom_1(79176) <= 12752094;
srom_1(79177) <= 13232185;
srom_1(79178) <= 13689563;
srom_1(79179) <= 14122083;
srom_1(79180) <= 14527716;
srom_1(79181) <= 14904562;
srom_1(79182) <= 15250851;
srom_1(79183) <= 15564962;
srom_1(79184) <= 15845420;
srom_1(79185) <= 16090910;
srom_1(79186) <= 16300282;
srom_1(79187) <= 16472553;
srom_1(79188) <= 16606916;
srom_1(79189) <= 16702740;
srom_1(79190) <= 16759576;
srom_1(79191) <= 16777158;
srom_1(79192) <= 16755403;
srom_1(79193) <= 16694414;
srom_1(79194) <= 16594475;
srom_1(79195) <= 16456057;
srom_1(79196) <= 16279807;
srom_1(79197) <= 16066553;
srom_1(79198) <= 15817295;
srom_1(79199) <= 15533200;
srom_1(79200) <= 15215603;
srom_1(79201) <= 14865991;
srom_1(79202) <= 14486004;
srom_1(79203) <= 14077425;
srom_1(79204) <= 13642169;
srom_1(79205) <= 13182277;
srom_1(79206) <= 12699906;
srom_1(79207) <= 12197317;
srom_1(79208) <= 11676869;
srom_1(79209) <= 11141000;
srom_1(79210) <= 10592225;
srom_1(79211) <= 10033116;
srom_1(79212) <= 9466296;
srom_1(79213) <= 8894421;
srom_1(79214) <= 8320175;
srom_1(79215) <= 7746250;
srom_1(79216) <= 7175337;
srom_1(79217) <= 6610114;
srom_1(79218) <= 6053230;
srom_1(79219) <= 5507298;
srom_1(79220) <= 4974877;
srom_1(79221) <= 4458464;
srom_1(79222) <= 3960482;
srom_1(79223) <= 3483264;
srom_1(79224) <= 3029049;
srom_1(79225) <= 2599967;
srom_1(79226) <= 2198029;
srom_1(79227) <= 1825122;
srom_1(79228) <= 1482993;
srom_1(79229) <= 1173246;
srom_1(79230) <= 897335;
srom_1(79231) <= 656554;
srom_1(79232) <= 452030;
srom_1(79233) <= 284724;
srom_1(79234) <= 155419;
srom_1(79235) <= 64723;
srom_1(79236) <= 13061;
srom_1(79237) <= 674;
srom_1(79238) <= 27621;
srom_1(79239) <= 93776;
srom_1(79240) <= 198828;
srom_1(79241) <= 342284;
srom_1(79242) <= 523473;
srom_1(79243) <= 741544;
srom_1(79244) <= 995475;
srom_1(79245) <= 1284074;
srom_1(79246) <= 1605989;
srom_1(79247) <= 1959711;
srom_1(79248) <= 2343579;
srom_1(79249) <= 2755795;
srom_1(79250) <= 3194425;
srom_1(79251) <= 3657412;
srom_1(79252) <= 4142585;
srom_1(79253) <= 4647670;
srom_1(79254) <= 5170297;
srom_1(79255) <= 5708016;
srom_1(79256) <= 6258305;
srom_1(79257) <= 6818583;
srom_1(79258) <= 7386224;
srom_1(79259) <= 7958566;
srom_1(79260) <= 8532924;
srom_1(79261) <= 9106605;
srom_1(79262) <= 9676920;
srom_1(79263) <= 10241193;
srom_1(79264) <= 10796779;
srom_1(79265) <= 11341072;
srom_1(79266) <= 11871520;
srom_1(79267) <= 12385635;
srom_1(79268) <= 12881007;
srom_1(79269) <= 13355312;
srom_1(79270) <= 13806327;
srom_1(79271) <= 14231936;
srom_1(79272) <= 14630144;
srom_1(79273) <= 14999083;
srom_1(79274) <= 15337024;
srom_1(79275) <= 15642381;
srom_1(79276) <= 15913722;
srom_1(79277) <= 16149776;
srom_1(79278) <= 16349434;
srom_1(79279) <= 16511762;
srom_1(79280) <= 16635998;
srom_1(79281) <= 16721558;
srom_1(79282) <= 16768043;
srom_1(79283) <= 16775233;
srom_1(79284) <= 16743096;
srom_1(79285) <= 16671782;
srom_1(79286) <= 16561625;
srom_1(79287) <= 16413142;
srom_1(79288) <= 16227029;
srom_1(79289) <= 16004159;
srom_1(79290) <= 15745577;
srom_1(79291) <= 15452496;
srom_1(79292) <= 15126289;
srom_1(79293) <= 14768488;
srom_1(79294) <= 14380769;
srom_1(79295) <= 13964950;
srom_1(79296) <= 13522983;
srom_1(79297) <= 13056938;
srom_1(79298) <= 12569002;
srom_1(79299) <= 12061463;
srom_1(79300) <= 11536700;
srom_1(79301) <= 10997175;
srom_1(79302) <= 10445418;
srom_1(79303) <= 9884015;
srom_1(79304) <= 9315600;
srom_1(79305) <= 8742838;
srom_1(79306) <= 8168414;
srom_1(79307) <= 7595024;
srom_1(79308) <= 7025354;
srom_1(79309) <= 6462078;
srom_1(79310) <= 5907836;
srom_1(79311) <= 5365226;
srom_1(79312) <= 4836795;
srom_1(79313) <= 4325019;
srom_1(79314) <= 3832299;
srom_1(79315) <= 3360944;
srom_1(79316) <= 2913167;
srom_1(79317) <= 2491065;
srom_1(79318) <= 2096619;
srom_1(79319) <= 1731678;
srom_1(79320) <= 1397954;
srom_1(79321) <= 1097012;
srom_1(79322) <= 830262;
srom_1(79323) <= 598956;
srom_1(79324) <= 404179;
srom_1(79325) <= 246843;
srom_1(79326) <= 127686;
srom_1(79327) <= 47268;
srom_1(79328) <= 5965;
srom_1(79329) <= 3972;
srom_1(79330) <= 41297;
srom_1(79331) <= 117765;
srom_1(79332) <= 233018;
srom_1(79333) <= 386515;
srom_1(79334) <= 577537;
srom_1(79335) <= 805188;
srom_1(79336) <= 1068400;
srom_1(79337) <= 1365939;
srom_1(79338) <= 1696409;
srom_1(79339) <= 2058262;
srom_1(79340) <= 2449800;
srom_1(79341) <= 2869187;
srom_1(79342) <= 3314456;
srom_1(79343) <= 3783520;
srom_1(79344) <= 4274179;
srom_1(79345) <= 4784131;
srom_1(79346) <= 5310986;
srom_1(79347) <= 5852274;
srom_1(79348) <= 6405455;
srom_1(79349) <= 6967935;
srom_1(79350) <= 7537078;
srom_1(79351) <= 8110214;
srom_1(79352) <= 8684655;
srom_1(79353) <= 9257708;
srom_1(79354) <= 9826686;
srom_1(79355) <= 10388919;
srom_1(79356) <= 10941773;
srom_1(79357) <= 11482654;
srom_1(79358) <= 12009026;
srom_1(79359) <= 12518421;
srom_1(79360) <= 13008449;
srom_1(79361) <= 13476813;
srom_1(79362) <= 13921318;
srom_1(79363) <= 14339877;
srom_1(79364) <= 14730529;
srom_1(79365) <= 15091441;
srom_1(79366) <= 15420921;
srom_1(79367) <= 15717425;
srom_1(79368) <= 15979561;
srom_1(79369) <= 16206100;
srom_1(79370) <= 16395981;
srom_1(79371) <= 16548312;
srom_1(79372) <= 16662380;
srom_1(79373) <= 16737649;
srom_1(79374) <= 16773766;
srom_1(79375) <= 16770563;
srom_1(79376) <= 16728054;
srom_1(79377) <= 16646438;
srom_1(79378) <= 16526098;
srom_1(79379) <= 16367599;
srom_1(79380) <= 16171684;
srom_1(79381) <= 15939271;
srom_1(79382) <= 15671450;
srom_1(79383) <= 15369478;
srom_1(79384) <= 15034770;
srom_1(79385) <= 14668896;
srom_1(79386) <= 14273572;
srom_1(79387) <= 13850650;
srom_1(79388) <= 13402116;
srom_1(79389) <= 12930071;
srom_1(79390) <= 12436730;
srom_1(79391) <= 11924406;
srom_1(79392) <= 11395501;
srom_1(79393) <= 10852496;
srom_1(79394) <= 10297937;
srom_1(79395) <= 9734424;
srom_1(79396) <= 9164600;
srom_1(79397) <= 8591138;
srom_1(79398) <= 8016726;
srom_1(79399) <= 7444057;
srom_1(79400) <= 6875818;
srom_1(79401) <= 6314673;
srom_1(79402) <= 5763253;
srom_1(79403) <= 5224145;
srom_1(79404) <= 4699875;
srom_1(79405) <= 4192904;
srom_1(79406) <= 3705607;
srom_1(79407) <= 3240271;
srom_1(79408) <= 2799077;
srom_1(79409) <= 2384094;
srom_1(79410) <= 1997269;
srom_1(79411) <= 1640415;
srom_1(79412) <= 1315205;
srom_1(79413) <= 1023165;
srom_1(79414) <= 765664;
srom_1(79415) <= 543909;
srom_1(79416) <= 358941;
srom_1(79417) <= 211627;
srom_1(79418) <= 102658;
srom_1(79419) <= 32544;
srom_1(79420) <= 1614;
srom_1(79421) <= 10015;
srom_1(79422) <= 57705;
srom_1(79423) <= 144461;
srom_1(79424) <= 269878;
srom_1(79425) <= 433366;
srom_1(79426) <= 634158;
srom_1(79427) <= 871314;
srom_1(79428) <= 1143721;
srom_1(79429) <= 1450102;
srom_1(79430) <= 1789020;
srom_1(79431) <= 2158886;
srom_1(79432) <= 2557965;
srom_1(79433) <= 2984386;
srom_1(79434) <= 3436149;
srom_1(79435) <= 3911136;
srom_1(79436) <= 4407119;
srom_1(79437) <= 4921773;
srom_1(79438) <= 5452684;
srom_1(79439) <= 5997362;
srom_1(79440) <= 6553254;
srom_1(79441) <= 7117753;
srom_1(79442) <= 7688211;
srom_1(79443) <= 8261953;
srom_1(79444) <= 8836289;
srom_1(79445) <= 9408526;
srom_1(79446) <= 9975980;
srom_1(79447) <= 10535991;
srom_1(79448) <= 11085931;
srom_1(79449) <= 11623223;
srom_1(79450) <= 12145347;
srom_1(79451) <= 12649854;
srom_1(79452) <= 13134379;
srom_1(79453) <= 13596649;
srom_1(79454) <= 14034497;
srom_1(79455) <= 14445869;
srom_1(79456) <= 14828837;
srom_1(79457) <= 15181604;
srom_1(79458) <= 15502516;
srom_1(79459) <= 15790069;
srom_1(79460) <= 16042914;
srom_1(79461) <= 16259865;
srom_1(79462) <= 16439906;
srom_1(79463) <= 16582191;
srom_1(79464) <= 16686053;
srom_1(79465) <= 16751006;
srom_1(79466) <= 16776744;
srom_1(79467) <= 16763148;
srom_1(79468) <= 16710281;
srom_1(79469) <= 16618390;
srom_1(79470) <= 16487908;
srom_1(79471) <= 16319444;
srom_1(79472) <= 16113791;
srom_1(79473) <= 15871911;
srom_1(79474) <= 15594940;
srom_1(79475) <= 15284175;
srom_1(79476) <= 14941075;
srom_1(79477) <= 14567248;
srom_1(79478) <= 14164448;
srom_1(79479) <= 13734562;
srom_1(79480) <= 13279607;
srom_1(79481) <= 12801717;
srom_1(79482) <= 12303133;
srom_1(79483) <= 11786191;
srom_1(79484) <= 11253317;
srom_1(79485) <= 10707010;
srom_1(79486) <= 10149831;
srom_1(79487) <= 9584393;
srom_1(79488) <= 9013347;
srom_1(79489) <= 8439372;
srom_1(79490) <= 7865159;
srom_1(79491) <= 7293400;
srom_1(79492) <= 6726777;
srom_1(79493) <= 6167947;
srom_1(79494) <= 5619531;
srom_1(79495) <= 5084099;
srom_1(79496) <= 4564164;
srom_1(79497) <= 4062162;
srom_1(79498) <= 3580449;
srom_1(79499) <= 3121283;
srom_1(79500) <= 2686818;
srom_1(79501) <= 2279090;
srom_1(79502) <= 1900011;
srom_1(79503) <= 1551360;
srom_1(79504) <= 1234771;
srom_1(79505) <= 951729;
srom_1(79506) <= 703561;
srom_1(79507) <= 491430;
srom_1(79508) <= 316333;
srom_1(79509) <= 179088;
srom_1(79510) <= 80342;
srom_1(79511) <= 20555;
srom_1(79512) <= 9;
srom_1(79513) <= 18800;
srom_1(79514) <= 76841;
srom_1(79515) <= 173857;
srom_1(79516) <= 309396;
srom_1(79517) <= 482821;
srom_1(79518) <= 693318;
srom_1(79519) <= 939902;
srom_1(79520) <= 1221415;
srom_1(79521) <= 1536538;
srom_1(79522) <= 1883792;
srom_1(79523) <= 2261549;
srom_1(79524) <= 2668039;
srom_1(79525) <= 3101354;
srom_1(79526) <= 3559463;
srom_1(79527) <= 4040217;
srom_1(79528) <= 4541363;
srom_1(79529) <= 5060549;
srom_1(79530) <= 5595342;
srom_1(79531) <= 6143234;
srom_1(79532) <= 6701654;
srom_1(79533) <= 7267986;
srom_1(79534) <= 7839572;
srom_1(79535) <= 8413733;
srom_1(79536) <= 8987777;
srom_1(79537) <= 9559010;
srom_1(79538) <= 10124755;
srom_1(79539) <= 10682359;
srom_1(79540) <= 11229207;
srom_1(79541) <= 11762734;
srom_1(79542) <= 12280438;
srom_1(79543) <= 12779893;
srom_1(79544) <= 13258755;
srom_1(79545) <= 13714779;
srom_1(79546) <= 14145827;
srom_1(79547) <= 14549878;
srom_1(79548) <= 14925036;
srom_1(79549) <= 15269543;
srom_1(79550) <= 15581782;
srom_1(79551) <= 15860291;
srom_1(79552) <= 16103762;
srom_1(79553) <= 16311054;
srom_1(79554) <= 16481195;
srom_1(79555) <= 16613387;
srom_1(79556) <= 16707010;
srom_1(79557) <= 16761625;
srom_1(79558) <= 16776976;
srom_1(79559) <= 16752992;
srom_1(79560) <= 16689784;
srom_1(79561) <= 16587649;
srom_1(79562) <= 16447065;
srom_1(79563) <= 16268693;
srom_1(79564) <= 16053369;
srom_1(79565) <= 15802101;
srom_1(79566) <= 15516070;
srom_1(79567) <= 15196615;
srom_1(79568) <= 14845235;
srom_1(79569) <= 14463578;
srom_1(79570) <= 14053433;
srom_1(79571) <= 13616723;
srom_1(79572) <= 13155498;
srom_1(79573) <= 12671919;
srom_1(79574) <= 12168253;
srom_1(79575) <= 11646864;
srom_1(79576) <= 11110196;
srom_1(79577) <= 10560765;
srom_1(79578) <= 10001148;
srom_1(79579) <= 9433970;
srom_1(79580) <= 8861889;
srom_1(79581) <= 8287589;
srom_1(79582) <= 7713763;
srom_1(79583) <= 7143101;
srom_1(79584) <= 6578280;
srom_1(79585) <= 6021948;
srom_1(79586) <= 5476714;
srom_1(79587) <= 4945135;
srom_1(79588) <= 4429704;
srom_1(79589) <= 3932837;
srom_1(79590) <= 3456865;
srom_1(79591) <= 3004020;
srom_1(79592) <= 2576425;
srom_1(79593) <= 2176085;
srom_1(79594) <= 1804878;
srom_1(79595) <= 1464544;
srom_1(79596) <= 1156679;
srom_1(79597) <= 882728;
srom_1(79598) <= 643974;
srom_1(79599) <= 441537;
srom_1(79600) <= 276367;
srom_1(79601) <= 149238;
srom_1(79602) <= 60746;
srom_1(79603) <= 11306;
srom_1(79604) <= 1151;
srom_1(79605) <= 30327;
srom_1(79606) <= 98697;
srom_1(79607) <= 205943;
srom_1(79608) <= 351559;
srom_1(79609) <= 534864;
srom_1(79610) <= 754998;
srom_1(79611) <= 1010928;
srom_1(79612) <= 1301455;
srom_1(79613) <= 1625216;
srom_1(79614) <= 1980693;
srom_1(79615) <= 2366219;
srom_1(79616) <= 2779986;
srom_1(79617) <= 3220053;
srom_1(79618) <= 3684358;
srom_1(79619) <= 4170722;
srom_1(79620) <= 4676866;
srom_1(79621) <= 5200415;
srom_1(79622) <= 5738915;
srom_1(79623) <= 6289840;
srom_1(79624) <= 6850607;
srom_1(79625) <= 7418586;
srom_1(79626) <= 7991114;
srom_1(79627) <= 8565506;
srom_1(79628) <= 9139068;
srom_1(79629) <= 9709111;
srom_1(79630) <= 10272962;
srom_1(79631) <= 10827977;
srom_1(79632) <= 11371552;
srom_1(79633) <= 11901139;
srom_1(79634) <= 12414255;
srom_1(79635) <= 12908494;
srom_1(79636) <= 13381537;
srom_1(79637) <= 13831166;
srom_1(79638) <= 14255273;
srom_1(79639) <= 14651870;
srom_1(79640) <= 15019096;
srom_1(79641) <= 15355229;
srom_1(79642) <= 15658693;
srom_1(79643) <= 15928066;
srom_1(79644) <= 16162083;
srom_1(79645) <= 16359648;
srom_1(79646) <= 16519834;
srom_1(79647) <= 16641890;
srom_1(79648) <= 16725243;
srom_1(79649) <= 16769503;
srom_1(79650) <= 16774462;
srom_1(79651) <= 16740097;
srom_1(79652) <= 16666569;
srom_1(79653) <= 16554222;
srom_1(79654) <= 16403585;
srom_1(79655) <= 16215362;
srom_1(79656) <= 15990437;
srom_1(79657) <= 15729864;
srom_1(79658) <= 15434866;
srom_1(79659) <= 15106825;
srom_1(79660) <= 14747281;
srom_1(79661) <= 14357918;
srom_1(79662) <= 13940563;
srom_1(79663) <= 13497173;
srom_1(79664) <= 13029828;
srom_1(79665) <= 12540718;
srom_1(79666) <= 12032137;
srom_1(79667) <= 11506471;
srom_1(79668) <= 10966183;
srom_1(79669) <= 10413809;
srom_1(79670) <= 9851938;
srom_1(79671) <= 9283205;
srom_1(79672) <= 8710276;
srom_1(79673) <= 8135840;
srom_1(79674) <= 7562588;
srom_1(79675) <= 6993210;
srom_1(79676) <= 6430376;
srom_1(79677) <= 5876724;
srom_1(79678) <= 5334852;
srom_1(79679) <= 4807299;
srom_1(79680) <= 4296541;
srom_1(79681) <= 3804971;
srom_1(79682) <= 3334896;
srom_1(79683) <= 2888520;
srom_1(79684) <= 2467935;
srom_1(79685) <= 2075114;
srom_1(79686) <= 1711900;
srom_1(79687) <= 1379994;
srom_1(79688) <= 1080955;
srom_1(79689) <= 816184;
srom_1(79690) <= 586922;
srom_1(79691) <= 394245;
srom_1(79692) <= 239057;
srom_1(79693) <= 122084;
srom_1(79694) <= 43876;
srom_1(79695) <= 4800;
srom_1(79696) <= 5038;
srom_1(79697) <= 44589;
srom_1(79698) <= 123268;
srom_1(79699) <= 240707;
srom_1(79700) <= 396353;
srom_1(79701) <= 589479;
srom_1(79702) <= 819176;
srom_1(79703) <= 1084370;
srom_1(79704) <= 1383815;
srom_1(79705) <= 1716109;
srom_1(79706) <= 2079692;
srom_1(79707) <= 2472860;
srom_1(79708) <= 2893769;
srom_1(79709) <= 3340444;
srom_1(79710) <= 3810793;
srom_1(79711) <= 4302608;
srom_1(79712) <= 4813584;
srom_1(79713) <= 5341325;
srom_1(79714) <= 5883355;
srom_1(79715) <= 6437134;
srom_1(79716) <= 7000063;
srom_1(79717) <= 7569504;
srom_1(79718) <= 8142786;
srom_1(79719) <= 8717220;
srom_1(79720) <= 9290114;
srom_1(79721) <= 9858780;
srom_1(79722) <= 10420552;
srom_1(79723) <= 10972795;
srom_1(79724) <= 11512921;
srom_1(79725) <= 12038395;
srom_1(79726) <= 12546754;
srom_1(79727) <= 13035615;
srom_1(79728) <= 13502683;
srom_1(79729) <= 13945771;
srom_1(79730) <= 14362798;
srom_1(79731) <= 14751811;
srom_1(79732) <= 15110985;
srom_1(79733) <= 15438634;
srom_1(79734) <= 15733224;
srom_1(79735) <= 15993373;
srom_1(79736) <= 16217860;
srom_1(79737) <= 16405633;
srom_1(79738) <= 16555811;
srom_1(79739) <= 16667691;
srom_1(79740) <= 16740747;
srom_1(79741) <= 16774637;
srom_1(79742) <= 16769202;
srom_1(79743) <= 16724468;
srom_1(79744) <= 16640644;
srom_1(79745) <= 16518123;
srom_1(79746) <= 16357480;
srom_1(79747) <= 16159469;
srom_1(79748) <= 15925017;
srom_1(79749) <= 15655224;
srom_1(79750) <= 15351356;
srom_1(79751) <= 15014837;
srom_1(79752) <= 14647245;
srom_1(79753) <= 14250304;
srom_1(79754) <= 13825876;
srom_1(79755) <= 13375951;
srom_1(79756) <= 12902638;
srom_1(79757) <= 12408157;
srom_1(79758) <= 11894828;
srom_1(79759) <= 11365056;
srom_1(79760) <= 10821327;
srom_1(79761) <= 10266190;
srom_1(79762) <= 9702248;
srom_1(79763) <= 9132147;
srom_1(79764) <= 8558558;
srom_1(79765) <= 7984173;
srom_1(79766) <= 7411684;
srom_1(79767) <= 6843776;
srom_1(79768) <= 6283113;
srom_1(79769) <= 5732322;
srom_1(79770) <= 5193989;
srom_1(79771) <= 4670635;
srom_1(79772) <= 4164717;
srom_1(79773) <= 3678606;
srom_1(79774) <= 3214581;
srom_1(79775) <= 2774820;
srom_1(79776) <= 2361383;
srom_1(79777) <= 1976210;
srom_1(79778) <= 1621108;
srom_1(79779) <= 1297740;
srom_1(79780) <= 1007623;
srom_1(79781) <= 752119;
srom_1(79782) <= 532425;
srom_1(79783) <= 349571;
srom_1(79784) <= 204415;
srom_1(79785) <= 97637;
srom_1(79786) <= 29739;
srom_1(79787) <= 1038;
srom_1(79788) <= 11670;
srom_1(79789) <= 61583;
srom_1(79790) <= 150545;
srom_1(79791) <= 278139;
srom_1(79792) <= 443764;
srom_1(79793) <= 646646;
srom_1(79794) <= 885833;
srom_1(79795) <= 1160203;
srom_1(79796) <= 1468469;
srom_1(79797) <= 1809186;
srom_1(79798) <= 2180757;
srom_1(79799) <= 2581438;
srom_1(79800) <= 3009350;
srom_1(79801) <= 3462489;
srom_1(79802) <= 3938727;
srom_1(79803) <= 4435832;
srom_1(79804) <= 4951473;
srom_1(79805) <= 5483232;
srom_1(79806) <= 6028616;
srom_1(79807) <= 6585066;
srom_1(79808) <= 7149974;
srom_1(79809) <= 7720690;
srom_1(79810) <= 8294538;
srom_1(79811) <= 8868827;
srom_1(79812) <= 9440864;
srom_1(79813) <= 10007967;
srom_1(79814) <= 10567477;
srom_1(79815) <= 11116768;
srom_1(79816) <= 11653267;
srom_1(79817) <= 12174456;
srom_1(79818) <= 12677892;
srom_1(79819) <= 13161214;
srom_1(79820) <= 13622156;
srom_1(79821) <= 14058556;
srom_1(79822) <= 14468368;
srom_1(79823) <= 14849669;
srom_1(79824) <= 15200672;
srom_1(79825) <= 15519732;
srom_1(79826) <= 15805351;
srom_1(79827) <= 16056190;
srom_1(79828) <= 16271073;
srom_1(79829) <= 16448993;
srom_1(79830) <= 16589115;
srom_1(79831) <= 16690782;
srom_1(79832) <= 16753517;
srom_1(79833) <= 16777026;
srom_1(79834) <= 16761199;
srom_1(79835) <= 16706110;
srom_1(79836) <= 16612017;
srom_1(79837) <= 16479362;
srom_1(79838) <= 16308767;
srom_1(79839) <= 16101031;
srom_1(79840) <= 15857129;
srom_1(79841) <= 15578205;
srom_1(79842) <= 15265566;
srom_1(79843) <= 14920678;
srom_1(79844) <= 14545160;
srom_1(79845) <= 14140771;
srom_1(79846) <= 13709409;
srom_1(79847) <= 13253095;
srom_1(79848) <= 12773970;
srom_1(79849) <= 12274281;
srom_1(79850) <= 11756370;
srom_1(79851) <= 11222667;
srom_1(79852) <= 10675674;
srom_1(79853) <= 10117956;
srom_1(79854) <= 9552129;
srom_1(79855) <= 8980845;
srom_1(79856) <= 8406784;
srom_1(79857) <= 7832638;
srom_1(79858) <= 7261099;
srom_1(79859) <= 6694848;
srom_1(79860) <= 6136539;
srom_1(79861) <= 5588790;
srom_1(79862) <= 5054171;
srom_1(79863) <= 4535189;
srom_1(79864) <= 4034276;
srom_1(79865) <= 3553782;
srom_1(79866) <= 3095961;
srom_1(79867) <= 2662958;
srom_1(79868) <= 2256805;
srom_1(79869) <= 1879406;
srom_1(79870) <= 1532531;
srom_1(79871) <= 1217807;
srom_1(79872) <= 936708;
srom_1(79873) <= 690555;
srom_1(79874) <= 480500;
srom_1(79875) <= 307529;
srom_1(79876) <= 172453;
srom_1(79877) <= 75905;
srom_1(79878) <= 18338;
srom_1(79879) <= 23;
srom_1(79880) <= 21044;
srom_1(79881) <= 81304;
srom_1(79882) <= 180520;
srom_1(79883) <= 318226;
srom_1(79884) <= 493777;
srom_1(79885) <= 706349;
srom_1(79886) <= 954946;
srom_1(79887) <= 1238402;
srom_1(79888) <= 1555388;
srom_1(79889) <= 1904418;
srom_1(79890) <= 2283854;
srom_1(79891) <= 2691917;
srom_1(79892) <= 3126694;
srom_1(79893) <= 3586145;
srom_1(79894) <= 4068118;
srom_1(79895) <= 4570350;
srom_1(79896) <= 5090488;
srom_1(79897) <= 5626091;
srom_1(79898) <= 6174649;
srom_1(79899) <= 6733589;
srom_1(79900) <= 7300290;
srom_1(79901) <= 7872094;
srom_1(79902) <= 8446321;
srom_1(79903) <= 9020277;
srom_1(79904) <= 9591271;
srom_1(79905) <= 10156625;
srom_1(79906) <= 10713688;
srom_1(79907) <= 11259848;
srom_1(79908) <= 11792544;
srom_1(79909) <= 12309277;
srom_1(79910) <= 12807626;
srom_1(79911) <= 13285251;
srom_1(79912) <= 13739915;
srom_1(79913) <= 14169485;
srom_1(79914) <= 14571946;
srom_1(79915) <= 14945412;
srom_1(79916) <= 15288130;
srom_1(79917) <= 15598494;
srom_1(79918) <= 15875049;
srom_1(79919) <= 16116497;
srom_1(79920) <= 16321706;
srom_1(79921) <= 16489714;
srom_1(79922) <= 16619733;
srom_1(79923) <= 16711154;
srom_1(79924) <= 16763548;
srom_1(79925) <= 16776668;
srom_1(79926) <= 16750454;
srom_1(79927) <= 16685028;
srom_1(79928) <= 16580698;
srom_1(79929) <= 16437952;
srom_1(79930) <= 16257460;
srom_1(79931) <= 16040068;
srom_1(79932) <= 15786796;
srom_1(79933) <= 15498831;
srom_1(79934) <= 15177524;
srom_1(79935) <= 14824382;
srom_1(79936) <= 14441059;
srom_1(79937) <= 14029355;
srom_1(79938) <= 13591199;
srom_1(79939) <= 13128647;
srom_1(79940) <= 12643867;
srom_1(79941) <= 12139132;
srom_1(79942) <= 11616811;
srom_1(79943) <= 11079350;
srom_1(79944) <= 10529272;
srom_1(79945) <= 9969156;
srom_1(79946) <= 9401628;
srom_1(79947) <= 8829350;
srom_1(79948) <= 8255005;
srom_1(79949) <= 7681286;
srom_1(79950) <= 7110884;
srom_1(79951) <= 6546474;
srom_1(79952) <= 5990702;
srom_1(79953) <= 5446175;
srom_1(79954) <= 4915446;
srom_1(79955) <= 4401004;
srom_1(79956) <= 3905261;
srom_1(79957) <= 3430542;
srom_1(79958) <= 2979073;
srom_1(79959) <= 2552971;
srom_1(79960) <= 2154234;
srom_1(79961) <= 1784733;
srom_1(79962) <= 1446199;
srom_1(79963) <= 1140221;
srom_1(79964) <= 868233;
srom_1(79965) <= 631510;
srom_1(79966) <= 431164;
srom_1(79967) <= 268132;
srom_1(79968) <= 143180;
srom_1(79969) <= 56894;
srom_1(79970) <= 9678;
srom_1(79971) <= 1754;
srom_1(79972) <= 33158;
srom_1(79973) <= 103744;
srom_1(79974) <= 213181;
srom_1(79975) <= 360955;
srom_1(79976) <= 546373;
srom_1(79977) <= 768567;
srom_1(79978) <= 1026493;
srom_1(79979) <= 1318943;
srom_1(79980) <= 1644545;
srom_1(79981) <= 2001772;
srom_1(79982) <= 2388949;
srom_1(79983) <= 2804261;
srom_1(79984) <= 3245759;
srom_1(79985) <= 3711375;
srom_1(79986) <= 4198923;
srom_1(79987) <= 4706118;
srom_1(79988) <= 5230582;
srom_1(79989) <= 5769854;
srom_1(79990) <= 6321407;
srom_1(79991) <= 6882654;
srom_1(79992) <= 7450963;
srom_1(79993) <= 8023668;
srom_1(79994) <= 8598085;
srom_1(79995) <= 9171520;
srom_1(79996) <= 9741283;
srom_1(79997) <= 10304703;
srom_1(79998) <= 10859138;
srom_1(79999) <= 11401987;
srom_1(80000) <= 11930706;
srom_1(80001) <= 12442815;
srom_1(80002) <= 12935912;
srom_1(80003) <= 13407686;
srom_1(80004) <= 13855923;
srom_1(80005) <= 14278522;
srom_1(80006) <= 14673501;
srom_1(80007) <= 15039008;
srom_1(80008) <= 15373329;
srom_1(80009) <= 15674896;
srom_1(80010) <= 15942296;
srom_1(80011) <= 16174273;
srom_1(80012) <= 16369741;
srom_1(80013) <= 16527783;
srom_1(80014) <= 16647657;
srom_1(80015) <= 16728802;
srom_1(80016) <= 16770837;
srom_1(80017) <= 16773564;
srom_1(80018) <= 16736972;
srom_1(80019) <= 16661231;
srom_1(80020) <= 16546697;
srom_1(80021) <= 16393907;
srom_1(80022) <= 16203577;
srom_1(80023) <= 15976601;
srom_1(80024) <= 15714041;
srom_1(80025) <= 15417130;
srom_1(80026) <= 15087260;
srom_1(80027) <= 14725978;
srom_1(80028) <= 14334977;
srom_1(80029) <= 13916092;
srom_1(80030) <= 13471287;
srom_1(80031) <= 13002647;
srom_1(80032) <= 12512370;
srom_1(80033) <= 12002756;
srom_1(80034) <= 11476194;
srom_1(80035) <= 10935153;
srom_1(80036) <= 10382170;
srom_1(80037) <= 9819839;
srom_1(80038) <= 9250796;
srom_1(80039) <= 8677710;
srom_1(80040) <= 8103269;
srom_1(80041) <= 7530165;
srom_1(80042) <= 6961087;
srom_1(80043) <= 6398703;
srom_1(80044) <= 5845651;
srom_1(80045) <= 5304523;
srom_1(80046) <= 4777857;
srom_1(80047) <= 4268124;
srom_1(80048) <= 3777713;
srom_1(80049) <= 3308924;
srom_1(80050) <= 2863956;
srom_1(80051) <= 2444894;
srom_1(80052) <= 2053705;
srom_1(80053) <= 1692222;
srom_1(80054) <= 1362140;
srom_1(80055) <= 1065009;
srom_1(80056) <= 802220;
srom_1(80057) <= 575006;
srom_1(80058) <= 384433;
srom_1(80059) <= 231394;
srom_1(80060) <= 116607;
srom_1(80061) <= 40611;
srom_1(80062) <= 3761;
srom_1(80063) <= 6230;
srom_1(80064) <= 48008;
srom_1(80065) <= 128897;
srom_1(80066) <= 248519;
srom_1(80067) <= 406312;
srom_1(80068) <= 601538;
srom_1(80069) <= 833279;
srom_1(80070) <= 1100450;
srom_1(80071) <= 1401798;
srom_1(80072) <= 1735909;
srom_1(80073) <= 2101217;
srom_1(80074) <= 2496009;
srom_1(80075) <= 2918433;
srom_1(80076) <= 3366509;
srom_1(80077) <= 3838135;
srom_1(80078) <= 4331100;
srom_1(80079) <= 4843092;
srom_1(80080) <= 5371710;
srom_1(80081) <= 5914475;
srom_1(80082) <= 6468842;
srom_1(80083) <= 7032212;
srom_1(80084) <= 7601942;
srom_1(80085) <= 8175361;
srom_1(80086) <= 8749781;
srom_1(80087) <= 9322506;
srom_1(80088) <= 9890852;
srom_1(80089) <= 10452154;
srom_1(80090) <= 11003779;
srom_1(80091) <= 11543140;
srom_1(80092) <= 12067709;
srom_1(80093) <= 12575025;
srom_1(80094) <= 13062710;
srom_1(80095) <= 13528476;
srom_1(80096) <= 13970140;
srom_1(80097) <= 14385630;
srom_1(80098) <= 14772998;
srom_1(80099) <= 15130427;
srom_1(80100) <= 15456241;
srom_1(80101) <= 15748913;
srom_1(80102) <= 16007070;
srom_1(80103) <= 16229501;
srom_1(80104) <= 16415164;
srom_1(80105) <= 16563187;
srom_1(80106) <= 16672877;
srom_1(80107) <= 16743719;
srom_1(80108) <= 16775381;
srom_1(80109) <= 16767715;
srom_1(80110) <= 16720756;
srom_1(80111) <= 16634725;
srom_1(80112) <= 16510025;
srom_1(80113) <= 16347241;
srom_1(80114) <= 16147136;
srom_1(80115) <= 15910649;
srom_1(80116) <= 15638888;
srom_1(80117) <= 15333128;
srom_1(80118) <= 14994803;
srom_1(80119) <= 14625499;
srom_1(80120) <= 14226948;
srom_1(80121) <= 13801020;
srom_1(80122) <= 13349710;
srom_1(80123) <= 12875137;
srom_1(80124) <= 12379524;
srom_1(80125) <= 11865197;
srom_1(80126) <= 11334566;
srom_1(80127) <= 10790121;
srom_1(80128) <= 10234415;
srom_1(80129) <= 9670053;
srom_1(80130) <= 9099682;
srom_1(80131) <= 8525976;
srom_1(80132) <= 7951626;
srom_1(80133) <= 7379325;
srom_1(80134) <= 6811757;
srom_1(80135) <= 6251584;
srom_1(80136) <= 5701432;
srom_1(80137) <= 5163881;
srom_1(80138) <= 4641451;
srom_1(80139) <= 4136594;
srom_1(80140) <= 3651675;
srom_1(80141) <= 3188970;
srom_1(80142) <= 2750647;
srom_1(80143) <= 2338763;
srom_1(80144) <= 1955249;
srom_1(80145) <= 1601903;
srom_1(80146) <= 1280382;
srom_1(80147) <= 992194;
srom_1(80148) <= 738690;
srom_1(80149) <= 521059;
srom_1(80150) <= 340322;
srom_1(80151) <= 197327;
srom_1(80152) <= 92742;
srom_1(80153) <= 27061;
srom_1(80154) <= 589;
srom_1(80155) <= 13451;
srom_1(80156) <= 65588;
srom_1(80157) <= 156754;
srom_1(80158) <= 286522;
srom_1(80159) <= 454283;
srom_1(80160) <= 659251;
srom_1(80161) <= 900465;
srom_1(80162) <= 1176793;
srom_1(80163) <= 1486940;
srom_1(80164) <= 1829452;
srom_1(80165) <= 2202721;
srom_1(80166) <= 2604998;
srom_1(80167) <= 3034396;
srom_1(80168) <= 3488903;
srom_1(80169) <= 3966385;
srom_1(80170) <= 4464605;
srom_1(80171) <= 4981226;
srom_1(80172) <= 5513825;
srom_1(80173) <= 6059905;
srom_1(80174) <= 6616905;
srom_1(80175) <= 7182214;
srom_1(80176) <= 7753179;
srom_1(80177) <= 8327124;
srom_1(80178) <= 8901358;
srom_1(80179) <= 9473187;
srom_1(80180) <= 10039930;
srom_1(80181) <= 10598929;
srom_1(80182) <= 11147564;
srom_1(80183) <= 11683261;
srom_1(80184) <= 12203508;
srom_1(80185) <= 12705865;
srom_1(80186) <= 13187978;
srom_1(80187) <= 13647584;
srom_1(80188) <= 14082530;
srom_1(80189) <= 14490775;
srom_1(80190) <= 14870404;
srom_1(80191) <= 15219638;
srom_1(80192) <= 15536839;
srom_1(80193) <= 15820520;
srom_1(80194) <= 16069350;
srom_1(80195) <= 16282162;
srom_1(80196) <= 16457959;
srom_1(80197) <= 16595915;
srom_1(80198) <= 16695385;
srom_1(80199) <= 16755901;
srom_1(80200) <= 16777180;
srom_1(80201) <= 16759123;
srom_1(80202) <= 16701813;
srom_1(80203) <= 16605520;
srom_1(80204) <= 16470694;
srom_1(80205) <= 16297969;
srom_1(80206) <= 16088155;
srom_1(80207) <= 15842234;
srom_1(80208) <= 15561361;
srom_1(80209) <= 15246852;
srom_1(80210) <= 14900183;
srom_1(80211) <= 14522979;
srom_1(80212) <= 14117008;
srom_1(80213) <= 13684175;
srom_1(80214) <= 13226509;
srom_1(80215) <= 12746157;
srom_1(80216) <= 12245371;
srom_1(80217) <= 11726499;
srom_1(80218) <= 11191974;
srom_1(80219) <= 10644304;
srom_1(80220) <= 10086055;
srom_1(80221) <= 9519847;
srom_1(80222) <= 8948334;
srom_1(80223) <= 8374197;
srom_1(80224) <= 7800126;
srom_1(80225) <= 7228816;
srom_1(80226) <= 6662944;
srom_1(80227) <= 6105164;
srom_1(80228) <= 5558092;
srom_1(80229) <= 5024294;
srom_1(80230) <= 4506272;
srom_1(80231) <= 4006455;
srom_1(80232) <= 3527188;
srom_1(80233) <= 3070718;
srom_1(80234) <= 2639185;
srom_1(80235) <= 2234613;
srom_1(80236) <= 1858899;
srom_1(80237) <= 1513806;
srom_1(80238) <= 1200950;
srom_1(80239) <= 921800;
srom_1(80240) <= 677665;
srom_1(80241) <= 469689;
srom_1(80242) <= 298847;
srom_1(80243) <= 165941;
srom_1(80244) <= 71594;
srom_1(80245) <= 16248;
srom_1(80246) <= 163;
srom_1(80247) <= 23414;
srom_1(80248) <= 85893;
srom_1(80249) <= 187306;
srom_1(80250) <= 327177;
srom_1(80251) <= 504852;
srom_1(80252) <= 719496;
srom_1(80253) <= 970103;
srom_1(80254) <= 1255498;
srom_1(80255) <= 1574342;
srom_1(80256) <= 1925141;
srom_1(80257) <= 2306250;
srom_1(80258) <= 2715881;
srom_1(80259) <= 3152113;
srom_1(80260) <= 3612901;
srom_1(80261) <= 4096083;
srom_1(80262) <= 4599395;
srom_1(80263) <= 5120476;
srom_1(80264) <= 5656882;
srom_1(80265) <= 6206098;
srom_1(80266) <= 6765549;
srom_1(80267) <= 7332611;
srom_1(80268) <= 7904624;
srom_1(80269) <= 8478907;
srom_1(80270) <= 9052767;
srom_1(80271) <= 9623513;
srom_1(80272) <= 10188467;
srom_1(80273) <= 10744981;
srom_1(80274) <= 11290446;
srom_1(80275) <= 11822302;
srom_1(80276) <= 12338057;
srom_1(80277) <= 12835292;
srom_1(80278) <= 13311674;
srom_1(80279) <= 13764971;
srom_1(80280) <= 14193056;
srom_1(80281) <= 14593922;
srom_1(80282) <= 14965689;
srom_1(80283) <= 15306613;
srom_1(80284) <= 15615097;
srom_1(80285) <= 15889694;
srom_1(80286) <= 16129115;
srom_1(80287) <= 16332238;
srom_1(80288) <= 16498111;
srom_1(80289) <= 16625956;
srom_1(80290) <= 16715173;
srom_1(80291) <= 16765344;
srom_1(80292) <= 16776233;
srom_1(80293) <= 16747790;
srom_1(80294) <= 16680148;
srom_1(80295) <= 16573624;
srom_1(80296) <= 16428717;
srom_1(80297) <= 16246108;
srom_1(80298) <= 16026652;
srom_1(80299) <= 15771379;
srom_1(80300) <= 15481486;
srom_1(80301) <= 15158331;
srom_1(80302) <= 14803431;
srom_1(80303) <= 14418450;
srom_1(80304) <= 14005192;
srom_1(80305) <= 13565597;
srom_1(80306) <= 13101725;
srom_1(80307) <= 12615751;
srom_1(80308) <= 12109955;
srom_1(80309) <= 11586708;
srom_1(80310) <= 11048464;
srom_1(80311) <= 10497747;
srom_1(80312) <= 9937140;
srom_1(80313) <= 9369271;
srom_1(80314) <= 8796804;
srom_1(80315) <= 8222422;
srom_1(80316) <= 7648820;
srom_1(80317) <= 7078686;
srom_1(80318) <= 6514696;
srom_1(80319) <= 5959492;
srom_1(80320) <= 5415680;
srom_1(80321) <= 4885809;
srom_1(80322) <= 4372363;
srom_1(80323) <= 3877751;
srom_1(80324) <= 3404293;
srom_1(80325) <= 2954207;
srom_1(80326) <= 2529605;
srom_1(80327) <= 2132478;
srom_1(80328) <= 1764688;
srom_1(80329) <= 1427960;
srom_1(80330) <= 1123872;
srom_1(80331) <= 853852;
srom_1(80332) <= 619164;
srom_1(80333) <= 420911;
srom_1(80334) <= 260020;
srom_1(80335) <= 137247;
srom_1(80336) <= 53168;
srom_1(80337) <= 8176;
srom_1(80338) <= 2483;
srom_1(80339) <= 36116;
srom_1(80340) <= 108916;
srom_1(80341) <= 220543;
srom_1(80342) <= 370472;
srom_1(80343) <= 558001;
srom_1(80344) <= 782251;
srom_1(80345) <= 1042169;
srom_1(80346) <= 1336537;
srom_1(80347) <= 1663975;
srom_1(80348) <= 2022947;
srom_1(80349) <= 2411770;
srom_1(80350) <= 2828620;
srom_1(80351) <= 3271543;
srom_1(80352) <= 3738462;
srom_1(80353) <= 4227187;
srom_1(80354) <= 4735426;
srom_1(80355) <= 5260796;
srom_1(80356) <= 5800833;
srom_1(80357) <= 6353006;
srom_1(80358) <= 6914724;
srom_1(80359) <= 7483353;
srom_1(80360) <= 8056228;
srom_1(80361) <= 8630661;
srom_1(80362) <= 9203959;
srom_1(80363) <= 9773434;
srom_1(80364) <= 10336415;
srom_1(80365) <= 10890262;
srom_1(80366) <= 11432377;
srom_1(80367) <= 11960220;
srom_1(80368) <= 12471314;
srom_1(80369) <= 12963262;
srom_1(80370) <= 13433759;
srom_1(80371) <= 13880597;
srom_1(80372) <= 14301681;
srom_1(80373) <= 14695037;
srom_1(80374) <= 15058820;
srom_1(80375) <= 15391324;
srom_1(80376) <= 15690989;
srom_1(80377) <= 15956412;
srom_1(80378) <= 16186346;
srom_1(80379) <= 16379714;
srom_1(80380) <= 16535609;
srom_1(80381) <= 16653300;
srom_1(80382) <= 16732235;
srom_1(80383) <= 16772044;
srom_1(80384) <= 16772540;
srom_1(80385) <= 16733721;
srom_1(80386) <= 16655768;
srom_1(80387) <= 16539048;
srom_1(80388) <= 16384108;
srom_1(80389) <= 16191675;
srom_1(80390) <= 15962650;
srom_1(80391) <= 15698107;
srom_1(80392) <= 15399288;
srom_1(80393) <= 15067594;
srom_1(80394) <= 14704579;
srom_1(80395) <= 14311947;
srom_1(80396) <= 13891538;
srom_1(80397) <= 13445324;
srom_1(80398) <= 12975397;
srom_1(80399) <= 12483961;
srom_1(80400) <= 11973321;
srom_1(80401) <= 11445870;
srom_1(80402) <= 10904084;
srom_1(80403) <= 10350501;
srom_1(80404) <= 9787718;
srom_1(80405) <= 9218374;
srom_1(80406) <= 8645140;
srom_1(80407) <= 8070702;
srom_1(80408) <= 7497755;
srom_1(80409) <= 6928985;
srom_1(80410) <= 6367061;
srom_1(80411) <= 5814615;
srom_1(80412) <= 5274241;
srom_1(80413) <= 4748470;
srom_1(80414) <= 4239770;
srom_1(80415) <= 3750525;
srom_1(80416) <= 3283029;
srom_1(80417) <= 2839475;
srom_1(80418) <= 2421943;
srom_1(80419) <= 2032390;
srom_1(80420) <= 1672645;
srom_1(80421) <= 1344392;
srom_1(80422) <= 1049172;
srom_1(80423) <= 788370;
srom_1(80424) <= 563207;
srom_1(80425) <= 374741;
srom_1(80426) <= 223854;
srom_1(80427) <= 111255;
srom_1(80428) <= 37471;
srom_1(80429) <= 2848;
srom_1(80430) <= 7549;
srom_1(80431) <= 51552;
srom_1(80432) <= 134650;
srom_1(80433) <= 256454;
srom_1(80434) <= 416392;
srom_1(80435) <= 613714;
srom_1(80436) <= 847496;
srom_1(80437) <= 1116641;
srom_1(80438) <= 1419886;
srom_1(80439) <= 1755810;
srom_1(80440) <= 2122837;
srom_1(80441) <= 2519247;
srom_1(80442) <= 2943180;
srom_1(80443) <= 3392649;
srom_1(80444) <= 3865546;
srom_1(80445) <= 4359652;
srom_1(80446) <= 4872652;
srom_1(80447) <= 5402140;
srom_1(80448) <= 5945632;
srom_1(80449) <= 6500579;
srom_1(80450) <= 7064381;
srom_1(80451) <= 7634392;
srom_1(80452) <= 8207940;
srom_1(80453) <= 8782335;
srom_1(80454) <= 9354884;
srom_1(80455) <= 9922902;
srom_1(80456) <= 10483725;
srom_1(80457) <= 11034723;
srom_1(80458) <= 11573312;
srom_1(80459) <= 12096968;
srom_1(80460) <= 12603233;
srom_1(80461) <= 13089735;
srom_1(80462) <= 13554192;
srom_1(80463) <= 13994425;
srom_1(80464) <= 14408371;
srom_1(80465) <= 14794088;
srom_1(80466) <= 15149767;
srom_1(80467) <= 15473741;
srom_1(80468) <= 15764491;
srom_1(80469) <= 16020652;
srom_1(80470) <= 16241024;
srom_1(80471) <= 16424574;
srom_1(80472) <= 16570440;
srom_1(80473) <= 16677938;
srom_1(80474) <= 16746565;
srom_1(80475) <= 16775999;
srom_1(80476) <= 16766102;
srom_1(80477) <= 16716919;
srom_1(80478) <= 16628682;
srom_1(80479) <= 16501805;
srom_1(80480) <= 16336882;
srom_1(80481) <= 16134686;
srom_1(80482) <= 15896167;
srom_1(80483) <= 15622442;
srom_1(80484) <= 15314796;
srom_1(80485) <= 14974670;
srom_1(80486) <= 14603659;
srom_1(80487) <= 14203504;
srom_1(80488) <= 13776082;
srom_1(80489) <= 13323395;
srom_1(80490) <= 12847567;
srom_1(80491) <= 12350830;
srom_1(80492) <= 11835513;
srom_1(80493) <= 11304032;
srom_1(80494) <= 10758879;
srom_1(80495) <= 10202612;
srom_1(80496) <= 9637838;
srom_1(80497) <= 9067206;
srom_1(80498) <= 8493391;
srom_1(80499) <= 7919086;
srom_1(80500) <= 7346982;
srom_1(80501) <= 6779762;
srom_1(80502) <= 6220087;
srom_1(80503) <= 5670581;
srom_1(80504) <= 5133821;
srom_1(80505) <= 4612324;
srom_1(80506) <= 4108535;
srom_1(80507) <= 3624816;
srom_1(80508) <= 3163437;
srom_1(80509) <= 2726560;
srom_1(80510) <= 2316234;
srom_1(80511) <= 1934384;
srom_1(80512) <= 1582800;
srom_1(80513) <= 1263131;
srom_1(80514) <= 976876;
srom_1(80515) <= 725376;
srom_1(80516) <= 509813;
srom_1(80517) <= 331195;
srom_1(80518) <= 190362;
srom_1(80519) <= 87973;
srom_1(80520) <= 24508;
srom_1(80521) <= 266;
srom_1(80522) <= 15359;
srom_1(80523) <= 69718;
srom_1(80524) <= 163086;
srom_1(80525) <= 295027;
srom_1(80526) <= 464922;
srom_1(80527) <= 671973;
srom_1(80528) <= 915210;
srom_1(80529) <= 1193493;
srom_1(80530) <= 1505516;
srom_1(80531) <= 1849816;
srom_1(80532) <= 2224779;
srom_1(80533) <= 2628646;
srom_1(80534) <= 3059523;
srom_1(80535) <= 3515391;
srom_1(80536) <= 3994110;
srom_1(80537) <= 4493437;
srom_1(80538) <= 5011030;
srom_1(80539) <= 5544461;
srom_1(80540) <= 6091230;
srom_1(80541) <= 6648771;
srom_1(80542) <= 7214472;
srom_1(80543) <= 7785678;
srom_1(80544) <= 8359712;
srom_1(80545) <= 8933881;
srom_1(80546) <= 9505493;
srom_1(80547) <= 10071868;
srom_1(80548) <= 10630349;
srom_1(80549) <= 11178318;
srom_1(80550) <= 11713205;
srom_1(80551) <= 12232502;
srom_1(80552) <= 12733773;
srom_1(80553) <= 13214669;
srom_1(80554) <= 13672933;
srom_1(80555) <= 14106418;
srom_1(80556) <= 14513090;
srom_1(80557) <= 14891041;
srom_1(80558) <= 15238501;
srom_1(80559) <= 15553839;
srom_1(80560) <= 15835577;
srom_1(80561) <= 16082394;
srom_1(80562) <= 16293132;
srom_1(80563) <= 16466802;
srom_1(80564) <= 16602592;
srom_1(80565) <= 16699863;
srom_1(80566) <= 16758160;
srom_1(80567) <= 16777209;
srom_1(80568) <= 16756921;
srom_1(80569) <= 16697391;
srom_1(80570) <= 16598898;
srom_1(80571) <= 16461905;
srom_1(80572) <= 16287053;
srom_1(80573) <= 16075162;
srom_1(80574) <= 15827227;
srom_1(80575) <= 15544409;
srom_1(80576) <= 15228035;
srom_1(80577) <= 14879589;
srom_1(80578) <= 14500705;
srom_1(80579) <= 14093158;
srom_1(80580) <= 13658862;
srom_1(80581) <= 13199851;
srom_1(80582) <= 12718278;
srom_1(80583) <= 12216402;
srom_1(80584) <= 11696577;
srom_1(80585) <= 11161239;
srom_1(80586) <= 10612899;
srom_1(80587) <= 10054129;
srom_1(80588) <= 9487549;
srom_1(80589) <= 8915815;
srom_1(80590) <= 8341609;
srom_1(80591) <= 7767623;
srom_1(80592) <= 7196550;
srom_1(80593) <= 6631066;
srom_1(80594) <= 6073824;
srom_1(80595) <= 5527437;
srom_1(80596) <= 4994467;
srom_1(80597) <= 4477413;
srom_1(80598) <= 3978701;
srom_1(80599) <= 3500667;
srom_1(80600) <= 3045555;
srom_1(80601) <= 2615498;
srom_1(80602) <= 2212514;
srom_1(80603) <= 1838491;
srom_1(80604) <= 1495184;
srom_1(80605) <= 1184203;
srom_1(80606) <= 907005;
srom_1(80607) <= 664892;
srom_1(80608) <= 458997;
srom_1(80609) <= 290287;
srom_1(80610) <= 159553;
srom_1(80611) <= 67408;
srom_1(80612) <= 14284;
srom_1(80613) <= 430;
srom_1(80614) <= 25910;
srom_1(80615) <= 90607;
srom_1(80616) <= 194216;
srom_1(80617) <= 336250;
srom_1(80618) <= 516046;
srom_1(80619) <= 732758;
srom_1(80620) <= 985371;
srom_1(80621) <= 1272701;
srom_1(80622) <= 1593399;
srom_1(80623) <= 1945963;
srom_1(80624) <= 2328738;
srom_1(80625) <= 2739930;
srom_1(80626) <= 3177611;
srom_1(80627) <= 3639728;
srom_1(80628) <= 4124114;
srom_1(80629) <= 4628497;
srom_1(80630) <= 5150513;
srom_1(80631) <= 5687714;
srom_1(80632) <= 6237580;
srom_1(80633) <= 6797533;
srom_1(80634) <= 7364947;
srom_1(80635) <= 7937161;
srom_1(80636) <= 8511493;
srom_1(80637) <= 9085248;
srom_1(80638) <= 9655736;
srom_1(80639) <= 10220282;
srom_1(80640) <= 10776239;
srom_1(80641) <= 11320999;
srom_1(80642) <= 11852009;
srom_1(80643) <= 12366777;
srom_1(80644) <= 12862891;
srom_1(80645) <= 13338023;
srom_1(80646) <= 13789945;
srom_1(80647) <= 14216539;
srom_1(80648) <= 14615803;
srom_1(80649) <= 14985866;
srom_1(80650) <= 15324992;
srom_1(80651) <= 15631592;
srom_1(80652) <= 15904226;
srom_1(80653) <= 16141617;
srom_1(80654) <= 16342651;
srom_1(80655) <= 16506386;
srom_1(80656) <= 16632054;
srom_1(80657) <= 16719066;
srom_1(80658) <= 16767014;
srom_1(80659) <= 16775672;
srom_1(80660) <= 16745000;
srom_1(80661) <= 16675142;
srom_1(80662) <= 16566426;
srom_1(80663) <= 16419361;
srom_1(80664) <= 16234638;
srom_1(80665) <= 16013121;
srom_1(80666) <= 15755851;
srom_1(80667) <= 15464033;
srom_1(80668) <= 15139036;
srom_1(80669) <= 14782384;
srom_1(80670) <= 14395749;
srom_1(80671) <= 13980945;
srom_1(80672) <= 13539916;
srom_1(80673) <= 13074731;
srom_1(80674) <= 12587571;
srom_1(80675) <= 12080721;
srom_1(80676) <= 11556557;
srom_1(80677) <= 11017538;
srom_1(80678) <= 10466191;
srom_1(80679) <= 9905101;
srom_1(80680) <= 9336900;
srom_1(80681) <= 8764251;
srom_1(80682) <= 8189842;
srom_1(80683) <= 7616364;
srom_1(80684) <= 7046508;
srom_1(80685) <= 6482945;
srom_1(80686) <= 5928319;
srom_1(80687) <= 5385230;
srom_1(80688) <= 4856224;
srom_1(80689) <= 4343784;
srom_1(80690) <= 3850310;
srom_1(80691) <= 3378119;
srom_1(80692) <= 2929423;
srom_1(80693) <= 2506327;
srom_1(80694) <= 2110815;
srom_1(80695) <= 1744742;
srom_1(80696) <= 1409825;
srom_1(80697) <= 1107633;
srom_1(80698) <= 839584;
srom_1(80699) <= 606936;
srom_1(80700) <= 410778;
srom_1(80701) <= 252031;
srom_1(80702) <= 131439;
srom_1(80703) <= 49568;
srom_1(80704) <= 6801;
srom_1(80705) <= 3340;
srom_1(80706) <= 39200;
srom_1(80707) <= 114213;
srom_1(80708) <= 228028;
srom_1(80709) <= 380110;
srom_1(80710) <= 569747;
srom_1(80711) <= 796049;
srom_1(80712) <= 1057956;
srom_1(80713) <= 1354238;
srom_1(80714) <= 1683507;
srom_1(80715) <= 2044219;
srom_1(80716) <= 2434681;
srom_1(80717) <= 2853064;
srom_1(80718) <= 3297404;
srom_1(80719) <= 3765619;
srom_1(80720) <= 4255513;
srom_1(80721) <= 4764788;
srom_1(80722) <= 5291057;
srom_1(80723) <= 5831851;
srom_1(80724) <= 6384635;
srom_1(80725) <= 6946815;
srom_1(80726) <= 7515757;
srom_1(80727) <= 8088792;
srom_1(80728) <= 8663233;
srom_1(80729) <= 9236386;
srom_1(80730) <= 9805564;
srom_1(80731) <= 10368097;
srom_1(80732) <= 10921348;
srom_1(80733) <= 11462721;
srom_1(80734) <= 11989679;
srom_1(80735) <= 12499750;
srom_1(80736) <= 12990543;
srom_1(80737) <= 13459756;
srom_1(80738) <= 13905188;
srom_1(80739) <= 14324751;
srom_1(80740) <= 14716478;
srom_1(80741) <= 15078531;
srom_1(80742) <= 15409213;
srom_1(80743) <= 15706972;
srom_1(80744) <= 15970414;
srom_1(80745) <= 16198301;
srom_1(80746) <= 16389566;
srom_1(80747) <= 16543312;
srom_1(80748) <= 16658818;
srom_1(80749) <= 16735542;
srom_1(80750) <= 16773124;
srom_1(80751) <= 16771389;
srom_1(80752) <= 16730343;
srom_1(80753) <= 16650181;
srom_1(80754) <= 16531277;
srom_1(80755) <= 16374189;
srom_1(80756) <= 16179654;
srom_1(80757) <= 15948584;
srom_1(80758) <= 15682063;
srom_1(80759) <= 15381341;
srom_1(80760) <= 15047827;
srom_1(80761) <= 14683085;
srom_1(80762) <= 14288827;
srom_1(80763) <= 13866900;
srom_1(80764) <= 13419284;
srom_1(80765) <= 12948078;
srom_1(80766) <= 12455490;
srom_1(80767) <= 11943831;
srom_1(80768) <= 11415501;
srom_1(80769) <= 10872977;
srom_1(80770) <= 10318802;
srom_1(80771) <= 9755576;
srom_1(80772) <= 9185940;
srom_1(80773) <= 8612565;
srom_1(80774) <= 8038140;
srom_1(80775) <= 7465358;
srom_1(80776) <= 6896906;
srom_1(80777) <= 6335448;
srom_1(80778) <= 5783619;
srom_1(80779) <= 5244006;
srom_1(80780) <= 4719138;
srom_1(80781) <= 4211478;
srom_1(80782) <= 3723406;
srom_1(80783) <= 3257211;
srom_1(80784) <= 2815078;
srom_1(80785) <= 2399082;
srom_1(80786) <= 2011172;
srom_1(80787) <= 1653169;
srom_1(80788) <= 1326750;
srom_1(80789) <= 1033447;
srom_1(80790) <= 774635;
srom_1(80791) <= 551527;
srom_1(80792) <= 365170;
srom_1(80793) <= 216438;
srom_1(80794) <= 106028;
srom_1(80795) <= 34457;
srom_1(80796) <= 2062;
srom_1(80797) <= 8995;
srom_1(80798) <= 55222;
srom_1(80799) <= 140528;
srom_1(80800) <= 264511;
srom_1(80801) <= 426591;
srom_1(80802) <= 626008;
srom_1(80803) <= 861827;
srom_1(80804) <= 1132941;
srom_1(80805) <= 1438079;
srom_1(80806) <= 1775811;
srom_1(80807) <= 2144552;
srom_1(80808) <= 2542574;
srom_1(80809) <= 2968010;
srom_1(80810) <= 3418865;
srom_1(80811) <= 3893025;
srom_1(80812) <= 4388266;
srom_1(80813) <= 4902266;
srom_1(80814) <= 5432615;
srom_1(80815) <= 5976825;
srom_1(80816) <= 6532345;
srom_1(80817) <= 7096570;
srom_1(80818) <= 7666854;
srom_1(80819) <= 8240522;
srom_1(80820) <= 8814884;
srom_1(80821) <= 9387248;
srom_1(80822) <= 9954928;
srom_1(80823) <= 10515264;
srom_1(80824) <= 11065627;
srom_1(80825) <= 11603436;
srom_1(80826) <= 12126170;
srom_1(80827) <= 12631378;
srom_1(80828) <= 13116689;
srom_1(80829) <= 13579829;
srom_1(80830) <= 14018625;
srom_1(80831) <= 14431021;
srom_1(80832) <= 14815081;
srom_1(80833) <= 15169006;
srom_1(80834) <= 15491135;
srom_1(80835) <= 15779957;
srom_1(80836) <= 16034119;
srom_1(80837) <= 16252429;
srom_1(80838) <= 16433862;
srom_1(80839) <= 16577569;
srom_1(80840) <= 16682875;
srom_1(80841) <= 16749286;
srom_1(80842) <= 16776490;
srom_1(80843) <= 16764362;
srom_1(80844) <= 16712956;
srom_1(80845) <= 16622515;
srom_1(80846) <= 16493462;
srom_1(80847) <= 16326402;
srom_1(80848) <= 16122120;
srom_1(80849) <= 15881572;
srom_1(80850) <= 15605888;
srom_1(80851) <= 15296359;
srom_1(80852) <= 14954437;
srom_1(80853) <= 14581726;
srom_1(80854) <= 14179973;
srom_1(80855) <= 13751062;
srom_1(80856) <= 13297005;
srom_1(80857) <= 12819931;
srom_1(80858) <= 12322077;
srom_1(80859) <= 11805777;
srom_1(80860) <= 11273454;
srom_1(80861) <= 10727602;
srom_1(80862) <= 10170781;
srom_1(80863) <= 9605604;
srom_1(80864) <= 9034720;
srom_1(80865) <= 8460805;
srom_1(80866) <= 7886553;
srom_1(80867) <= 7314654;
srom_1(80868) <= 6747792;
srom_1(80869) <= 6188624;
srom_1(80870) <= 5639772;
srom_1(80871) <= 5103811;
srom_1(80872) <= 4583253;
srom_1(80873) <= 4080540;
srom_1(80874) <= 3598029;
srom_1(80875) <= 3137982;
srom_1(80876) <= 2702558;
srom_1(80877) <= 2293797;
srom_1(80878) <= 1913617;
srom_1(80879) <= 1563801;
srom_1(80880) <= 1245988;
srom_1(80881) <= 961669;
srom_1(80882) <= 712178;
srom_1(80883) <= 498685;
srom_1(80884) <= 322190;
srom_1(80885) <= 183521;
srom_1(80886) <= 83328;
srom_1(80887) <= 22082;
srom_1(80888) <= 69;
srom_1(80889) <= 17394;
srom_1(80890) <= 73973;
srom_1(80891) <= 169543;
srom_1(80892) <= 303655;
srom_1(80893) <= 475680;
srom_1(80894) <= 684811;
srom_1(80895) <= 930068;
srom_1(80896) <= 1210301;
srom_1(80897) <= 1524195;
srom_1(80898) <= 1870279;
srom_1(80899) <= 2246929;
srom_1(80900) <= 2652380;
srom_1(80901) <= 3084731;
srom_1(80902) <= 3541952;
srom_1(80903) <= 4021902;
srom_1(80904) <= 4522328;
srom_1(80905) <= 5040885;
srom_1(80906) <= 5575140;
srom_1(80907) <= 6122589;
srom_1(80908) <= 6680664;
srom_1(80909) <= 7246748;
srom_1(80910) <= 7818186;
srom_1(80911) <= 8392299;
srom_1(80912) <= 8966395;
srom_1(80913) <= 9537782;
srom_1(80914) <= 10103780;
srom_1(80915) <= 10661734;
srom_1(80916) <= 11209030;
srom_1(80917) <= 11743099;
srom_1(80918) <= 12261438;
srom_1(80919) <= 12761616;
srom_1(80920) <= 13241287;
srom_1(80921) <= 13698203;
srom_1(80922) <= 14130219;
srom_1(80923) <= 14535312;
srom_1(80924) <= 14911581;
srom_1(80925) <= 15257261;
srom_1(80926) <= 15570731;
srom_1(80927) <= 15850522;
srom_1(80928) <= 16095322;
srom_1(80929) <= 16303982;
srom_1(80930) <= 16475524;
srom_1(80931) <= 16609144;
srom_1(80932) <= 16704215;
srom_1(80933) <= 16760292;
srom_1(80934) <= 16777110;
srom_1(80935) <= 16754592;
srom_1(80936) <= 16692843;
srom_1(80937) <= 16592153;
srom_1(80938) <= 16452993;
srom_1(80939) <= 16276017;
srom_1(80940) <= 16062054;
srom_1(80941) <= 15812107;
srom_1(80942) <= 15527349;
srom_1(80943) <= 15209115;
srom_1(80944) <= 14858898;
srom_1(80945) <= 14478339;
srom_1(80946) <= 14069223;
srom_1(80947) <= 13633469;
srom_1(80948) <= 13173119;
srom_1(80949) <= 12690334;
srom_1(80950) <= 12187376;
srom_1(80951) <= 11666605;
srom_1(80952) <= 11130462;
srom_1(80953) <= 10581461;
srom_1(80954) <= 10022177;
srom_1(80955) <= 9455233;
srom_1(80956) <= 8883288;
srom_1(80957) <= 8309022;
srom_1(80958) <= 7735130;
srom_1(80959) <= 7164302;
srom_1(80960) <= 6599215;
srom_1(80961) <= 6042519;
srom_1(80962) <= 5496825;
srom_1(80963) <= 4964692;
srom_1(80964) <= 4448614;
srom_1(80965) <= 3951012;
srom_1(80966) <= 3474220;
srom_1(80967) <= 3020473;
srom_1(80968) <= 2591899;
srom_1(80969) <= 2190508;
srom_1(80970) <= 1818182;
srom_1(80971) <= 1476667;
srom_1(80972) <= 1167564;
srom_1(80973) <= 892323;
srom_1(80974) <= 652235;
srom_1(80975) <= 448425;
srom_1(80976) <= 281850;
srom_1(80977) <= 153290;
srom_1(80978) <= 63348;
srom_1(80979) <= 12446;
srom_1(80980) <= 823;
srom_1(80981) <= 28533;
srom_1(80982) <= 95446;
srom_1(80983) <= 201249;
srom_1(80984) <= 345445;
srom_1(80985) <= 527358;
srom_1(80986) <= 746136;
srom_1(80987) <= 1000751;
srom_1(80988) <= 1290011;
srom_1(80989) <= 1612559;
srom_1(80990) <= 1966881;
srom_1(80991) <= 2351318;
srom_1(80992) <= 2764065;
srom_1(80993) <= 3203188;
srom_1(80994) <= 3666627;
srom_1(80995) <= 4152208;
srom_1(80996) <= 4657656;
srom_1(80997) <= 5180600;
srom_1(80998) <= 5718587;
srom_1(80999) <= 6269094;
srom_1(81000) <= 6829541;
srom_1(81001) <= 7397299;
srom_1(81002) <= 7969705;
srom_1(81003) <= 8544076;
srom_1(81004) <= 9117718;
srom_1(81005) <= 9687940;
srom_1(81006) <= 10252070;
srom_1(81007) <= 10807461;
srom_1(81008) <= 11351509;
srom_1(81009) <= 11881663;
srom_1(81010) <= 12395438;
srom_1(81011) <= 12890422;
srom_1(81012) <= 13364296;
srom_1(81013) <= 13814838;
srom_1(81014) <= 14239934;
srom_1(81015) <= 14637591;
srom_1(81016) <= 15005944;
srom_1(81017) <= 15343267;
srom_1(81018) <= 15647976;
srom_1(81019) <= 15918644;
srom_1(81020) <= 16154001;
srom_1(81021) <= 16352944;
srom_1(81022) <= 16514539;
srom_1(81023) <= 16638028;
srom_1(81024) <= 16722834;
srom_1(81025) <= 16768557;
srom_1(81026) <= 16774984;
srom_1(81027) <= 16742084;
srom_1(81028) <= 16670012;
srom_1(81029) <= 16559105;
srom_1(81030) <= 16409884;
srom_1(81031) <= 16223049;
srom_1(81032) <= 15999475;
srom_1(81033) <= 15740211;
srom_1(81034) <= 15446474;
srom_1(81035) <= 15119639;
srom_1(81036) <= 14761240;
srom_1(81037) <= 14372958;
srom_1(81038) <= 13956613;
srom_1(81039) <= 13514158;
srom_1(81040) <= 13047667;
srom_1(81041) <= 12559328;
srom_1(81042) <= 12051432;
srom_1(81043) <= 11526359;
srom_1(81044) <= 10986572;
srom_1(81045) <= 10434603;
srom_1(81046) <= 9873039;
srom_1(81047) <= 9304514;
srom_1(81048) <= 8731694;
srom_1(81049) <= 8157265;
srom_1(81050) <= 7583921;
srom_1(81051) <= 7014350;
srom_1(81052) <= 6451224;
srom_1(81053) <= 5897183;
srom_1(81054) <= 5354825;
srom_1(81055) <= 4826693;
srom_1(81056) <= 4315265;
srom_1(81057) <= 3822938;
srom_1(81058) <= 3352020;
srom_1(81059) <= 2904721;
srom_1(81060) <= 2483138;
srom_1(81061) <= 2089248;
srom_1(81062) <= 1724898;
srom_1(81063) <= 1391795;
srom_1(81064) <= 1091504;
srom_1(81065) <= 825431;
srom_1(81066) <= 594824;
srom_1(81067) <= 400765;
srom_1(81068) <= 244164;
srom_1(81069) <= 125755;
srom_1(81070) <= 46093;
srom_1(81071) <= 5552;
srom_1(81072) <= 4322;
srom_1(81073) <= 42409;
srom_1(81074) <= 119634;
srom_1(81075) <= 235636;
srom_1(81076) <= 389869;
srom_1(81077) <= 581611;
srom_1(81078) <= 809963;
srom_1(81079) <= 1073853;
srom_1(81080) <= 1372045;
srom_1(81081) <= 1703141;
srom_1(81082) <= 2065586;
srom_1(81083) <= 2457682;
srom_1(81084) <= 2877591;
srom_1(81085) <= 3323342;
srom_1(81086) <= 3792847;
srom_1(81087) <= 4283902;
srom_1(81088) <= 4794206;
srom_1(81089) <= 5321365;
srom_1(81090) <= 5862908;
srom_1(81091) <= 6416294;
srom_1(81092) <= 6978929;
srom_1(81093) <= 7548175;
srom_1(81094) <= 8121362;
srom_1(81095) <= 8695802;
srom_1(81096) <= 9268801;
srom_1(81097) <= 9837673;
srom_1(81098) <= 10399750;
srom_1(81099) <= 10952395;
srom_1(81100) <= 11493019;
srom_1(81101) <= 12019084;
srom_1(81102) <= 12528125;
srom_1(81103) <= 13017755;
srom_1(81104) <= 13485677;
srom_1(81105) <= 13929696;
srom_1(81106) <= 14347732;
srom_1(81107) <= 14737824;
srom_1(81108) <= 15098141;
srom_1(81109) <= 15426996;
srom_1(81110) <= 15722845;
srom_1(81111) <= 15984301;
srom_1(81112) <= 16210138;
srom_1(81113) <= 16399298;
srom_1(81114) <= 16550893;
srom_1(81115) <= 16664212;
srom_1(81116) <= 16738723;
srom_1(81117) <= 16774079;
srom_1(81118) <= 16770111;
srom_1(81119) <= 16726840;
srom_1(81120) <= 16644469;
srom_1(81121) <= 16523382;
srom_1(81122) <= 16364149;
srom_1(81123) <= 16167516;
srom_1(81124) <= 15934405;
srom_1(81125) <= 15665909;
srom_1(81126) <= 15363287;
srom_1(81127) <= 15027959;
srom_1(81128) <= 14661496;
srom_1(81129) <= 14265618;
srom_1(81130) <= 13842180;
srom_1(81131) <= 13393169;
srom_1(81132) <= 12920689;
srom_1(81133) <= 12426957;
srom_1(81134) <= 11914288;
srom_1(81135) <= 11385086;
srom_1(81136) <= 10841832;
srom_1(81137) <= 10287074;
srom_1(81138) <= 9723414;
srom_1(81139) <= 9153494;
srom_1(81140) <= 8579987;
srom_1(81141) <= 8005583;
srom_1(81142) <= 7432975;
srom_1(81143) <= 6864849;
srom_1(81144) <= 6303867;
srom_1(81145) <= 5752662;
srom_1(81146) <= 5213818;
srom_1(81147) <= 4689861;
srom_1(81148) <= 4183249;
srom_1(81149) <= 3696358;
srom_1(81150) <= 3231470;
srom_1(81151) <= 2790765;
srom_1(81152) <= 2376311;
srom_1(81153) <= 1990050;
srom_1(81154) <= 1633795;
srom_1(81155) <= 1309215;
srom_1(81156) <= 1017833;
srom_1(81157) <= 761015;
srom_1(81158) <= 539965;
srom_1(81159) <= 355720;
srom_1(81160) <= 209145;
srom_1(81161) <= 100925;
srom_1(81162) <= 31570;
srom_1(81163) <= 1403;
srom_1(81164) <= 10567;
srom_1(81165) <= 59018;
srom_1(81166) <= 146530;
srom_1(81167) <= 272691;
srom_1(81168) <= 436911;
srom_1(81169) <= 638419;
srom_1(81170) <= 876271;
srom_1(81171) <= 1149350;
srom_1(81172) <= 1456377;
srom_1(81173) <= 1795911;
srom_1(81174) <= 2166361;
srom_1(81175) <= 2565989;
srom_1(81176) <= 2992921;
srom_1(81177) <= 3445156;
srom_1(81178) <= 3920572;
srom_1(81179) <= 4416940;
srom_1(81180) <= 4931932;
srom_1(81181) <= 5463135;
srom_1(81182) <= 6008055;
srom_1(81183) <= 6564139;
srom_1(81184) <= 7128779;
srom_1(81185) <= 7699326;
srom_1(81186) <= 8273105;
srom_1(81187) <= 8847427;
srom_1(81188) <= 9419596;
srom_1(81189) <= 9986931;
srom_1(81190) <= 10546771;
srom_1(81191) <= 11096490;
srom_1(81192) <= 11633512;
srom_1(81193) <= 12155317;
srom_1(81194) <= 12659458;
srom_1(81195) <= 13143572;
srom_1(81196) <= 13605388;
srom_1(81197) <= 14042741;
srom_1(81198) <= 14453580;
srom_1(81199) <= 14835978;
srom_1(81200) <= 15188142;
srom_1(81201) <= 15508421;
srom_1(81202) <= 15795312;
srom_1(81203) <= 16047471;
srom_1(81204) <= 16263715;
srom_1(81205) <= 16443030;
srom_1(81206) <= 16584574;
srom_1(81207) <= 16687686;
srom_1(81208) <= 16751879;
srom_1(81209) <= 16776855;
srom_1(81210) <= 16762495;
srom_1(81211) <= 16708867;
srom_1(81212) <= 16616223;
srom_1(81213) <= 16484996;
srom_1(81214) <= 16315803;
srom_1(81215) <= 16109437;
srom_1(81216) <= 15866864;
srom_1(81217) <= 15589224;
srom_1(81218) <= 15277818;
srom_1(81219) <= 14934105;
srom_1(81220) <= 14559699;
srom_1(81221) <= 14156354;
srom_1(81222) <= 13725962;
srom_1(81223) <= 13270541;
srom_1(81224) <= 12792228;
srom_1(81225) <= 12293264;
srom_1(81226) <= 11775990;
srom_1(81227) <= 11242832;
srom_1(81228) <= 10696289;
srom_1(81229) <= 10138924;
srom_1(81230) <= 9573352;
srom_1(81231) <= 9002224;
srom_1(81232) <= 8428218;
srom_1(81233) <= 7854027;
srom_1(81234) <= 7282343;
srom_1(81235) <= 6715846;
srom_1(81236) <= 6157193;
srom_1(81237) <= 5609005;
srom_1(81238) <= 5073850;
srom_1(81239) <= 4554240;
srom_1(81240) <= 4052610;
srom_1(81241) <= 3571314;
srom_1(81242) <= 3112607;
srom_1(81243) <= 2678642;
srom_1(81244) <= 2271452;
srom_1(81245) <= 1892948;
srom_1(81246) <= 1544904;
srom_1(81247) <= 1228952;
srom_1(81248) <= 946575;
srom_1(81249) <= 699096;
srom_1(81250) <= 487676;
srom_1(81251) <= 313306;
srom_1(81252) <= 176803;
srom_1(81253) <= 78809;
srom_1(81254) <= 19782;
srom_1(81255) <= 0;
srom_1(81256) <= 19554;
srom_1(81257) <= 78354;
srom_1(81258) <= 176124;
srom_1(81259) <= 312404;
srom_1(81260) <= 486557;
srom_1(81261) <= 697765;
srom_1(81262) <= 945038;
srom_1(81263) <= 1227217;
srom_1(81264) <= 1542978;
srom_1(81265) <= 1890840;
srom_1(81266) <= 2269173;
srom_1(81267) <= 2676202;
srom_1(81268) <= 3110018;
srom_1(81269) <= 3568587;
srom_1(81270) <= 4049759;
srom_1(81271) <= 4551277;
srom_1(81272) <= 5070790;
srom_1(81273) <= 5605862;
srom_1(81274) <= 6153982;
srom_1(81275) <= 6712582;
srom_1(81276) <= 7279041;
srom_1(81277) <= 7850703;
srom_1(81278) <= 8424887;
srom_1(81279) <= 8998901;
srom_1(81280) <= 9570054;
srom_1(81281) <= 10135666;
srom_1(81282) <= 10693086;
srom_1(81283) <= 11239699;
srom_1(81284) <= 11772942;
srom_1(81285) <= 12290316;
srom_1(81286) <= 12789392;
srom_1(81287) <= 13267832;
srom_1(81288) <= 13723392;
srom_1(81289) <= 14153934;
srom_1(81290) <= 14557442;
srom_1(81291) <= 14932021;
srom_1(81292) <= 15275916;
srom_1(81293) <= 15587515;
srom_1(81294) <= 15865355;
srom_1(81295) <= 16108134;
srom_1(81296) <= 16314713;
srom_1(81297) <= 16484124;
srom_1(81298) <= 16615573;
srom_1(81299) <= 16708442;
srom_1(81300) <= 16762297;
srom_1(81301) <= 16776885;
srom_1(81302) <= 16752137;
srom_1(81303) <= 16688170;
srom_1(81304) <= 16585284;
srom_1(81305) <= 16443960;
srom_1(81306) <= 16264862;
srom_1(81307) <= 16048829;
srom_1(81308) <= 15796875;
srom_1(81309) <= 15510182;
srom_1(81310) <= 15190092;
srom_1(81311) <= 14838108;
srom_1(81312) <= 14455881;
srom_1(81313) <= 14045201;
srom_1(81314) <= 13607996;
srom_1(81315) <= 13146316;
srom_1(81316) <= 12662325;
srom_1(81317) <= 12158293;
srom_1(81318) <= 11636583;
srom_1(81319) <= 11099643;
srom_1(81320) <= 10549990;
srom_1(81321) <= 9990201;
srom_1(81322) <= 9422902;
srom_1(81323) <= 8850753;
srom_1(81324) <= 8276436;
srom_1(81325) <= 7702646;
srom_1(81326) <= 7132072;
srom_1(81327) <= 6567391;
srom_1(81328) <= 6011250;
srom_1(81329) <= 5466257;
srom_1(81330) <= 4934968;
srom_1(81331) <= 4419874;
srom_1(81332) <= 3923391;
srom_1(81333) <= 3447847;
srom_1(81334) <= 2995472;
srom_1(81335) <= 2568387;
srom_1(81336) <= 2168596;
srom_1(81337) <= 1797972;
srom_1(81338) <= 1458253;
srom_1(81339) <= 1151034;
srom_1(81340) <= 877754;
srom_1(81341) <= 639695;
srom_1(81342) <= 437973;
srom_1(81343) <= 273535;
srom_1(81344) <= 147150;
srom_1(81345) <= 59413;
srom_1(81346) <= 10735;
srom_1(81347) <= 1343;
srom_1(81348) <= 31282;
srom_1(81349) <= 100411;
srom_1(81350) <= 208406;
srom_1(81351) <= 354761;
srom_1(81352) <= 538790;
srom_1(81353) <= 759629;
srom_1(81354) <= 1016243;
srom_1(81355) <= 1307429;
srom_1(81356) <= 1631820;
srom_1(81357) <= 1987897;
srom_1(81358) <= 2373988;
srom_1(81359) <= 2788285;
srom_1(81360) <= 3228843;
srom_1(81361) <= 3693597;
srom_1(81362) <= 4180367;
srom_1(81363) <= 4686872;
srom_1(81364) <= 5210735;
srom_1(81365) <= 5749500;
srom_1(81366) <= 6300641;
srom_1(81367) <= 6861573;
srom_1(81368) <= 7429666;
srom_1(81369) <= 8002256;
srom_1(81370) <= 8576657;
srom_1(81371) <= 9150177;
srom_1(81372) <= 9720125;
srom_1(81373) <= 10283829;
srom_1(81374) <= 10838646;
srom_1(81375) <= 11381974;
srom_1(81376) <= 11911265;
srom_1(81377) <= 12424037;
srom_1(81378) <= 12917886;
srom_1(81379) <= 13390495;
srom_1(81380) <= 13839649;
srom_1(81381) <= 14263240;
srom_1(81382) <= 14659284;
srom_1(81383) <= 15025922;
srom_1(81384) <= 15361436;
srom_1(81385) <= 15664252;
srom_1(81386) <= 15932949;
srom_1(81387) <= 16166269;
srom_1(81388) <= 16363116;
srom_1(81389) <= 16522568;
srom_1(81390) <= 16643878;
srom_1(81391) <= 16726475;
srom_1(81392) <= 16769974;
srom_1(81393) <= 16774169;
srom_1(81394) <= 16739041;
srom_1(81395) <= 16664756;
srom_1(81396) <= 16551661;
srom_1(81397) <= 16400286;
srom_1(81398) <= 16211342;
srom_1(81399) <= 15985714;
srom_1(81400) <= 15724461;
srom_1(81401) <= 15428808;
srom_1(81402) <= 15100140;
srom_1(81403) <= 14740000;
srom_1(81404) <= 14350076;
srom_1(81405) <= 13932197;
srom_1(81406) <= 13488322;
srom_1(81407) <= 13020532;
srom_1(81408) <= 12531022;
srom_1(81409) <= 12022087;
srom_1(81410) <= 11496113;
srom_1(81411) <= 10955567;
srom_1(81412) <= 10402983;
srom_1(81413) <= 9840954;
srom_1(81414) <= 9272114;
srom_1(81415) <= 8699131;
srom_1(81416) <= 8124691;
srom_1(81417) <= 7551489;
srom_1(81418) <= 6982213;
srom_1(81419) <= 6419532;
srom_1(81420) <= 5866084;
srom_1(81421) <= 5324466;
srom_1(81422) <= 4797216;
srom_1(81423) <= 4286808;
srom_1(81424) <= 3795634;
srom_1(81425) <= 3325998;
srom_1(81426) <= 2880103;
srom_1(81427) <= 2460039;
srom_1(81428) <= 2067776;
srom_1(81429) <= 1705153;
srom_1(81430) <= 1373872;
srom_1(81431) <= 1075485;
srom_1(81432) <= 811391;
srom_1(81433) <= 582830;
srom_1(81434) <= 390873;
srom_1(81435) <= 236420;
srom_1(81436) <= 120196;
srom_1(81437) <= 42745;
srom_1(81438) <= 4430;
srom_1(81439) <= 5432;
srom_1(81440) <= 45745;
srom_1(81441) <= 125181;
srom_1(81442) <= 243367;
srom_1(81443) <= 399748;
srom_1(81444) <= 593593;
srom_1(81445) <= 823990;
srom_1(81446) <= 1089861;
srom_1(81447) <= 1389958;
srom_1(81448) <= 1722875;
srom_1(81449) <= 2087049;
srom_1(81450) <= 2480773;
srom_1(81451) <= 2902201;
srom_1(81452) <= 3349357;
srom_1(81453) <= 3820143;
srom_1(81454) <= 4312353;
srom_1(81455) <= 4823678;
srom_1(81456) <= 5351719;
srom_1(81457) <= 5894002;
srom_1(81458) <= 6447983;
srom_1(81459) <= 7011064;
srom_1(81460) <= 7580605;
srom_1(81461) <= 8153935;
srom_1(81462) <= 8728365;
srom_1(81463) <= 9301202;
srom_1(81464) <= 9869760;
srom_1(81465) <= 10431372;
srom_1(81466) <= 10983404;
srom_1(81467) <= 11523269;
srom_1(81468) <= 12048435;
srom_1(81469) <= 12556438;
srom_1(81470) <= 13044896;
srom_1(81471) <= 13511520;
srom_1(81472) <= 13954121;
srom_1(81473) <= 14370623;
srom_1(81474) <= 14759073;
srom_1(81475) <= 15117650;
srom_1(81476) <= 15444673;
srom_1(81477) <= 15738607;
srom_1(81478) <= 15998074;
srom_1(81479) <= 16221858;
srom_1(81480) <= 16408909;
srom_1(81481) <= 16558350;
srom_1(81482) <= 16669480;
srom_1(81483) <= 16741779;
srom_1(81484) <= 16774906;
srom_1(81485) <= 16768707;
srom_1(81486) <= 16723212;
srom_1(81487) <= 16638632;
srom_1(81488) <= 16515365;
srom_1(81489) <= 16353989;
srom_1(81490) <= 16155261;
srom_1(81491) <= 15920112;
srom_1(81492) <= 15649645;
srom_1(81493) <= 15345129;
srom_1(81494) <= 15007991;
srom_1(81495) <= 14639813;
srom_1(81496) <= 14242320;
srom_1(81497) <= 13817378;
srom_1(81498) <= 13366978;
srom_1(81499) <= 12893233;
srom_1(81500) <= 12398364;
srom_1(81501) <= 11884692;
srom_1(81502) <= 11354625;
srom_1(81503) <= 10810650;
srom_1(81504) <= 10255318;
srom_1(81505) <= 9691231;
srom_1(81506) <= 9121036;
srom_1(81507) <= 8547407;
srom_1(81508) <= 7973032;
srom_1(81509) <= 7400607;
srom_1(81510) <= 6832815;
srom_1(81511) <= 6272318;
srom_1(81512) <= 5721745;
srom_1(81513) <= 5183678;
srom_1(81514) <= 4660640;
srom_1(81515) <= 4155084;
srom_1(81516) <= 3669380;
srom_1(81517) <= 3205807;
srom_1(81518) <= 2766537;
srom_1(81519) <= 2353631;
srom_1(81520) <= 1969025;
srom_1(81521) <= 1614523;
srom_1(81522) <= 1291787;
srom_1(81523) <= 1002330;
srom_1(81524) <= 747510;
srom_1(81525) <= 528522;
srom_1(81526) <= 346392;
srom_1(81527) <= 201975;
srom_1(81528) <= 95948;
srom_1(81529) <= 28808;
srom_1(81530) <= 870;
srom_1(81531) <= 12265;
srom_1(81532) <= 62940;
srom_1(81533) <= 152656;
srom_1(81534) <= 280994;
srom_1(81535) <= 447351;
srom_1(81536) <= 650948;
srom_1(81537) <= 890828;
srom_1(81538) <= 1165869;
srom_1(81539) <= 1474779;
srom_1(81540) <= 1816111;
srom_1(81541) <= 2188264;
srom_1(81542) <= 2589492;
srom_1(81543) <= 3017914;
srom_1(81544) <= 3471521;
srom_1(81545) <= 3948186;
srom_1(81546) <= 4445673;
srom_1(81547) <= 4961651;
srom_1(81548) <= 5493698;
srom_1(81549) <= 6039321;
srom_1(81550) <= 6595961;
srom_1(81551) <= 7161006;
srom_1(81552) <= 7731809;
srom_1(81553) <= 8305691;
srom_1(81554) <= 8879962;
srom_1(81555) <= 9451929;
srom_1(81556) <= 10018910;
srom_1(81557) <= 10578246;
srom_1(81558) <= 11127313;
srom_1(81559) <= 11663538;
srom_1(81560) <= 12184406;
srom_1(81561) <= 12687474;
srom_1(81562) <= 13170383;
srom_1(81563) <= 13630868;
srom_1(81564) <= 14066771;
srom_1(81565) <= 14476047;
srom_1(81566) <= 14856777;
srom_1(81567) <= 15207175;
srom_1(81568) <= 15525599;
srom_1(81569) <= 15810555;
srom_1(81570) <= 16060707;
srom_1(81571) <= 16274882;
srom_1(81572) <= 16452075;
srom_1(81573) <= 16591456;
srom_1(81574) <= 16692371;
srom_1(81575) <= 16754347;
srom_1(81576) <= 16777093;
srom_1(81577) <= 16760502;
srom_1(81578) <= 16704653;
srom_1(81579) <= 16609807;
srom_1(81580) <= 16476409;
srom_1(81581) <= 16305085;
srom_1(81582) <= 16096637;
srom_1(81583) <= 15852044;
srom_1(81584) <= 15572452;
srom_1(81585) <= 15259172;
srom_1(81586) <= 14913675;
srom_1(81587) <= 14537578;
srom_1(81588) <= 14132648;
srom_1(81589) <= 13700781;
srom_1(81590) <= 13244004;
srom_1(81591) <= 12764458;
srom_1(81592) <= 12264393;
srom_1(81593) <= 11746152;
srom_1(81594) <= 11212167;
srom_1(81595) <= 10664941;
srom_1(81596) <= 10107041;
srom_1(81597) <= 9541082;
srom_1(81598) <= 8969719;
srom_1(81599) <= 8395631;
srom_1(81600) <= 7821510;
srom_1(81601) <= 7250048;
srom_1(81602) <= 6683925;
srom_1(81603) <= 6125796;
srom_1(81604) <= 5578279;
srom_1(81605) <= 5043940;
srom_1(81606) <= 4525285;
srom_1(81607) <= 4024746;
srom_1(81608) <= 3544672;
srom_1(81609) <= 3087312;
srom_1(81610) <= 2654812;
srom_1(81611) <= 2249199;
srom_1(81612) <= 1872376;
srom_1(81613) <= 1526110;
srom_1(81614) <= 1212025;
srom_1(81615) <= 931593;
srom_1(81616) <= 686130;
srom_1(81617) <= 476786;
srom_1(81618) <= 304544;
srom_1(81619) <= 170210;
srom_1(81620) <= 74415;
srom_1(81621) <= 17609;
srom_1(81622) <= 56;
srom_1(81623) <= 21841;
srom_1(81624) <= 82860;
srom_1(81625) <= 182828;
srom_1(81626) <= 321276;
srom_1(81627) <= 497554;
srom_1(81628) <= 710836;
srom_1(81629) <= 960121;
srom_1(81630) <= 1244241;
srom_1(81631) <= 1561864;
srom_1(81632) <= 1911500;
srom_1(81633) <= 2291509;
srom_1(81634) <= 2700109;
srom_1(81635) <= 3135385;
srom_1(81636) <= 3595295;
srom_1(81637) <= 4077682;
srom_1(81638) <= 4580285;
srom_1(81639) <= 5100746;
srom_1(81640) <= 5636625;
srom_1(81641) <= 6185409;
srom_1(81642) <= 6744525;
srom_1(81643) <= 7311350;
srom_1(81644) <= 7883227;
srom_1(81645) <= 8457474;
srom_1(81646) <= 9031398;
srom_1(81647) <= 9602308;
srom_1(81648) <= 10167526;
srom_1(81649) <= 10724402;
srom_1(81650) <= 11270325;
srom_1(81651) <= 11802735;
srom_1(81652) <= 12319134;
srom_1(81653) <= 12817102;
srom_1(81654) <= 13294303;
srom_1(81655) <= 13748500;
srom_1(81656) <= 14177562;
srom_1(81657) <= 14579478;
srom_1(81658) <= 14952363;
srom_1(81659) <= 15294468;
srom_1(81660) <= 15604189;
srom_1(81661) <= 15880074;
srom_1(81662) <= 16120829;
srom_1(81663) <= 16325324;
srom_1(81664) <= 16492602;
srom_1(81665) <= 16621877;
srom_1(81666) <= 16712544;
srom_1(81667) <= 16764177;
srom_1(81668) <= 16776533;
srom_1(81669) <= 16749556;
srom_1(81670) <= 16683372;
srom_1(81671) <= 16578291;
srom_1(81672) <= 16434805;
srom_1(81673) <= 16253588;
srom_1(81674) <= 16035489;
srom_1(81675) <= 15781532;
srom_1(81676) <= 15492907;
srom_1(81677) <= 15170967;
srom_1(81678) <= 14817222;
srom_1(81679) <= 14433331;
srom_1(81680) <= 14021095;
srom_1(81681) <= 13582445;
srom_1(81682) <= 13119440;
srom_1(81683) <= 12634251;
srom_1(81684) <= 12129152;
srom_1(81685) <= 11606513;
srom_1(81686) <= 11068784;
srom_1(81687) <= 10518486;
srom_1(81688) <= 9958201;
srom_1(81689) <= 9390555;
srom_1(81690) <= 8818211;
srom_1(81691) <= 8243852;
srom_1(81692) <= 7670173;
srom_1(81693) <= 7099862;
srom_1(81694) <= 6535594;
srom_1(81695) <= 5980016;
srom_1(81696) <= 5435733;
srom_1(81697) <= 4905296;
srom_1(81698) <= 4391194;
srom_1(81699) <= 3895838;
srom_1(81700) <= 3421549;
srom_1(81701) <= 2970553;
srom_1(81702) <= 2544963;
srom_1(81703) <= 2146777;
srom_1(81704) <= 1777861;
srom_1(81705) <= 1439945;
srom_1(81706) <= 1134613;
srom_1(81707) <= 863298;
srom_1(81708) <= 627272;
srom_1(81709) <= 427641;
srom_1(81710) <= 265342;
srom_1(81711) <= 141136;
srom_1(81712) <= 55604;
srom_1(81713) <= 9150;
srom_1(81714) <= 1989;
srom_1(81715) <= 34156;
srom_1(81716) <= 105500;
srom_1(81717) <= 215687;
srom_1(81718) <= 364199;
srom_1(81719) <= 550340;
srom_1(81720) <= 773237;
srom_1(81721) <= 1031846;
srom_1(81722) <= 1324953;
srom_1(81723) <= 1651184;
srom_1(81724) <= 2009009;
srom_1(81725) <= 2396750;
srom_1(81726) <= 2812589;
srom_1(81727) <= 3254576;
srom_1(81728) <= 3720638;
srom_1(81729) <= 4208589;
srom_1(81730) <= 4716143;
srom_1(81731) <= 5240918;
srom_1(81732) <= 5780453;
srom_1(81733) <= 6332219;
srom_1(81734) <= 6893628;
srom_1(81735) <= 7462047;
srom_1(81736) <= 8034812;
srom_1(81737) <= 8609235;
srom_1(81738) <= 9182624;
srom_1(81739) <= 9752289;
srom_1(81740) <= 10315560;
srom_1(81741) <= 10869795;
srom_1(81742) <= 11412394;
srom_1(81743) <= 11940814;
srom_1(81744) <= 12452576;
srom_1(81745) <= 12945281;
srom_1(81746) <= 13416618;
srom_1(81747) <= 13864377;
srom_1(81748) <= 14286458;
srom_1(81749) <= 14680883;
srom_1(81750) <= 15045800;
srom_1(81751) <= 15379500;
srom_1(81752) <= 15680417;
srom_1(81753) <= 15947140;
srom_1(81754) <= 16178419;
srom_1(81755) <= 16373168;
srom_1(81756) <= 16530476;
srom_1(81757) <= 16649603;
srom_1(81758) <= 16729991;
srom_1(81759) <= 16771264;
srom_1(81760) <= 16773228;
srom_1(81761) <= 16735873;
srom_1(81762) <= 16659375;
srom_1(81763) <= 16544093;
srom_1(81764) <= 16390567;
srom_1(81765) <= 16199517;
srom_1(81766) <= 15971839;
srom_1(81767) <= 15708600;
srom_1(81768) <= 15411035;
srom_1(81769) <= 15080540;
srom_1(81770) <= 14718664;
srom_1(81771) <= 14327105;
srom_1(81772) <= 13907697;
srom_1(81773) <= 13462409;
srom_1(81774) <= 12993328;
srom_1(81775) <= 12502654;
srom_1(81776) <= 11992688;
srom_1(81777) <= 11465820;
srom_1(81778) <= 10924523;
srom_1(81779) <= 10371334;
srom_1(81780) <= 9808847;
srom_1(81781) <= 9239701;
srom_1(81782) <= 8666563;
srom_1(81783) <= 8092122;
srom_1(81784) <= 7519071;
srom_1(81785) <= 6950097;
srom_1(81786) <= 6387870;
srom_1(81787) <= 5835024;
srom_1(81788) <= 5294153;
srom_1(81789) <= 4767793;
srom_1(81790) <= 4258412;
srom_1(81791) <= 3768400;
srom_1(81792) <= 3300052;
srom_1(81793) <= 2855567;
srom_1(81794) <= 2437028;
srom_1(81795) <= 2046399;
srom_1(81796) <= 1685510;
srom_1(81797) <= 1356054;
srom_1(81798) <= 1059576;
srom_1(81799) <= 797466;
srom_1(81800) <= 570954;
srom_1(81801) <= 381102;
srom_1(81802) <= 228800;
srom_1(81803) <= 114761;
srom_1(81804) <= 39522;
srom_1(81805) <= 3434;
srom_1(81806) <= 6668;
srom_1(81807) <= 49207;
srom_1(81808) <= 130852;
srom_1(81809) <= 251221;
srom_1(81810) <= 409749;
srom_1(81811) <= 605692;
srom_1(81812) <= 838132;
srom_1(81813) <= 1105979;
srom_1(81814) <= 1407977;
srom_1(81815) <= 1742709;
srom_1(81816) <= 2108606;
srom_1(81817) <= 2503953;
srom_1(81818) <= 2926894;
srom_1(81819) <= 3375447;
srom_1(81820) <= 3847509;
srom_1(81821) <= 4340865;
srom_1(81822) <= 4853203;
srom_1(81823) <= 5382120;
srom_1(81824) <= 5925134;
srom_1(81825) <= 6479701;
srom_1(81826) <= 7043220;
srom_1(81827) <= 7613047;
srom_1(81828) <= 8186512;
srom_1(81829) <= 8760924;
srom_1(81830) <= 9333590;
srom_1(81831) <= 9901824;
srom_1(81832) <= 10462963;
srom_1(81833) <= 11014374;
srom_1(81834) <= 11553473;
srom_1(81835) <= 12077730;
srom_1(81836) <= 12584687;
srom_1(81837) <= 13071968;
srom_1(81838) <= 13537287;
srom_1(81839) <= 13978461;
srom_1(81840) <= 14393423;
srom_1(81841) <= 14780227;
srom_1(81842) <= 15137058;
srom_1(81843) <= 15462243;
srom_1(81844) <= 15754257;
srom_1(81845) <= 16011732;
srom_1(81846) <= 16233459;
srom_1(81847) <= 16418398;
srom_1(81848) <= 16565683;
srom_1(81849) <= 16674624;
srom_1(81850) <= 16744708;
srom_1(81851) <= 16775607;
srom_1(81852) <= 16767177;
srom_1(81853) <= 16719457;
srom_1(81854) <= 16632671;
srom_1(81855) <= 16507225;
srom_1(81856) <= 16343709;
srom_1(81857) <= 16142888;
srom_1(81858) <= 15905705;
srom_1(81859) <= 15633271;
srom_1(81860) <= 15326865;
srom_1(81861) <= 14987923;
srom_1(81862) <= 14618035;
srom_1(81863) <= 14218934;
srom_1(81864) <= 13792493;
srom_1(81865) <= 13340712;
srom_1(81866) <= 12865708;
srom_1(81867) <= 12369710;
srom_1(81868) <= 11855043;
srom_1(81869) <= 11324120;
srom_1(81870) <= 10779432;
srom_1(81871) <= 10223533;
srom_1(81872) <= 9659029;
srom_1(81873) <= 9088567;
srom_1(81874) <= 8514823;
srom_1(81875) <= 7940488;
srom_1(81876) <= 7368253;
srom_1(81877) <= 6800804;
srom_1(81878) <= 6240800;
srom_1(81879) <= 5690868;
srom_1(81880) <= 5153587;
srom_1(81881) <= 4631475;
srom_1(81882) <= 4126983;
srom_1(81883) <= 3642474;
srom_1(81884) <= 3180222;
srom_1(81885) <= 2742393;
srom_1(81886) <= 2331042;
srom_1(81887) <= 1948097;
srom_1(81888) <= 1595353;
srom_1(81889) <= 1274465;
srom_1(81890) <= 986938;
srom_1(81891) <= 734120;
srom_1(81892) <= 517197;
srom_1(81893) <= 337185;
srom_1(81894) <= 194929;
srom_1(81895) <= 91096;
srom_1(81896) <= 26173;
srom_1(81897) <= 464;
srom_1(81898) <= 14090;
srom_1(81899) <= 66987;
srom_1(81900) <= 158907;
srom_1(81901) <= 289419;
srom_1(81902) <= 457911;
srom_1(81903) <= 663592;
srom_1(81904) <= 905499;
srom_1(81905) <= 1182497;
srom_1(81906) <= 1493286;
srom_1(81907) <= 1836411;
srom_1(81908) <= 2210260;
srom_1(81909) <= 2613082;
srom_1(81910) <= 3042987;
srom_1(81911) <= 3497960;
srom_1(81912) <= 3975867;
srom_1(81913) <= 4474467;
srom_1(81914) <= 4991421;
srom_1(81915) <= 5524306;
srom_1(81916) <= 6070623;
srom_1(81917) <= 6627809;
srom_1(81918) <= 7193252;
srom_1(81919) <= 7764301;
srom_1(81920) <= 8338278;
srom_1(81921) <= 8912490;
srom_1(81922) <= 9484246;
srom_1(81923) <= 10050864;
srom_1(81924) <= 10609687;
srom_1(81925) <= 11158095;
srom_1(81926) <= 11693515;
srom_1(81927) <= 12213438;
srom_1(81928) <= 12715425;
srom_1(81929) <= 13197121;
srom_1(81930) <= 13656269;
srom_1(81931) <= 14090716;
srom_1(81932) <= 14498423;
srom_1(81933) <= 14877479;
srom_1(81934) <= 15226106;
srom_1(81935) <= 15542670;
srom_1(81936) <= 15825686;
srom_1(81937) <= 16073827;
srom_1(81938) <= 16285930;
srom_1(81939) <= 16460999;
srom_1(81940) <= 16598214;
srom_1(81941) <= 16696932;
srom_1(81942) <= 16756688;
srom_1(81943) <= 16777204;
srom_1(81944) <= 16758383;
srom_1(81945) <= 16700313;
srom_1(81946) <= 16603267;
srom_1(81947) <= 16467700;
srom_1(81948) <= 16294246;
srom_1(81949) <= 16083721;
srom_1(81950) <= 15837110;
srom_1(81951) <= 15555571;
srom_1(81952) <= 15240424;
srom_1(81953) <= 14893145;
srom_1(81954) <= 14515365;
srom_1(81955) <= 14108855;
srom_1(81956) <= 13675520;
srom_1(81957) <= 13217393;
srom_1(81958) <= 12736622;
srom_1(81959) <= 12235462;
srom_1(81960) <= 11716263;
srom_1(81961) <= 11181459;
srom_1(81962) <= 10633559;
srom_1(81963) <= 10075131;
srom_1(81964) <= 9508794;
srom_1(81965) <= 8937205;
srom_1(81966) <= 8363043;
srom_1(81967) <= 7789001;
srom_1(81968) <= 7217770;
srom_1(81969) <= 6652030;
srom_1(81970) <= 6094434;
srom_1(81971) <= 5547595;
srom_1(81972) <= 5014079;
srom_1(81973) <= 4496388;
srom_1(81974) <= 3996948;
srom_1(81975) <= 3518103;
srom_1(81976) <= 3062096;
srom_1(81977) <= 2631068;
srom_1(81978) <= 2227039;
srom_1(81979) <= 1851903;
srom_1(81980) <= 1507420;
srom_1(81981) <= 1195206;
srom_1(81982) <= 916724;
srom_1(81983) <= 673280;
srom_1(81984) <= 466016;
srom_1(81985) <= 295903;
srom_1(81986) <= 163741;
srom_1(81987) <= 70147;
srom_1(81988) <= 15561;
srom_1(81989) <= 240;
srom_1(81990) <= 24254;
srom_1(81991) <= 87492;
srom_1(81992) <= 189657;
srom_1(81993) <= 330269;
srom_1(81994) <= 508670;
srom_1(81995) <= 724022;
srom_1(81996) <= 975316;
srom_1(81997) <= 1261374;
srom_1(81998) <= 1580853;
srom_1(81999) <= 1932257;
srom_1(82000) <= 2313937;
srom_1(82001) <= 2724102;
srom_1(82002) <= 3160831;
srom_1(82003) <= 3622074;
srom_1(82004) <= 4105670;
srom_1(82005) <= 4609349;
srom_1(82006) <= 5130751;
srom_1(82007) <= 5667430;
srom_1(82008) <= 6216870;
srom_1(82009) <= 6776493;
srom_1(82010) <= 7343676;
srom_1(82011) <= 7915760;
srom_1(82012) <= 8490060;
srom_1(82013) <= 9063885;
srom_1(82014) <= 9634544;
srom_1(82015) <= 10199359;
srom_1(82016) <= 10755684;
srom_1(82017) <= 11300908;
srom_1(82018) <= 11832476;
srom_1(82019) <= 12347894;
srom_1(82020) <= 12844745;
srom_1(82021) <= 13320701;
srom_1(82022) <= 13773528;
srom_1(82023) <= 14201103;
srom_1(82024) <= 14601421;
srom_1(82025) <= 14972606;
srom_1(82026) <= 15312916;
srom_1(82027) <= 15620755;
srom_1(82028) <= 15894680;
srom_1(82029) <= 16133407;
srom_1(82030) <= 16335816;
srom_1(82031) <= 16500957;
srom_1(82032) <= 16628057;
srom_1(82033) <= 16716520;
srom_1(82034) <= 16765930;
srom_1(82035) <= 16776055;
srom_1(82036) <= 16746849;
srom_1(82037) <= 16678449;
srom_1(82038) <= 16571174;
srom_1(82039) <= 16425529;
srom_1(82040) <= 16242196;
srom_1(82041) <= 16022034;
srom_1(82042) <= 15766077;
srom_1(82043) <= 15475524;
srom_1(82044) <= 15151739;
srom_1(82045) <= 14796238;
srom_1(82046) <= 14410690;
srom_1(82047) <= 13996903;
srom_1(82048) <= 13556816;
srom_1(82049) <= 13092494;
srom_1(82050) <= 12606113;
srom_1(82051) <= 12099956;
srom_1(82052) <= 11576394;
srom_1(82053) <= 11037884;
srom_1(82054) <= 10486950;
srom_1(82055) <= 9926177;
srom_1(82056) <= 9358193;
srom_1(82057) <= 8785663;
srom_1(82058) <= 8211271;
srom_1(82059) <= 7637710;
srom_1(82060) <= 7067670;
srom_1(82061) <= 6503825;
srom_1(82062) <= 5948819;
srom_1(82063) <= 5405253;
srom_1(82064) <= 4875677;
srom_1(82065) <= 4362575;
srom_1(82066) <= 3868352;
srom_1(82067) <= 3395326;
srom_1(82068) <= 2945715;
srom_1(82069) <= 2521628;
srom_1(82070) <= 2125053;
srom_1(82071) <= 1757850;
srom_1(82072) <= 1421741;
srom_1(82073) <= 1118302;
srom_1(82074) <= 848956;
srom_1(82075) <= 614966;
srom_1(82076) <= 417429;
srom_1(82077) <= 257272;
srom_1(82078) <= 135245;
srom_1(82079) <= 51921;
srom_1(82080) <= 7691;
srom_1(82081) <= 2762;
srom_1(82082) <= 37157;
srom_1(82083) <= 110715;
srom_1(82084) <= 223091;
srom_1(82085) <= 373757;
srom_1(82086) <= 562008;
srom_1(82087) <= 786961;
srom_1(82088) <= 1047560;
srom_1(82089) <= 1342584;
srom_1(82090) <= 1670649;
srom_1(82091) <= 2030217;
srom_1(82092) <= 2419602;
srom_1(82093) <= 2836977;
srom_1(82094) <= 3280386;
srom_1(82095) <= 3747749;
srom_1(82096) <= 4236875;
srom_1(82097) <= 4745469;
srom_1(82098) <= 5271148;
srom_1(82099) <= 5811445;
srom_1(82100) <= 6363828;
srom_1(82101) <= 6925705;
srom_1(82102) <= 7494443;
srom_1(82103) <= 8067373;
srom_1(82104) <= 8641810;
srom_1(82105) <= 9215059;
srom_1(82106) <= 9784433;
srom_1(82107) <= 10347262;
srom_1(82108) <= 10900905;
srom_1(82109) <= 11442768;
srom_1(82110) <= 11970309;
srom_1(82111) <= 12481054;
srom_1(82112) <= 12972607;
srom_1(82113) <= 13442665;
srom_1(82114) <= 13889023;
srom_1(82115) <= 14309587;
srom_1(82116) <= 14702386;
srom_1(82117) <= 15065578;
srom_1(82118) <= 15397458;
srom_1(82119) <= 15696472;
srom_1(82120) <= 15961217;
srom_1(82121) <= 16190451;
srom_1(82122) <= 16383100;
srom_1(82123) <= 16538260;
srom_1(82124) <= 16655203;
srom_1(82125) <= 16733381;
srom_1(82126) <= 16772428;
srom_1(82127) <= 16772160;
srom_1(82128) <= 16732579;
srom_1(82129) <= 16653870;
srom_1(82130) <= 16536402;
srom_1(82131) <= 16380727;
srom_1(82132) <= 16187574;
srom_1(82133) <= 15957848;
srom_1(82134) <= 15692628;
srom_1(82135) <= 15393157;
srom_1(82136) <= 15060839;
srom_1(82137) <= 14697233;
srom_1(82138) <= 14304044;
srom_1(82139) <= 13883115;
srom_1(82140) <= 13436420;
srom_1(82141) <= 12966054;
srom_1(82142) <= 12474223;
srom_1(82143) <= 11963234;
srom_1(82144) <= 11435481;
srom_1(82145) <= 10893441;
srom_1(82146) <= 10339655;
srom_1(82147) <= 9776719;
srom_1(82148) <= 9207275;
srom_1(82149) <= 8633991;
srom_1(82150) <= 8059556;
srom_1(82151) <= 7486665;
srom_1(82152) <= 6918003;
srom_1(82153) <= 6356237;
srom_1(82154) <= 5804002;
srom_1(82155) <= 5263887;
srom_1(82156) <= 4738425;
srom_1(82157) <= 4230079;
srom_1(82158) <= 3741235;
srom_1(82159) <= 3274183;
srom_1(82160) <= 2831115;
srom_1(82161) <= 2414108;
srom_1(82162) <= 2025117;
srom_1(82163) <= 1665967;
srom_1(82164) <= 1338342;
srom_1(82165) <= 1043778;
srom_1(82166) <= 783656;
srom_1(82167) <= 559196;
srom_1(82168) <= 371452;
srom_1(82169) <= 221302;
srom_1(82170) <= 109452;
srom_1(82171) <= 36425;
srom_1(82172) <= 2565;
srom_1(82173) <= 8030;
srom_1(82174) <= 52794;
srom_1(82175) <= 136648;
srom_1(82176) <= 259198;
srom_1(82177) <= 419869;
srom_1(82178) <= 617909;
srom_1(82179) <= 852388;
srom_1(82180) <= 1122207;
srom_1(82181) <= 1426101;
srom_1(82182) <= 1762644;
srom_1(82183) <= 2130259;
srom_1(82184) <= 2527221;
srom_1(82185) <= 2951670;
srom_1(82186) <= 3401613;
srom_1(82187) <= 3874943;
srom_1(82188) <= 4369439;
srom_1(82189) <= 4882782;
srom_1(82190) <= 5412565;
srom_1(82191) <= 5956304;
srom_1(82192) <= 6511449;
srom_1(82193) <= 7075396;
srom_1(82194) <= 7645501;
srom_1(82195) <= 8219091;
srom_1(82196) <= 8793476;
srom_1(82197) <= 9365963;
srom_1(82198) <= 9933866;
srom_1(82199) <= 10494523;
srom_1(82200) <= 11045305;
srom_1(82201) <= 11583628;
srom_1(82202) <= 12106969;
srom_1(82203) <= 12612873;
srom_1(82204) <= 13098969;
srom_1(82205) <= 13562975;
srom_1(82206) <= 14002718;
srom_1(82207) <= 14416133;
srom_1(82208) <= 14801284;
srom_1(82209) <= 15156363;
srom_1(82210) <= 15479707;
srom_1(82211) <= 15769797;
srom_1(82212) <= 16025275;
srom_1(82213) <= 16244941;
srom_1(82214) <= 16427767;
srom_1(82215) <= 16572894;
srom_1(82216) <= 16679642;
srom_1(82217) <= 16747511;
srom_1(82218) <= 16776182;
srom_1(82219) <= 16765520;
srom_1(82220) <= 16715577;
srom_1(82221) <= 16626585;
srom_1(82222) <= 16498963;
srom_1(82223) <= 16333308;
srom_1(82224) <= 16130398;
srom_1(82225) <= 15891185;
srom_1(82226) <= 15616789;
srom_1(82227) <= 15308497;
srom_1(82228) <= 14967756;
srom_1(82229) <= 14596163;
srom_1(82230) <= 14195460;
srom_1(82231) <= 13767527;
srom_1(82232) <= 13314371;
srom_1(82233) <= 12838116;
srom_1(82234) <= 12340996;
srom_1(82235) <= 11825341;
srom_1(82236) <= 11293571;
srom_1(82237) <= 10748178;
srom_1(82238) <= 10191720;
srom_1(82239) <= 9626807;
srom_1(82240) <= 9056088;
srom_1(82241) <= 8482238;
srom_1(82242) <= 7907950;
srom_1(82243) <= 7335915;
srom_1(82244) <= 6768817;
srom_1(82245) <= 6209315;
srom_1(82246) <= 5660032;
srom_1(82247) <= 5123544;
srom_1(82248) <= 4602367;
srom_1(82249) <= 4098946;
srom_1(82250) <= 3615640;
srom_1(82251) <= 3154716;
srom_1(82252) <= 2718335;
srom_1(82253) <= 2308545;
srom_1(82254) <= 1927265;
srom_1(82255) <= 1576286;
srom_1(82256) <= 1257251;
srom_1(82257) <= 971658;
srom_1(82258) <= 720846;
srom_1(82259) <= 505990;
srom_1(82260) <= 328099;
srom_1(82261) <= 188006;
srom_1(82262) <= 86369;
srom_1(82263) <= 23664;
srom_1(82264) <= 184;
srom_1(82265) <= 16041;
srom_1(82266) <= 71160;
srom_1(82267) <= 165282;
srom_1(82268) <= 297966;
srom_1(82269) <= 468590;
srom_1(82270) <= 676354;
srom_1(82271) <= 920283;
srom_1(82272) <= 1199233;
srom_1(82273) <= 1511897;
srom_1(82274) <= 1856809;
srom_1(82275) <= 2232350;
srom_1(82276) <= 2636760;
srom_1(82277) <= 3068142;
srom_1(82278) <= 3524474;
srom_1(82279) <= 4003615;
srom_1(82280) <= 4503319;
srom_1(82281) <= 5021243;
srom_1(82282) <= 5554957;
srom_1(82283) <= 6101959;
srom_1(82284) <= 6659684;
srom_1(82285) <= 7225517;
srom_1(82286) <= 7796803;
srom_1(82287) <= 8370865;
srom_1(82288) <= 8945010;
srom_1(82289) <= 9516546;
srom_1(82290) <= 10082793;
srom_1(82291) <= 10641095;
srom_1(82292) <= 11188834;
srom_1(82293) <= 11723442;
srom_1(82294) <= 12242412;
srom_1(82295) <= 12743310;
srom_1(82296) <= 13223788;
srom_1(82297) <= 13681591;
srom_1(82298) <= 14114574;
srom_1(82299) <= 14520706;
srom_1(82300) <= 14898082;
srom_1(82301) <= 15244934;
srom_1(82302) <= 15559633;
srom_1(82303) <= 15840705;
srom_1(82304) <= 16086832;
srom_1(82305) <= 16296859;
srom_1(82306) <= 16469801;
srom_1(82307) <= 16604848;
srom_1(82308) <= 16701367;
srom_1(82309) <= 16758904;
srom_1(82310) <= 16777189;
srom_1(82311) <= 16756138;
srom_1(82312) <= 16695848;
srom_1(82313) <= 16596603;
srom_1(82314) <= 16458868;
srom_1(82315) <= 16283289;
srom_1(82316) <= 16070689;
srom_1(82317) <= 15822064;
srom_1(82318) <= 15538582;
srom_1(82319) <= 15221571;
srom_1(82320) <= 14872518;
srom_1(82321) <= 14493060;
srom_1(82322) <= 14084976;
srom_1(82323) <= 13650179;
srom_1(82324) <= 13190710;
srom_1(82325) <= 12708721;
srom_1(82326) <= 12206474;
srom_1(82327) <= 11686324;
srom_1(82328) <= 11150710;
srom_1(82329) <= 10602143;
srom_1(82330) <= 10043196;
srom_1(82331) <= 9476490;
srom_1(82332) <= 8904683;
srom_1(82333) <= 8330455;
srom_1(82334) <= 7756501;
srom_1(82335) <= 7185510;
srom_1(82336) <= 6620162;
srom_1(82337) <= 6063106;
srom_1(82338) <= 5516955;
srom_1(82339) <= 4984270;
srom_1(82340) <= 4467550;
srom_1(82341) <= 3969216;
srom_1(82342) <= 3491607;
srom_1(82343) <= 3036961;
srom_1(82344) <= 2607411;
srom_1(82345) <= 2204972;
srom_1(82346) <= 1831529;
srom_1(82347) <= 1488834;
srom_1(82348) <= 1178496;
srom_1(82349) <= 901967;
srom_1(82350) <= 660546;
srom_1(82351) <= 455365;
srom_1(82352) <= 287386;
srom_1(82353) <= 157395;
srom_1(82354) <= 66004;
srom_1(82355) <= 13641;
srom_1(82356) <= 550;
srom_1(82357) <= 26794;
srom_1(82358) <= 92249;
srom_1(82359) <= 196609;
srom_1(82360) <= 339384;
srom_1(82361) <= 519904;
srom_1(82362) <= 737324;
srom_1(82363) <= 990623;
srom_1(82364) <= 1278613;
srom_1(82365) <= 1599945;
srom_1(82366) <= 1953112;
srom_1(82367) <= 2336456;
srom_1(82368) <= 2748181;
srom_1(82369) <= 3186356;
srom_1(82370) <= 3648926;
srom_1(82371) <= 4133722;
srom_1(82372) <= 4638471;
srom_1(82373) <= 5160806;
srom_1(82374) <= 5698276;
srom_1(82375) <= 6248363;
srom_1(82376) <= 6808486;
srom_1(82377) <= 7376018;
srom_1(82378) <= 7948299;
srom_1(82379) <= 8522645;
srom_1(82380) <= 9096362;
srom_1(82381) <= 9666761;
srom_1(82382) <= 10231165;
srom_1(82383) <= 10786929;
srom_1(82384) <= 11331447;
srom_1(82385) <= 11862165;
srom_1(82386) <= 12376594;
srom_1(82387) <= 12872321;
srom_1(82388) <= 13347024;
srom_1(82389) <= 13798474;
srom_1(82390) <= 14224556;
srom_1(82391) <= 14623271;
srom_1(82392) <= 14992749;
srom_1(82393) <= 15331259;
srom_1(82394) <= 15637212;
srom_1(82395) <= 15909174;
srom_1(82396) <= 16145869;
srom_1(82397) <= 16346187;
srom_1(82398) <= 16509190;
srom_1(82399) <= 16634113;
srom_1(82400) <= 16720370;
srom_1(82401) <= 16767556;
srom_1(82402) <= 16775450;
srom_1(82403) <= 16744016;
srom_1(82404) <= 16673400;
srom_1(82405) <= 16563934;
srom_1(82406) <= 16416131;
srom_1(82407) <= 16230685;
srom_1(82408) <= 16008464;
srom_1(82409) <= 15750511;
srom_1(82410) <= 15458035;
srom_1(82411) <= 15132408;
srom_1(82412) <= 14775158;
srom_1(82413) <= 14387959;
srom_1(82414) <= 13972626;
srom_1(82415) <= 13531109;
srom_1(82416) <= 13065476;
srom_1(82417) <= 12577912;
srom_1(82418) <= 12070703;
srom_1(82419) <= 11546227;
srom_1(82420) <= 11006944;
srom_1(82421) <= 10455383;
srom_1(82422) <= 9894130;
srom_1(82423) <= 9325817;
srom_1(82424) <= 8753109;
srom_1(82425) <= 8178691;
srom_1(82426) <= 7605259;
srom_1(82427) <= 7035499;
srom_1(82428) <= 6472085;
srom_1(82429) <= 5917658;
srom_1(82430) <= 5374818;
srom_1(82431) <= 4846111;
srom_1(82432) <= 4334016;
srom_1(82433) <= 3840934;
srom_1(82434) <= 3369178;
srom_1(82435) <= 2920959;
srom_1(82436) <= 2498380;
srom_1(82437) <= 2103423;
srom_1(82438) <= 1737939;
srom_1(82439) <= 1403642;
srom_1(82440) <= 1102100;
srom_1(82441) <= 834727;
srom_1(82442) <= 602777;
srom_1(82443) <= 407337;
srom_1(82444) <= 249324;
srom_1(82445) <= 129479;
srom_1(82446) <= 48364;
srom_1(82447) <= 6359;
srom_1(82448) <= 3662;
srom_1(82449) <= 40284;
srom_1(82450) <= 116054;
srom_1(82451) <= 230618;
srom_1(82452) <= 383437;
srom_1(82453) <= 573794;
srom_1(82454) <= 800799;
srom_1(82455) <= 1063385;
srom_1(82456) <= 1360321;
srom_1(82457) <= 1690216;
srom_1(82458) <= 2051521;
srom_1(82459) <= 2442544;
srom_1(82460) <= 2861449;
srom_1(82461) <= 3306274;
srom_1(82462) <= 3774931;
srom_1(82463) <= 4265223;
srom_1(82464) <= 4774851;
srom_1(82465) <= 5301425;
srom_1(82466) <= 5842476;
srom_1(82467) <= 6395467;
srom_1(82468) <= 6957805;
srom_1(82469) <= 7526851;
srom_1(82470) <= 8099939;
srom_1(82471) <= 8674381;
srom_1(82472) <= 9247482;
srom_1(82473) <= 9816556;
srom_1(82474) <= 10378934;
srom_1(82475) <= 10931978;
srom_1(82476) <= 11473096;
srom_1(82477) <= 11999750;
srom_1(82478) <= 12509469;
srom_1(82479) <= 12999865;
srom_1(82480) <= 13468636;
srom_1(82481) <= 13913586;
srom_1(82482) <= 14332627;
srom_1(82483) <= 14723795;
srom_1(82484) <= 15085254;
srom_1(82485) <= 15415311;
srom_1(82486) <= 15712417;
srom_1(82487) <= 15975180;
srom_1(82488) <= 16202366;
srom_1(82489) <= 16392911;
srom_1(82490) <= 16545921;
srom_1(82491) <= 16660678;
srom_1(82492) <= 16736645;
srom_1(82493) <= 16773465;
srom_1(82494) <= 16770966;
srom_1(82495) <= 16729159;
srom_1(82496) <= 16648240;
srom_1(82497) <= 16528589;
srom_1(82498) <= 16370766;
srom_1(82499) <= 16175513;
srom_1(82500) <= 15943744;
srom_1(82501) <= 15676547;
srom_1(82502) <= 15375173;
srom_1(82503) <= 15041038;
srom_1(82504) <= 14675707;
srom_1(82505) <= 14280893;
srom_1(82506) <= 13858449;
srom_1(82507) <= 13410354;
srom_1(82508) <= 12938711;
srom_1(82509) <= 12445731;
srom_1(82510) <= 11933726;
srom_1(82511) <= 11405096;
srom_1(82512) <= 10862321;
srom_1(82513) <= 10307946;
srom_1(82514) <= 9744570;
srom_1(82515) <= 9174836;
srom_1(82516) <= 8601415;
srom_1(82517) <= 8026996;
srom_1(82518) <= 7454273;
srom_1(82519) <= 6885931;
srom_1(82520) <= 6324636;
srom_1(82521) <= 5773019;
srom_1(82522) <= 5233668;
srom_1(82523) <= 4709111;
srom_1(82524) <= 4201809;
srom_1(82525) <= 3714140;
srom_1(82526) <= 3248392;
srom_1(82527) <= 2806747;
srom_1(82528) <= 2391278;
srom_1(82529) <= 2003932;
srom_1(82530) <= 1646526;
srom_1(82531) <= 1320737;
srom_1(82532) <= 1028090;
srom_1(82533) <= 769960;
srom_1(82534) <= 547557;
srom_1(82535) <= 361922;
srom_1(82536) <= 213928;
srom_1(82537) <= 104267;
srom_1(82538) <= 33455;
srom_1(82539) <= 1822;
srom_1(82540) <= 9519;
srom_1(82541) <= 56507;
srom_1(82542) <= 142568;
srom_1(82543) <= 267297;
srom_1(82544) <= 430110;
srom_1(82545) <= 630243;
srom_1(82546) <= 866758;
srom_1(82547) <= 1138545;
srom_1(82548) <= 1444330;
srom_1(82549) <= 1782679;
srom_1(82550) <= 2152006;
srom_1(82551) <= 2550578;
srom_1(82552) <= 2976527;
srom_1(82553) <= 3427855;
srom_1(82554) <= 3902445;
srom_1(82555) <= 4398073;
srom_1(82556) <= 4912414;
srom_1(82557) <= 5443056;
srom_1(82558) <= 5987510;
srom_1(82559) <= 6543224;
srom_1(82560) <= 7107592;
srom_1(82561) <= 7677967;
srom_1(82562) <= 8251674;
srom_1(82563) <= 8826023;
srom_1(82564) <= 9398321;
srom_1(82565) <= 9965885;
srom_1(82566) <= 10526051;
srom_1(82567) <= 11076195;
srom_1(82568) <= 11613736;
srom_1(82569) <= 12136152;
srom_1(82570) <= 12640996;
srom_1(82571) <= 13125898;
srom_1(82572) <= 13588586;
srom_1(82573) <= 14026889;
srom_1(82574) <= 14438752;
srom_1(82575) <= 14822244;
srom_1(82576) <= 15175567;
srom_1(82577) <= 15497063;
srom_1(82578) <= 15785225;
srom_1(82579) <= 16038702;
srom_1(82580) <= 16256305;
srom_1(82581) <= 16437014;
srom_1(82582) <= 16579981;
srom_1(82583) <= 16684535;
srom_1(82584) <= 16750188;
srom_1(82585) <= 16776629;
srom_1(82586) <= 16763737;
srom_1(82587) <= 16711571;
srom_1(82588) <= 16620375;
srom_1(82589) <= 16490578;
srom_1(82590) <= 16322788;
srom_1(82591) <= 16117792;
srom_1(82592) <= 15876551;
srom_1(82593) <= 15600197;
srom_1(82594) <= 15290024;
srom_1(82595) <= 14947489;
srom_1(82596) <= 14574197;
srom_1(82597) <= 14171899;
srom_1(82598) <= 13742480;
srom_1(82599) <= 13287956;
srom_1(82600) <= 12810457;
srom_1(82601) <= 12312222;
srom_1(82602) <= 11795588;
srom_1(82603) <= 11262978;
srom_1(82604) <= 10716888;
srom_1(82605) <= 10159881;
srom_1(82606) <= 9594567;
srom_1(82607) <= 9023598;
srom_1(82608) <= 8449652;
srom_1(82609) <= 7875419;
srom_1(82610) <= 7303593;
srom_1(82611) <= 6736855;
srom_1(82612) <= 6177862;
srom_1(82613) <= 5629237;
srom_1(82614) <= 5093551;
srom_1(82615) <= 4573316;
srom_1(82616) <= 4070973;
srom_1(82617) <= 3588877;
srom_1(82618) <= 3129288;
srom_1(82619) <= 2694362;
srom_1(82620) <= 2286139;
srom_1(82621) <= 1906532;
srom_1(82622) <= 1557321;
srom_1(82623) <= 1240145;
srom_1(82624) <= 956490;
srom_1(82625) <= 707688;
srom_1(82626) <= 494903;
srom_1(82627) <= 319135;
srom_1(82628) <= 181208;
srom_1(82629) <= 81767;
srom_1(82630) <= 21281;
srom_1(82631) <= 31;
srom_1(82632) <= 18119;
srom_1(82633) <= 75458;
srom_1(82634) <= 171781;
srom_1(82635) <= 306636;
srom_1(82636) <= 479389;
srom_1(82637) <= 689232;
srom_1(82638) <= 935179;
srom_1(82639) <= 1216079;
srom_1(82640) <= 1530612;
srom_1(82641) <= 1877305;
srom_1(82642) <= 2254532;
srom_1(82643) <= 2660524;
srom_1(82644) <= 3093377;
srom_1(82645) <= 3551060;
srom_1(82646) <= 4031429;
srom_1(82647) <= 4532230;
srom_1(82648) <= 5051115;
srom_1(82649) <= 5585650;
srom_1(82650) <= 6133330;
srom_1(82651) <= 6691585;
srom_1(82652) <= 7257798;
srom_1(82653) <= 7829314;
srom_1(82654) <= 8403453;
srom_1(82655) <= 8977522;
srom_1(82656) <= 9548830;
srom_1(82657) <= 10114696;
srom_1(82658) <= 10672469;
srom_1(82659) <= 11219532;
srom_1(82660) <= 11753319;
srom_1(82661) <= 12271328;
srom_1(82662) <= 12771130;
srom_1(82663) <= 13250381;
srom_1(82664) <= 13706833;
srom_1(82665) <= 14138346;
srom_1(82666) <= 14542897;
srom_1(82667) <= 14918588;
srom_1(82668) <= 15263657;
srom_1(82669) <= 15576488;
srom_1(82670) <= 15855612;
srom_1(82671) <= 16099720;
srom_1(82672) <= 16307668;
srom_1(82673) <= 16478482;
srom_1(82674) <= 16611359;
srom_1(82675) <= 16705676;
srom_1(82676) <= 16760992;
srom_1(82677) <= 16777047;
srom_1(82678) <= 16753766;
srom_1(82679) <= 16691258;
srom_1(82680) <= 16589816;
srom_1(82681) <= 16449915;
srom_1(82682) <= 16272212;
srom_1(82683) <= 16057540;
srom_1(82684) <= 15806906;
srom_1(82685) <= 15521485;
srom_1(82686) <= 15202616;
srom_1(82687) <= 14851793;
srom_1(82688) <= 14470662;
srom_1(82689) <= 14061011;
srom_1(82690) <= 13624759;
srom_1(82691) <= 13163953;
srom_1(82692) <= 12680755;
srom_1(82693) <= 12177428;
srom_1(82694) <= 11656335;
srom_1(82695) <= 11119918;
srom_1(82696) <= 10570693;
srom_1(82697) <= 10011236;
srom_1(82698) <= 9444169;
srom_1(82699) <= 8872153;
srom_1(82700) <= 8297869;
srom_1(82701) <= 7724010;
srom_1(82702) <= 7153269;
srom_1(82703) <= 6588320;
srom_1(82704) <= 6031813;
srom_1(82705) <= 5486358;
srom_1(82706) <= 4954512;
srom_1(82707) <= 4438771;
srom_1(82708) <= 3941551;
srom_1(82709) <= 3465185;
srom_1(82710) <= 3011907;
srom_1(82711) <= 2583842;
srom_1(82712) <= 2182998;
srom_1(82713) <= 1811253;
srom_1(82714) <= 1470353;
srom_1(82715) <= 1161894;
srom_1(82716) <= 887324;
srom_1(82717) <= 647930;
srom_1(82718) <= 444834;
srom_1(82719) <= 278990;
srom_1(82720) <= 151174;
srom_1(82721) <= 61987;
srom_1(82722) <= 11846;
srom_1(82723) <= 987;
srom_1(82724) <= 29459;
srom_1(82725) <= 97131;
srom_1(82726) <= 203685;
srom_1(82727) <= 348620;
srom_1(82728) <= 531258;
srom_1(82729) <= 750741;
srom_1(82730) <= 1006041;
srom_1(82731) <= 1295960;
srom_1(82732) <= 1619140;
srom_1(82733) <= 1974063;
srom_1(82734) <= 2359067;
srom_1(82735) <= 2772345;
srom_1(82736) <= 3211960;
srom_1(82737) <= 3675850;
srom_1(82738) <= 4161839;
srom_1(82739) <= 4667649;
srom_1(82740) <= 5190909;
srom_1(82741) <= 5729163;
srom_1(82742) <= 6279888;
srom_1(82743) <= 6840502;
srom_1(82744) <= 7408375;
srom_1(82745) <= 7980845;
srom_1(82746) <= 8555228;
srom_1(82747) <= 9128828;
srom_1(82748) <= 9698958;
srom_1(82749) <= 10262943;
srom_1(82750) <= 10818139;
srom_1(82751) <= 11361941;
srom_1(82752) <= 11891801;
srom_1(82753) <= 12405233;
srom_1(82754) <= 12899830;
srom_1(82755) <= 13373272;
srom_1(82756) <= 13823339;
srom_1(82757) <= 14247921;
srom_1(82758) <= 14645026;
srom_1(82759) <= 15012793;
srom_1(82760) <= 15349497;
srom_1(82761) <= 15653559;
srom_1(82762) <= 15923553;
srom_1(82763) <= 16158213;
srom_1(82764) <= 16356439;
srom_1(82765) <= 16517301;
srom_1(82766) <= 16640044;
srom_1(82767) <= 16724094;
srom_1(82768) <= 16769056;
srom_1(82769) <= 16774719;
srom_1(82770) <= 16741057;
srom_1(82771) <= 16668227;
srom_1(82772) <= 16556571;
srom_1(82773) <= 16406613;
srom_1(82774) <= 16219055;
srom_1(82775) <= 15994778;
srom_1(82776) <= 15734833;
srom_1(82777) <= 15440439;
srom_1(82778) <= 15112977;
srom_1(82779) <= 14753981;
srom_1(82780) <= 14365136;
srom_1(82781) <= 13948266;
srom_1(82782) <= 13505324;
srom_1(82783) <= 13038388;
srom_1(82784) <= 12549647;
srom_1(82785) <= 12041394;
srom_1(82786) <= 11516012;
srom_1(82787) <= 10975964;
srom_1(82788) <= 10423784;
srom_1(82789) <= 9862060;
srom_1(82790) <= 9293426;
srom_1(82791) <= 8720549;
srom_1(82792) <= 8146116;
srom_1(82793) <= 7572819;
srom_1(82794) <= 7003348;
srom_1(82795) <= 6440374;
srom_1(82796) <= 5886535;
srom_1(82797) <= 5344429;
srom_1(82798) <= 4816598;
srom_1(82799) <= 4305518;
srom_1(82800) <= 3813585;
srom_1(82801) <= 3343105;
srom_1(82802) <= 2896286;
srom_1(82803) <= 2475222;
srom_1(82804) <= 2081888;
srom_1(82805) <= 1718128;
srom_1(82806) <= 1385649;
srom_1(82807) <= 1086009;
srom_1(82808) <= 820613;
srom_1(82809) <= 590706;
srom_1(82810) <= 397366;
srom_1(82811) <= 241500;
srom_1(82812) <= 123838;
srom_1(82813) <= 44933;
srom_1(82814) <= 5154;
srom_1(82815) <= 4688;
srom_1(82816) <= 43537;
srom_1(82817) <= 121519;
srom_1(82818) <= 238268;
srom_1(82819) <= 393237;
srom_1(82820) <= 585699;
srom_1(82821) <= 814751;
srom_1(82822) <= 1079320;
srom_1(82823) <= 1378165;
srom_1(82824) <= 1709883;
srom_1(82825) <= 2072921;
srom_1(82826) <= 2465575;
srom_1(82827) <= 2886005;
srom_1(82828) <= 3332238;
srom_1(82829) <= 3802182;
srom_1(82830) <= 4293633;
srom_1(82831) <= 4804287;
srom_1(82832) <= 5331749;
srom_1(82833) <= 5873546;
srom_1(82834) <= 6427137;
srom_1(82835) <= 6989926;
srom_1(82836) <= 7559273;
srom_1(82837) <= 8132510;
srom_1(82838) <= 8706948;
srom_1(82839) <= 9279892;
srom_1(82840) <= 9848658;
srom_1(82841) <= 10410576;
srom_1(82842) <= 10963013;
srom_1(82843) <= 11503378;
srom_1(82844) <= 12029136;
srom_1(82845) <= 12537823;
srom_1(82846) <= 13027052;
srom_1(82847) <= 13494531;
srom_1(82848) <= 13938066;
srom_1(82849) <= 14355577;
srom_1(82850) <= 14745107;
srom_1(82851) <= 15104830;
srom_1(82852) <= 15433058;
srom_1(82853) <= 15728252;
srom_1(82854) <= 15989028;
srom_1(82855) <= 16214163;
srom_1(82856) <= 16402601;
srom_1(82857) <= 16553459;
srom_1(82858) <= 16666029;
srom_1(82859) <= 16739783;
srom_1(82860) <= 16774376;
srom_1(82861) <= 16769645;
srom_1(82862) <= 16725613;
srom_1(82863) <= 16642485;
srom_1(82864) <= 16520652;
srom_1(82865) <= 16360685;
srom_1(82866) <= 16163335;
srom_1(82867) <= 15929526;
srom_1(82868) <= 15660355;
srom_1(82869) <= 15357084;
srom_1(82870) <= 15021136;
srom_1(82871) <= 14654085;
srom_1(82872) <= 14257654;
srom_1(82873) <= 13833700;
srom_1(82874) <= 13384213;
srom_1(82875) <= 12911300;
srom_1(82876) <= 12417178;
srom_1(82877) <= 11904164;
srom_1(82878) <= 11374665;
srom_1(82879) <= 10831164;
srom_1(82880) <= 10276208;
srom_1(82881) <= 9712401;
srom_1(82882) <= 9142386;
srom_1(82883) <= 8568836;
srom_1(82884) <= 7994441;
srom_1(82885) <= 7421895;
srom_1(82886) <= 6853882;
srom_1(82887) <= 6293065;
srom_1(82888) <= 5742076;
srom_1(82889) <= 5203497;
srom_1(82890) <= 4679854;
srom_1(82891) <= 4173602;
srom_1(82892) <= 3687116;
srom_1(82893) <= 3222677;
srom_1(82894) <= 2782463;
srom_1(82895) <= 2368538;
srom_1(82896) <= 1982843;
srom_1(82897) <= 1627187;
srom_1(82898) <= 1303238;
srom_1(82899) <= 1012514;
srom_1(82900) <= 756380;
srom_1(82901) <= 536035;
srom_1(82902) <= 352514;
srom_1(82903) <= 206677;
srom_1(82904) <= 99208;
srom_1(82905) <= 30610;
srom_1(82906) <= 1206;
srom_1(82907) <= 11134;
srom_1(82908) <= 60346;
srom_1(82909) <= 148613;
srom_1(82910) <= 275519;
srom_1(82911) <= 440471;
srom_1(82912) <= 642694;
srom_1(82913) <= 881241;
srom_1(82914) <= 1154992;
srom_1(82915) <= 1462664;
srom_1(82916) <= 1802814;
srom_1(82917) <= 2173847;
srom_1(82918) <= 2574023;
srom_1(82919) <= 3001466;
srom_1(82920) <= 3454171;
srom_1(82921) <= 3930015;
srom_1(82922) <= 4426768;
srom_1(82923) <= 4942098;
srom_1(82924) <= 5473591;
srom_1(82925) <= 6018752;
srom_1(82926) <= 6575027;
srom_1(82927) <= 7139807;
srom_1(82928) <= 7710443;
srom_1(82929) <= 8284258;
srom_1(82930) <= 8858563;
srom_1(82931) <= 9430664;
srom_1(82932) <= 9997879;
srom_1(82933) <= 10557547;
srom_1(82934) <= 11107045;
srom_1(82935) <= 11643794;
srom_1(82936) <= 12165279;
srom_1(82937) <= 12669054;
srom_1(82938) <= 13152756;
srom_1(82939) <= 13614118;
srom_1(82940) <= 14050975;
srom_1(82941) <= 14461280;
srom_1(82942) <= 14843108;
srom_1(82943) <= 15194668;
srom_1(82944) <= 15514312;
srom_1(82945) <= 15800542;
srom_1(82946) <= 16052014;
srom_1(82947) <= 16267550;
srom_1(82948) <= 16446139;
srom_1(82949) <= 16586944;
srom_1(82950) <= 16689303;
srom_1(82951) <= 16752738;
srom_1(82952) <= 16776951;
srom_1(82953) <= 16761827;
srom_1(82954) <= 16707439;
srom_1(82955) <= 16614041;
srom_1(82956) <= 16482071;
srom_1(82957) <= 16312148;
srom_1(82958) <= 16105069;
srom_1(82959) <= 15861804;
srom_1(82960) <= 15583496;
srom_1(82961) <= 15271448;
srom_1(82962) <= 14927124;
srom_1(82963) <= 14552138;
srom_1(82964) <= 14148250;
srom_1(82965) <= 13717352;
srom_1(82966) <= 13261467;
srom_1(82967) <= 12782731;
srom_1(82968) <= 12283389;
srom_1(82969) <= 11765783;
srom_1(82970) <= 11232341;
srom_1(82971) <= 10685563;
srom_1(82972) <= 10128014;
srom_1(82973) <= 9562309;
srom_1(82974) <= 8991099;
srom_1(82975) <= 8417065;
srom_1(82976) <= 7842897;
srom_1(82977) <= 7271287;
srom_1(82978) <= 6704918;
srom_1(82979) <= 6146443;
srom_1(82980) <= 5598483;
srom_1(82981) <= 5063607;
srom_1(82982) <= 4544323;
srom_1(82983) <= 4043066;
srom_1(82984) <= 3562187;
srom_1(82985) <= 3103941;
srom_1(82986) <= 2670476;
srom_1(82987) <= 2263825;
srom_1(82988) <= 1885896;
srom_1(82989) <= 1538460;
srom_1(82990) <= 1223147;
srom_1(82991) <= 941435;
srom_1(82992) <= 694645;
srom_1(82993) <= 483935;
srom_1(82994) <= 310293;
srom_1(82995) <= 174533;
srom_1(82996) <= 77291;
srom_1(82997) <= 19024;
srom_1(82998) <= 5;
srom_1(82999) <= 20323;
srom_1(83000) <= 79882;
srom_1(83001) <= 178404;
srom_1(83002) <= 315427;
srom_1(83003) <= 490307;
srom_1(83004) <= 702226;
srom_1(83005) <= 950188;
srom_1(83006) <= 1233032;
srom_1(83007) <= 1549430;
srom_1(83008) <= 1897900;
srom_1(83009) <= 2276807;
srom_1(83010) <= 2684375;
srom_1(83011) <= 3118691;
srom_1(83012) <= 3577720;
srom_1(83013) <= 4059309;
srom_1(83014) <= 4561199;
srom_1(83015) <= 5081038;
srom_1(83016) <= 5616386;
srom_1(83017) <= 6164735;
srom_1(83018) <= 6723512;
srom_1(83019) <= 7290097;
srom_1(83020) <= 7861834;
srom_1(83021) <= 8436041;
srom_1(83022) <= 9010025;
srom_1(83023) <= 9581095;
srom_1(83024) <= 10146574;
srom_1(83025) <= 10703808;
srom_1(83026) <= 11250186;
srom_1(83027) <= 11783145;
srom_1(83028) <= 12300186;
srom_1(83029) <= 12798884;
srom_1(83030) <= 13276901;
srom_1(83031) <= 13731994;
srom_1(83032) <= 14162031;
srom_1(83033) <= 14564995;
srom_1(83034) <= 14938995;
srom_1(83035) <= 15282278;
srom_1(83036) <= 15593234;
srom_1(83037) <= 15870405;
srom_1(83038) <= 16112492;
srom_1(83039) <= 16318358;
srom_1(83040) <= 16487040;
srom_1(83041) <= 16617745;
srom_1(83042) <= 16709860;
srom_1(83043) <= 16762955;
srom_1(83044) <= 16776779;
srom_1(83045) <= 16751268;
srom_1(83046) <= 16686542;
srom_1(83047) <= 16582904;
srom_1(83048) <= 16440840;
srom_1(83049) <= 16261017;
srom_1(83050) <= 16044277;
srom_1(83051) <= 15791636;
srom_1(83052) <= 15504281;
srom_1(83053) <= 15183558;
srom_1(83054) <= 14830971;
srom_1(83055) <= 14448173;
srom_1(83056) <= 14036960;
srom_1(83057) <= 13599260;
srom_1(83058) <= 13137125;
srom_1(83059) <= 12652723;
srom_1(83060) <= 12148325;
srom_1(83061) <= 11626297;
srom_1(83062) <= 11089086;
srom_1(83063) <= 10539211;
srom_1(83064) <= 9979251;
srom_1(83065) <= 9411833;
srom_1(83066) <= 8839616;
srom_1(83067) <= 8265284;
srom_1(83068) <= 7691530;
srom_1(83069) <= 7121045;
srom_1(83070) <= 6556505;
srom_1(83071) <= 6000555;
srom_1(83072) <= 5455804;
srom_1(83073) <= 4924806;
srom_1(83074) <= 4410051;
srom_1(83075) <= 3913953;
srom_1(83076) <= 3438838;
srom_1(83077) <= 2986934;
srom_1(83078) <= 2560360;
srom_1(83079) <= 2161117;
srom_1(83080) <= 1791077;
srom_1(83081) <= 1451975;
srom_1(83082) <= 1145401;
srom_1(83083) <= 872793;
srom_1(83084) <= 635430;
srom_1(83085) <= 434423;
srom_1(83086) <= 270717;
srom_1(83087) <= 145078;
srom_1(83088) <= 58096;
srom_1(83089) <= 10178;
srom_1(83090) <= 1550;
srom_1(83091) <= 32251;
srom_1(83092) <= 102139;
srom_1(83093) <= 210884;
srom_1(83094) <= 357978;
srom_1(83095) <= 542730;
srom_1(83096) <= 764274;
srom_1(83097) <= 1021571;
srom_1(83098) <= 1313415;
srom_1(83099) <= 1638436;
srom_1(83100) <= 1995112;
srom_1(83101) <= 2381769;
srom_1(83102) <= 2796594;
srom_1(83103) <= 3237641;
srom_1(83104) <= 3702844;
srom_1(83105) <= 4190020;
srom_1(83106) <= 4696884;
srom_1(83107) <= 5221060;
srom_1(83108) <= 5760090;
srom_1(83109) <= 6311445;
srom_1(83110) <= 6872542;
srom_1(83111) <= 7440747;
srom_1(83112) <= 8013398;
srom_1(83113) <= 8587808;
srom_1(83114) <= 9161283;
srom_1(83115) <= 9731136;
srom_1(83116) <= 10294693;
srom_1(83117) <= 10849311;
srom_1(83118) <= 11392391;
srom_1(83119) <= 11921385;
srom_1(83120) <= 12433812;
srom_1(83121) <= 12927270;
srom_1(83122) <= 13399445;
srom_1(83123) <= 13848122;
srom_1(83124) <= 14271197;
srom_1(83125) <= 14666687;
srom_1(83126) <= 15032737;
srom_1(83127) <= 15367630;
srom_1(83128) <= 15669797;
srom_1(83129) <= 15937819;
srom_1(83130) <= 16170441;
srom_1(83131) <= 16366570;
srom_1(83132) <= 16525289;
srom_1(83133) <= 16645851;
srom_1(83134) <= 16727693;
srom_1(83135) <= 16770430;
srom_1(83136) <= 16773861;
srom_1(83137) <= 16737971;
srom_1(83138) <= 16662928;
srom_1(83139) <= 16549084;
srom_1(83140) <= 16396973;
srom_1(83141) <= 16207308;
srom_1(83142) <= 15980978;
srom_1(83143) <= 15719045;
srom_1(83144) <= 15422737;
srom_1(83145) <= 15093443;
srom_1(83146) <= 14732708;
srom_1(83147) <= 14342224;
srom_1(83148) <= 13923821;
srom_1(83149) <= 13479461;
srom_1(83150) <= 13011229;
srom_1(83151) <= 12521320;
srom_1(83152) <= 12012031;
srom_1(83153) <= 11485750;
srom_1(83154) <= 10944946;
srom_1(83155) <= 10392154;
srom_1(83156) <= 9829967;
srom_1(83157) <= 9261021;
srom_1(83158) <= 8687984;
srom_1(83159) <= 8113543;
srom_1(83160) <= 7540392;
srom_1(83161) <= 6971219;
srom_1(83162) <= 6408692;
srom_1(83163) <= 5855449;
srom_1(83164) <= 5314086;
srom_1(83165) <= 4787139;
srom_1(83166) <= 4277082;
srom_1(83167) <= 3786305;
srom_1(83168) <= 3317109;
srom_1(83169) <= 2871696;
srom_1(83170) <= 2452153;
srom_1(83171) <= 2060448;
srom_1(83172) <= 1698418;
srom_1(83173) <= 1367761;
srom_1(83174) <= 1070027;
srom_1(83175) <= 806613;
srom_1(83176) <= 578752;
srom_1(83177) <= 387515;
srom_1(83178) <= 233798;
srom_1(83179) <= 118322;
srom_1(83180) <= 41627;
srom_1(83181) <= 4075;
srom_1(83182) <= 5840;
srom_1(83183) <= 46916;
srom_1(83184) <= 127108;
srom_1(83185) <= 246041;
srom_1(83186) <= 403158;
srom_1(83187) <= 597721;
srom_1(83188) <= 828818;
srom_1(83189) <= 1095366;
srom_1(83190) <= 1396114;
srom_1(83191) <= 1729652;
srom_1(83192) <= 2094416;
srom_1(83193) <= 2488697;
srom_1(83194) <= 2910643;
srom_1(83195) <= 3358278;
srom_1(83196) <= 3829502;
srom_1(83197) <= 4322105;
srom_1(83198) <= 4833777;
srom_1(83199) <= 5362119;
srom_1(83200) <= 5904654;
srom_1(83201) <= 6458836;
srom_1(83202) <= 7022068;
srom_1(83203) <= 7591708;
srom_1(83204) <= 8165084;
srom_1(83205) <= 8739509;
srom_1(83206) <= 9312289;
srom_1(83207) <= 9880737;
srom_1(83208) <= 10442188;
srom_1(83209) <= 10994009;
srom_1(83210) <= 11533612;
srom_1(83211) <= 12058468;
srom_1(83212) <= 12566114;
srom_1(83213) <= 13054170;
srom_1(83214) <= 13520348;
srom_1(83215) <= 13962461;
srom_1(83216) <= 14378437;
srom_1(83217) <= 14766324;
srom_1(83218) <= 15124304;
srom_1(83219) <= 15450698;
srom_1(83220) <= 15743976;
srom_1(83221) <= 16002761;
srom_1(83222) <= 16225842;
srom_1(83223) <= 16412170;
srom_1(83224) <= 16560874;
srom_1(83225) <= 16671255;
srom_1(83226) <= 16742795;
srom_1(83227) <= 16775160;
srom_1(83228) <= 16768198;
srom_1(83229) <= 16721941;
srom_1(83230) <= 16636606;
srom_1(83231) <= 16512593;
srom_1(83232) <= 16350484;
srom_1(83233) <= 16151039;
srom_1(83234) <= 15915194;
srom_1(83235) <= 15644053;
srom_1(83236) <= 15338890;
srom_1(83237) <= 15001134;
srom_1(83238) <= 14632369;
srom_1(83239) <= 14234326;
srom_1(83240) <= 13808870;
srom_1(83241) <= 13357996;
srom_1(83242) <= 12883820;
srom_1(83243) <= 12388563;
srom_1(83244) <= 11874550;
srom_1(83245) <= 11344190;
srom_1(83246) <= 10799970;
srom_1(83247) <= 10244442;
srom_1(83248) <= 9680212;
srom_1(83249) <= 9109924;
srom_1(83250) <= 8536255;
srom_1(83251) <= 7961893;
srom_1(83252) <= 7389532;
srom_1(83253) <= 6821856;
srom_1(83254) <= 6261527;
srom_1(83255) <= 5711172;
srom_1(83256) <= 5173373;
srom_1(83257) <= 4650652;
srom_1(83258) <= 4145459;
srom_1(83259) <= 3660163;
srom_1(83260) <= 3197041;
srom_1(83261) <= 2758264;
srom_1(83262) <= 2345889;
srom_1(83263) <= 1961851;
srom_1(83264) <= 1607950;
srom_1(83265) <= 1285846;
srom_1(83266) <= 997049;
srom_1(83267) <= 742914;
srom_1(83268) <= 524632;
srom_1(83269) <= 343227;
srom_1(83270) <= 199549;
srom_1(83271) <= 94273;
srom_1(83272) <= 27892;
srom_1(83273) <= 717;
srom_1(83274) <= 12876;
srom_1(83275) <= 64311;
srom_1(83276) <= 154782;
srom_1(83277) <= 283864;
srom_1(83278) <= 450952;
srom_1(83279) <= 655262;
srom_1(83280) <= 895837;
srom_1(83281) <= 1171548;
srom_1(83282) <= 1481102;
srom_1(83283) <= 1823048;
srom_1(83284) <= 2195782;
srom_1(83285) <= 2597556;
srom_1(83286) <= 3026487;
srom_1(83287) <= 3480562;
srom_1(83288) <= 3957653;
srom_1(83289) <= 4455522;
srom_1(83290) <= 4971834;
srom_1(83291) <= 5504169;
srom_1(83292) <= 6050031;
srom_1(83293) <= 6606858;
srom_1(83294) <= 7172041;
srom_1(83295) <= 7742929;
srom_1(83296) <= 8316844;
srom_1(83297) <= 8891096;
srom_1(83298) <= 9462992;
srom_1(83299) <= 10029849;
srom_1(83300) <= 10589011;
srom_1(83301) <= 11137853;
srom_1(83302) <= 11673804;
srom_1(83303) <= 12194349;
srom_1(83304) <= 12697048;
srom_1(83305) <= 13179543;
srom_1(83306) <= 13639571;
srom_1(83307) <= 14074976;
srom_1(83308) <= 14483716;
srom_1(83309) <= 14863873;
srom_1(83310) <= 15213666;
srom_1(83311) <= 15531454;
srom_1(83312) <= 15815747;
srom_1(83313) <= 16065211;
srom_1(83314) <= 16278677;
srom_1(83315) <= 16455143;
srom_1(83316) <= 16593783;
srom_1(83317) <= 16693946;
srom_1(83318) <= 16755163;
srom_1(83319) <= 16777145;
srom_1(83320) <= 16759791;
srom_1(83321) <= 16703182;
srom_1(83322) <= 16607583;
srom_1(83323) <= 16473442;
srom_1(83324) <= 16301388;
srom_1(83325) <= 16092229;
srom_1(83326) <= 15846945;
srom_1(83327) <= 15566686;
srom_1(83328) <= 15252767;
srom_1(83329) <= 14906659;
srom_1(83330) <= 14529986;
srom_1(83331) <= 14124514;
srom_1(83332) <= 13692144;
srom_1(83333) <= 13234904;
srom_1(83334) <= 12754938;
srom_1(83335) <= 12254497;
srom_1(83336) <= 11735928;
srom_1(83337) <= 11201661;
srom_1(83338) <= 10654204;
srom_1(83339) <= 10096122;
srom_1(83340) <= 9530033;
srom_1(83341) <= 8958591;
srom_1(83342) <= 8384477;
srom_1(83343) <= 7810382;
srom_1(83344) <= 7238998;
srom_1(83345) <= 6673006;
srom_1(83346) <= 6115058;
srom_1(83347) <= 5567772;
srom_1(83348) <= 5033714;
srom_1(83349) <= 4515388;
srom_1(83350) <= 4015225;
srom_1(83351) <= 3535570;
srom_1(83352) <= 3078672;
srom_1(83353) <= 2646675;
srom_1(83354) <= 2241604;
srom_1(83355) <= 1865358;
srom_1(83356) <= 1519702;
srom_1(83357) <= 1206256;
srom_1(83358) <= 926491;
srom_1(83359) <= 681719;
srom_1(83360) <= 473086;
srom_1(83361) <= 301573;
srom_1(83362) <= 167982;
srom_1(83363) <= 72940;
srom_1(83364) <= 16894;
srom_1(83365) <= 105;
srom_1(83366) <= 22653;
srom_1(83367) <= 84432;
srom_1(83368) <= 185151;
srom_1(83369) <= 324340;
srom_1(83370) <= 501345;
srom_1(83371) <= 715336;
srom_1(83372) <= 965309;
srom_1(83373) <= 1250093;
srom_1(83374) <= 1568352;
srom_1(83375) <= 1918593;
srom_1(83376) <= 2299175;
srom_1(83377) <= 2708312;
srom_1(83378) <= 3144085;
srom_1(83379) <= 3604452;
srom_1(83380) <= 4087254;
srom_1(83381) <= 4590226;
srom_1(83382) <= 5111010;
srom_1(83383) <= 5647164;
srom_1(83384) <= 6196173;
srom_1(83385) <= 6755464;
srom_1(83386) <= 7322413;
srom_1(83387) <= 7894361;
srom_1(83388) <= 8468628;
srom_1(83389) <= 9042519;
srom_1(83390) <= 9613343;
srom_1(83391) <= 10178425;
srom_1(83392) <= 10735113;
srom_1(83393) <= 11280798;
srom_1(83394) <= 11812920;
srom_1(83395) <= 12328984;
srom_1(83396) <= 12826571;
srom_1(83397) <= 13303347;
srom_1(83398) <= 13757075;
srom_1(83399) <= 14185629;
srom_1(83400) <= 14586999;
srom_1(83401) <= 14959303;
srom_1(83402) <= 15300794;
srom_1(83403) <= 15609871;
srom_1(83404) <= 15885086;
srom_1(83405) <= 16125147;
srom_1(83406) <= 16328929;
srom_1(83407) <= 16495476;
srom_1(83408) <= 16624006;
srom_1(83409) <= 16713919;
srom_1(83410) <= 16764791;
srom_1(83411) <= 16776384;
srom_1(83412) <= 16748644;
srom_1(83413) <= 16681701;
srom_1(83414) <= 16575869;
srom_1(83415) <= 16431644;
srom_1(83416) <= 16249702;
srom_1(83417) <= 16030897;
srom_1(83418) <= 15776255;
srom_1(83419) <= 15486969;
srom_1(83420) <= 15164397;
srom_1(83421) <= 14810051;
srom_1(83422) <= 14425592;
srom_1(83423) <= 14012824;
srom_1(83424) <= 13573682;
srom_1(83425) <= 13110225;
srom_1(83426) <= 12624628;
srom_1(83427) <= 12119166;
srom_1(83428) <= 11596210;
srom_1(83429) <= 11058212;
srom_1(83430) <= 10507696;
srom_1(83431) <= 9947243;
srom_1(83432) <= 9379480;
srom_1(83433) <= 8807072;
srom_1(83434) <= 8232700;
srom_1(83435) <= 7659060;
srom_1(83436) <= 7088841;
srom_1(83437) <= 6524718;
srom_1(83438) <= 5969334;
srom_1(83439) <= 5425295;
srom_1(83440) <= 4895153;
srom_1(83441) <= 4381392;
srom_1(83442) <= 3886422;
srom_1(83443) <= 3412565;
srom_1(83444) <= 2962042;
srom_1(83445) <= 2536966;
srom_1(83446) <= 2139331;
srom_1(83447) <= 1771000;
srom_1(83448) <= 1433702;
srom_1(83449) <= 1129018;
srom_1(83450) <= 858376;
srom_1(83451) <= 623047;
srom_1(83452) <= 424132;
srom_1(83453) <= 262566;
srom_1(83454) <= 139105;
srom_1(83455) <= 54330;
srom_1(83456) <= 8636;
srom_1(83457) <= 2239;
srom_1(83458) <= 35169;
srom_1(83459) <= 107271;
srom_1(83460) <= 218207;
srom_1(83461) <= 367457;
srom_1(83462) <= 554320;
srom_1(83463) <= 777921;
srom_1(83464) <= 1037212;
srom_1(83465) <= 1330975;
srom_1(83466) <= 1657835;
srom_1(83467) <= 2016257;
srom_1(83468) <= 2404561;
srom_1(83469) <= 2820927;
srom_1(83470) <= 3263401;
srom_1(83471) <= 3729909;
srom_1(83472) <= 4218264;
srom_1(83473) <= 4726174;
srom_1(83474) <= 5251259;
srom_1(83475) <= 5791056;
srom_1(83476) <= 6343034;
srom_1(83477) <= 6904604;
srom_1(83478) <= 7473133;
srom_1(83479) <= 8045956;
srom_1(83480) <= 8620385;
srom_1(83481) <= 9193727;
srom_1(83482) <= 9763294;
srom_1(83483) <= 10326414;
srom_1(83484) <= 10880447;
srom_1(83485) <= 11422795;
srom_1(83486) <= 11950915;
srom_1(83487) <= 12462330;
srom_1(83488) <= 12954642;
srom_1(83489) <= 13425542;
srom_1(83490) <= 13872822;
srom_1(83491) <= 14294385;
srom_1(83492) <= 14688253;
srom_1(83493) <= 15052581;
srom_1(83494) <= 15385658;
srom_1(83495) <= 15685925;
srom_1(83496) <= 15951971;
srom_1(83497) <= 16182550;
srom_1(83498) <= 16376581;
srom_1(83499) <= 16533154;
srom_1(83500) <= 16651533;
srom_1(83501) <= 16731166;
srom_1(83502) <= 16771677;
srom_1(83503) <= 16772877;
srom_1(83504) <= 16734760;
srom_1(83505) <= 16657505;
srom_1(83506) <= 16541475;
srom_1(83507) <= 16387213;
srom_1(83508) <= 16195442;
srom_1(83509) <= 15967063;
srom_1(83510) <= 15703146;
srom_1(83511) <= 15404928;
srom_1(83512) <= 15073809;
srom_1(83513) <= 14711340;
srom_1(83514) <= 14319222;
srom_1(83515) <= 13899293;
srom_1(83516) <= 13453522;
srom_1(83517) <= 12984001;
srom_1(83518) <= 12492930;
srom_1(83519) <= 11982613;
srom_1(83520) <= 11455441;
srom_1(83521) <= 10913889;
srom_1(83522) <= 10360495;
srom_1(83523) <= 9797853;
srom_1(83524) <= 9228604;
srom_1(83525) <= 8655415;
srom_1(83526) <= 8080975;
srom_1(83527) <= 7507978;
srom_1(83528) <= 6939110;
srom_1(83529) <= 6377039;
srom_1(83530) <= 5824402;
srom_1(83531) <= 5283789;
srom_1(83532) <= 4757735;
srom_1(83533) <= 4248708;
srom_1(83534) <= 3759094;
srom_1(83535) <= 3291190;
srom_1(83536) <= 2847189;
srom_1(83537) <= 2429173;
srom_1(83538) <= 2039104;
srom_1(83539) <= 1678810;
srom_1(83540) <= 1349980;
srom_1(83541) <= 1054156;
srom_1(83542) <= 792727;
srom_1(83543) <= 566917;
srom_1(83544) <= 377785;
srom_1(83545) <= 226220;
srom_1(83546) <= 112930;
srom_1(83547) <= 38448;
srom_1(83548) <= 3122;
srom_1(83549) <= 7120;
srom_1(83550) <= 50420;
srom_1(83551) <= 132822;
srom_1(83552) <= 253937;
srom_1(83553) <= 413199;
srom_1(83554) <= 609860;
srom_1(83555) <= 842999;
srom_1(83556) <= 1111521;
srom_1(83557) <= 1414168;
srom_1(83558) <= 1749521;
srom_1(83559) <= 2116007;
srom_1(83560) <= 2511907;
srom_1(83561) <= 2935365;
srom_1(83562) <= 3384395;
srom_1(83563) <= 3856891;
srom_1(83564) <= 4350638;
srom_1(83565) <= 4863321;
srom_1(83566) <= 5392535;
srom_1(83567) <= 5935799;
srom_1(83568) <= 6490564;
srom_1(83569) <= 7054230;
srom_1(83570) <= 7624154;
srom_1(83571) <= 8197662;
srom_1(83572) <= 8772066;
srom_1(83573) <= 9344672;
srom_1(83574) <= 9912794;
srom_1(83575) <= 10473769;
srom_1(83576) <= 11024965;
srom_1(83577) <= 11563799;
srom_1(83578) <= 12087744;
srom_1(83579) <= 12594342;
srom_1(83580) <= 13081217;
srom_1(83581) <= 13546088;
srom_1(83582) <= 13986773;
srom_1(83583) <= 14401207;
srom_1(83584) <= 14787445;
srom_1(83585) <= 15143677;
srom_1(83586) <= 15468232;
srom_1(83587) <= 15759589;
srom_1(83588) <= 16016380;
srom_1(83589) <= 16237402;
srom_1(83590) <= 16421618;
srom_1(83591) <= 16568165;
srom_1(83592) <= 16676355;
srom_1(83593) <= 16745681;
srom_1(83594) <= 16775818;
srom_1(83595) <= 16766624;
srom_1(83596) <= 16718143;
srom_1(83597) <= 16630602;
srom_1(83598) <= 16504411;
srom_1(83599) <= 16340163;
srom_1(83600) <= 16138626;
srom_1(83601) <= 15900748;
srom_1(83602) <= 15627642;
srom_1(83603) <= 15320590;
srom_1(83604) <= 14981032;
srom_1(83605) <= 14610559;
srom_1(83606) <= 14210910;
srom_1(83607) <= 13783958;
srom_1(83608) <= 13331705;
srom_1(83609) <= 12856272;
srom_1(83610) <= 12359889;
srom_1(83611) <= 11844883;
srom_1(83612) <= 11313669;
srom_1(83613) <= 10768739;
srom_1(83614) <= 10212648;
srom_1(83615) <= 9648003;
srom_1(83616) <= 9077452;
srom_1(83617) <= 8503671;
srom_1(83618) <= 7929350;
srom_1(83619) <= 7357183;
srom_1(83620) <= 6789853;
srom_1(83621) <= 6230020;
srom_1(83622) <= 5680309;
srom_1(83623) <= 5143299;
srom_1(83624) <= 4621506;
srom_1(83625) <= 4117379;
srom_1(83626) <= 3633281;
srom_1(83627) <= 3171483;
srom_1(83628) <= 2734149;
srom_1(83629) <= 2323332;
srom_1(83630) <= 1940956;
srom_1(83631) <= 1588815;
srom_1(83632) <= 1268561;
srom_1(83633) <= 981696;
srom_1(83634) <= 729564;
srom_1(83635) <= 513348;
srom_1(83636) <= 334061;
srom_1(83637) <= 192546;
srom_1(83638) <= 89464;
srom_1(83639) <= 25300;
srom_1(83640) <= 354;
srom_1(83641) <= 14744;
srom_1(83642) <= 68401;
srom_1(83643) <= 161075;
srom_1(83644) <= 292331;
srom_1(83645) <= 461553;
srom_1(83646) <= 667947;
srom_1(83647) <= 910546;
srom_1(83648) <= 1188213;
srom_1(83649) <= 1499645;
srom_1(83650) <= 1843381;
srom_1(83651) <= 2217810;
srom_1(83652) <= 2621176;
srom_1(83653) <= 3051588;
srom_1(83654) <= 3507027;
srom_1(83655) <= 3985357;
srom_1(83656) <= 4484335;
srom_1(83657) <= 5001622;
srom_1(83658) <= 5534792;
srom_1(83659) <= 6081344;
srom_1(83660) <= 6638716;
srom_1(83661) <= 7204293;
srom_1(83662) <= 7775425;
srom_1(83663) <= 8349431;
srom_1(83664) <= 8923622;
srom_1(83665) <= 9495303;
srom_1(83666) <= 10061795;
srom_1(83667) <= 10620441;
srom_1(83668) <= 11168620;
srom_1(83669) <= 11703764;
srom_1(83670) <= 12223361;
srom_1(83671) <= 12724976;
srom_1(83672) <= 13206257;
srom_1(83673) <= 13664945;
srom_1(83674) <= 14098891;
srom_1(83675) <= 14506060;
srom_1(83676) <= 14884542;
srom_1(83677) <= 15232562;
srom_1(83678) <= 15548488;
srom_1(83679) <= 15830839;
srom_1(83680) <= 16078291;
srom_1(83681) <= 16289684;
srom_1(83682) <= 16464026;
srom_1(83683) <= 16600499;
srom_1(83684) <= 16698464;
srom_1(83685) <= 16757461;
srom_1(83686) <= 16777213;
srom_1(83687) <= 16757629;
srom_1(83688) <= 16698799;
srom_1(83689) <= 16601000;
srom_1(83690) <= 16464691;
srom_1(83691) <= 16290509;
srom_1(83692) <= 16079273;
srom_1(83693) <= 15831973;
srom_1(83694) <= 15549768;
srom_1(83695) <= 15233983;
srom_1(83696) <= 14886097;
srom_1(83697) <= 14507741;
srom_1(83698) <= 14100692;
srom_1(83699) <= 13666856;
srom_1(83700) <= 13208268;
srom_1(83701) <= 12727080;
srom_1(83702) <= 12225547;
srom_1(83703) <= 11706022;
srom_1(83704) <= 11170939;
srom_1(83705) <= 10622810;
srom_1(83706) <= 10064203;
srom_1(83707) <= 9497740;
srom_1(83708) <= 8926075;
srom_1(83709) <= 8351889;
srom_1(83710) <= 7777876;
srom_1(83711) <= 7206727;
srom_1(83712) <= 6641120;
srom_1(83713) <= 6083707;
srom_1(83714) <= 5537103;
srom_1(83715) <= 5003871;
srom_1(83716) <= 4486511;
srom_1(83717) <= 3987449;
srom_1(83718) <= 3509026;
srom_1(83719) <= 3053484;
srom_1(83720) <= 2622961;
srom_1(83721) <= 2219475;
srom_1(83722) <= 1844919;
srom_1(83723) <= 1501047;
srom_1(83724) <= 1189474;
srom_1(83725) <= 911660;
srom_1(83726) <= 668909;
srom_1(83727) <= 462357;
srom_1(83728) <= 292974;
srom_1(83729) <= 161555;
srom_1(83730) <= 68715;
srom_1(83731) <= 14890;
srom_1(83732) <= 332;
srom_1(83733) <= 25109;
srom_1(83734) <= 89106;
srom_1(83735) <= 192022;
srom_1(83736) <= 333375;
srom_1(83737) <= 512501;
srom_1(83738) <= 728562;
srom_1(83739) <= 980542;
srom_1(83740) <= 1267262;
srom_1(83741) <= 1587376;
srom_1(83742) <= 1939384;
srom_1(83743) <= 2321634;
srom_1(83744) <= 2732334;
srom_1(83745) <= 3169559;
srom_1(83746) <= 3631257;
srom_1(83747) <= 4115264;
srom_1(83748) <= 4619310;
srom_1(83749) <= 5141032;
srom_1(83750) <= 5677983;
srom_1(83751) <= 6227645;
srom_1(83752) <= 6787440;
srom_1(83753) <= 7354744;
srom_1(83754) <= 7926896;
srom_1(83755) <= 8501213;
srom_1(83756) <= 9075002;
srom_1(83757) <= 9645573;
srom_1(83758) <= 10210248;
srom_1(83759) <= 10766382;
srom_1(83760) <= 11311365;
srom_1(83761) <= 11842643;
srom_1(83762) <= 12357724;
srom_1(83763) <= 12854191;
srom_1(83764) <= 13329719;
srom_1(83765) <= 13782075;
srom_1(83766) <= 14209140;
srom_1(83767) <= 14608910;
srom_1(83768) <= 14979512;
srom_1(83769) <= 15319206;
srom_1(83770) <= 15626400;
srom_1(83771) <= 15899654;
srom_1(83772) <= 16137685;
srom_1(83773) <= 16339379;
srom_1(83774) <= 16503789;
srom_1(83775) <= 16630144;
srom_1(83776) <= 16717852;
srom_1(83777) <= 16766500;
srom_1(83778) <= 16775862;
srom_1(83779) <= 16745894;
srom_1(83780) <= 16676735;
srom_1(83781) <= 16568710;
srom_1(83782) <= 16422326;
srom_1(83783) <= 16238269;
srom_1(83784) <= 16017402;
srom_1(83785) <= 15760762;
srom_1(83786) <= 15469550;
srom_1(83787) <= 15145134;
srom_1(83788) <= 14789034;
srom_1(83789) <= 14402920;
srom_1(83790) <= 13988603;
srom_1(83791) <= 13548026;
srom_1(83792) <= 13083254;
srom_1(83793) <= 12596468;
srom_1(83794) <= 12089950;
srom_1(83795) <= 11566074;
srom_1(83796) <= 11027299;
srom_1(83797) <= 10476149;
srom_1(83798) <= 9915211;
srom_1(83799) <= 9347113;
srom_1(83800) <= 8774521;
srom_1(83801) <= 8200120;
srom_1(83802) <= 7626602;
srom_1(83803) <= 7056657;
srom_1(83804) <= 6492958;
srom_1(83805) <= 5938149;
srom_1(83806) <= 5394831;
srom_1(83807) <= 4865552;
srom_1(83808) <= 4352793;
srom_1(83809) <= 3858960;
srom_1(83810) <= 3386368;
srom_1(83811) <= 2937233;
srom_1(83812) <= 2513661;
srom_1(83813) <= 2117639;
srom_1(83814) <= 1751024;
srom_1(83815) <= 1415534;
srom_1(83816) <= 1112744;
srom_1(83817) <= 844073;
srom_1(83818) <= 610781;
srom_1(83819) <= 413961;
srom_1(83820) <= 254538;
srom_1(83821) <= 133258;
srom_1(83822) <= 50690;
srom_1(83823) <= 7221;
srom_1(83824) <= 3056;
srom_1(83825) <= 38213;
srom_1(83826) <= 112528;
srom_1(83827) <= 225653;
srom_1(83828) <= 377056;
srom_1(83829) <= 566029;
srom_1(83830) <= 791684;
srom_1(83831) <= 1052964;
srom_1(83832) <= 1348643;
srom_1(83833) <= 1677335;
srom_1(83834) <= 2037498;
srom_1(83835) <= 2427444;
srom_1(83836) <= 2845344;
srom_1(83837) <= 3289238;
srom_1(83838) <= 3757045;
srom_1(83839) <= 4246570;
srom_1(83840) <= 4755520;
srom_1(83841) <= 5281506;
srom_1(83842) <= 5822062;
srom_1(83843) <= 6374653;
srom_1(83844) <= 6936689;
srom_1(83845) <= 7505533;
srom_1(83846) <= 8078519;
srom_1(83847) <= 8652958;
srom_1(83848) <= 9226158;
srom_1(83849) <= 9795430;
srom_1(83850) <= 10358106;
srom_1(83851) <= 10911545;
srom_1(83852) <= 11453154;
srom_1(83853) <= 11980391;
srom_1(83854) <= 12490786;
srom_1(83855) <= 12981944;
srom_1(83856) <= 13451563;
srom_1(83857) <= 13897439;
srom_1(83858) <= 14317483;
srom_1(83859) <= 14709724;
srom_1(83860) <= 15072324;
srom_1(83861) <= 15403581;
srom_1(83862) <= 15701942;
srom_1(83863) <= 15966009;
srom_1(83864) <= 16194543;
srom_1(83865) <= 16386471;
srom_1(83866) <= 16540896;
srom_1(83867) <= 16657091;
srom_1(83868) <= 16734513;
srom_1(83869) <= 16772797;
srom_1(83870) <= 16771766;
srom_1(83871) <= 16731422;
srom_1(83872) <= 16651957;
srom_1(83873) <= 16533742;
srom_1(83874) <= 16377331;
srom_1(83875) <= 16183459;
srom_1(83876) <= 15953034;
srom_1(83877) <= 15687137;
srom_1(83878) <= 15387014;
srom_1(83879) <= 15054073;
srom_1(83880) <= 14689876;
srom_1(83881) <= 14296130;
srom_1(83882) <= 13874682;
srom_1(83883) <= 13427507;
srom_1(83884) <= 12956703;
srom_1(83885) <= 12464478;
srom_1(83886) <= 11953140;
srom_1(83887) <= 11425087;
srom_1(83888) <= 10882794;
srom_1(83889) <= 10328805;
srom_1(83890) <= 9765718;
srom_1(83891) <= 9196173;
srom_1(83892) <= 8622842;
srom_1(83893) <= 8048412;
srom_1(83894) <= 7475577;
srom_1(83895) <= 6907023;
srom_1(83896) <= 6345418;
srom_1(83897) <= 5793393;
srom_1(83898) <= 5253539;
srom_1(83899) <= 4728385;
srom_1(83900) <= 4220396;
srom_1(83901) <= 3731953;
srom_1(83902) <= 3265347;
srom_1(83903) <= 2822765;
srom_1(83904) <= 2406284;
srom_1(83905) <= 2017856;
srom_1(83906) <= 1659302;
srom_1(83907) <= 1332304;
srom_1(83908) <= 1038396;
srom_1(83909) <= 778955;
srom_1(83910) <= 555199;
srom_1(83911) <= 368176;
srom_1(83912) <= 218764;
srom_1(83913) <= 107663;
srom_1(83914) <= 35394;
srom_1(83915) <= 2297;
srom_1(83916) <= 8525;
srom_1(83917) <= 54051;
srom_1(83918) <= 138660;
srom_1(83919) <= 261956;
srom_1(83920) <= 423361;
srom_1(83921) <= 622117;
srom_1(83922) <= 857294;
srom_1(83923) <= 1127787;
srom_1(83924) <= 1432328;
srom_1(83925) <= 1769490;
srom_1(83926) <= 2137692;
srom_1(83927) <= 2535206;
srom_1(83928) <= 2960168;
srom_1(83929) <= 3410587;
srom_1(83930) <= 3884349;
srom_1(83931) <= 4379233;
srom_1(83932) <= 4892918;
srom_1(83933) <= 5422996;
srom_1(83934) <= 5966981;
srom_1(83935) <= 6522321;
srom_1(83936) <= 7086413;
srom_1(83937) <= 7656612;
srom_1(83938) <= 8230243;
srom_1(83939) <= 8804617;
srom_1(83940) <= 9377040;
srom_1(83941) <= 9944828;
srom_1(83942) <= 10505318;
srom_1(83943) <= 11055882;
srom_1(83944) <= 11593938;
srom_1(83945) <= 12116964;
srom_1(83946) <= 12622506;
srom_1(83947) <= 13108194;
srom_1(83948) <= 13571750;
srom_1(83949) <= 14011000;
srom_1(83950) <= 14423885;
srom_1(83951) <= 14808469;
srom_1(83952) <= 15162948;
srom_1(83953) <= 15485659;
srom_1(83954) <= 15775090;
srom_1(83955) <= 16029883;
srom_1(83956) <= 16248844;
srom_1(83957) <= 16430945;
srom_1(83958) <= 16575333;
srom_1(83959) <= 16681331;
srom_1(83960) <= 16748441;
srom_1(83961) <= 16776349;
srom_1(83962) <= 16764924;
srom_1(83963) <= 16714220;
srom_1(83964) <= 16624474;
srom_1(83965) <= 16496107;
srom_1(83966) <= 16329721;
srom_1(83967) <= 16126097;
srom_1(83968) <= 15886189;
srom_1(83969) <= 15611122;
srom_1(83970) <= 15302186;
srom_1(83971) <= 14960830;
srom_1(83972) <= 14588655;
srom_1(83973) <= 14187406;
srom_1(83974) <= 13758964;
srom_1(83975) <= 13305338;
srom_1(83976) <= 12828657;
srom_1(83977) <= 12331154;
srom_1(83978) <= 11815164;
srom_1(83979) <= 11283105;
srom_1(83980) <= 10737473;
srom_1(83981) <= 10180826;
srom_1(83982) <= 9615775;
srom_1(83983) <= 9044969;
srom_1(83984) <= 8471085;
srom_1(83985) <= 7896815;
srom_1(83986) <= 7324851;
srom_1(83987) <= 6757875;
srom_1(83988) <= 6198546;
srom_1(83989) <= 5649487;
srom_1(83990) <= 5113273;
srom_1(83991) <= 4592418;
srom_1(83992) <= 4089364;
srom_1(83993) <= 3606472;
srom_1(83994) <= 3146004;
srom_1(83995) <= 2710120;
srom_1(83996) <= 2300865;
srom_1(83997) <= 1920158;
srom_1(83998) <= 1569783;
srom_1(83999) <= 1251384;
srom_1(84000) <= 966454;
srom_1(84001) <= 716329;
srom_1(84002) <= 502182;
srom_1(84003) <= 325017;
srom_1(84004) <= 185665;
srom_1(84005) <= 84780;
srom_1(84006) <= 22834;
srom_1(84007) <= 118;
srom_1(84008) <= 16738;
srom_1(84009) <= 72617;
srom_1(84010) <= 167493;
srom_1(84011) <= 300920;
srom_1(84012) <= 472273;
srom_1(84013) <= 680748;
srom_1(84014) <= 925369;
srom_1(84015) <= 1204987;
srom_1(84016) <= 1518291;
srom_1(84017) <= 1863813;
srom_1(84018) <= 2239932;
srom_1(84019) <= 2644884;
srom_1(84020) <= 3076770;
srom_1(84021) <= 3533565;
srom_1(84022) <= 4013127;
srom_1(84023) <= 4513208;
srom_1(84024) <= 5031461;
srom_1(84025) <= 5565457;
srom_1(84026) <= 6112692;
srom_1(84027) <= 6670600;
srom_1(84028) <= 7236564;
srom_1(84029) <= 7807930;
srom_1(84030) <= 8382019;
srom_1(84031) <= 8956139;
srom_1(84032) <= 9527598;
srom_1(84033) <= 10093715;
srom_1(84034) <= 10651837;
srom_1(84035) <= 11199346;
srom_1(84036) <= 11733674;
srom_1(84037) <= 12252316;
srom_1(84038) <= 12752839;
srom_1(84039) <= 13232898;
srom_1(84040) <= 13690240;
srom_1(84041) <= 14122720;
srom_1(84042) <= 14528312;
srom_1(84043) <= 14905112;
srom_1(84044) <= 15251354;
srom_1(84045) <= 15565414;
srom_1(84046) <= 15845820;
srom_1(84047) <= 16091256;
srom_1(84048) <= 16300572;
srom_1(84049) <= 16472786;
srom_1(84050) <= 16607091;
srom_1(84051) <= 16702856;
srom_1(84052) <= 16759633;
srom_1(84053) <= 16777155;
srom_1(84054) <= 16755340;
srom_1(84055) <= 16694291;
srom_1(84056) <= 16594294;
srom_1(84057) <= 16455818;
srom_1(84058) <= 16279511;
srom_1(84059) <= 16066201;
srom_1(84060) <= 15816889;
srom_1(84061) <= 15532743;
srom_1(84062) <= 15215095;
srom_1(84063) <= 14865436;
srom_1(84064) <= 14485404;
srom_1(84065) <= 14076783;
srom_1(84066) <= 13641488;
srom_1(84067) <= 13181560;
srom_1(84068) <= 12699156;
srom_1(84069) <= 12196539;
srom_1(84070) <= 11676065;
srom_1(84071) <= 11140175;
srom_1(84072) <= 10591382;
srom_1(84073) <= 10032260;
srom_1(84074) <= 9465430;
srom_1(84075) <= 8893550;
srom_1(84076) <= 8319302;
srom_1(84077) <= 7745379;
srom_1(84078) <= 7174473;
srom_1(84079) <= 6609260;
srom_1(84080) <= 6052391;
srom_1(84081) <= 5506478;
srom_1(84082) <= 4974079;
srom_1(84083) <= 4457693;
srom_1(84084) <= 3959740;
srom_1(84085) <= 3482555;
srom_1(84086) <= 3028377;
srom_1(84087) <= 2599335;
srom_1(84088) <= 2197440;
srom_1(84089) <= 1824578;
srom_1(84090) <= 1482497;
srom_1(84091) <= 1172801;
srom_1(84092) <= 896943;
srom_1(84093) <= 656215;
srom_1(84094) <= 451747;
srom_1(84095) <= 284498;
srom_1(84096) <= 155252;
srom_1(84097) <= 64615;
srom_1(84098) <= 13012;
srom_1(84099) <= 685;
srom_1(84100) <= 27692;
srom_1(84101) <= 93906;
srom_1(84102) <= 199017;
srom_1(84103) <= 342531;
srom_1(84104) <= 523777;
srom_1(84105) <= 741903;
srom_1(84106) <= 995887;
srom_1(84107) <= 1284539;
srom_1(84108) <= 1606503;
srom_1(84109) <= 1960272;
srom_1(84110) <= 2344185;
srom_1(84111) <= 2756442;
srom_1(84112) <= 3195111;
srom_1(84113) <= 3658133;
srom_1(84114) <= 4143339;
srom_1(84115) <= 4648452;
srom_1(84116) <= 5171103;
srom_1(84117) <= 5708843;
srom_1(84118) <= 6259149;
srom_1(84119) <= 6819441;
srom_1(84120) <= 7387091;
srom_1(84121) <= 7959438;
srom_1(84122) <= 8533797;
srom_1(84123) <= 9107476;
srom_1(84124) <= 9677783;
srom_1(84125) <= 10242045;
srom_1(84126) <= 10797615;
srom_1(84127) <= 11341889;
srom_1(84128) <= 11872314;
srom_1(84129) <= 12386403;
srom_1(84130) <= 12881744;
srom_1(84131) <= 13356016;
srom_1(84132) <= 13806994;
srom_1(84133) <= 14232563;
srom_1(84134) <= 14630728;
srom_1(84135) <= 14999621;
srom_1(84136) <= 15337513;
srom_1(84137) <= 15642819;
srom_1(84138) <= 15914108;
srom_1(84139) <= 16150107;
srom_1(84140) <= 16349710;
srom_1(84141) <= 16511980;
srom_1(84142) <= 16636157;
srom_1(84143) <= 16721659;
srom_1(84144) <= 16768084;
srom_1(84145) <= 16775214;
srom_1(84146) <= 16743017;
srom_1(84147) <= 16671644;
srom_1(84148) <= 16561428;
srom_1(84149) <= 16412887;
srom_1(84150) <= 16226718;
srom_1(84151) <= 16003793;
srom_1(84152) <= 15745157;
srom_1(84153) <= 15452025;
srom_1(84154) <= 15125769;
srom_1(84155) <= 14767921;
srom_1(84156) <= 14380158;
srom_1(84157) <= 13964298;
srom_1(84158) <= 13522292;
srom_1(84159) <= 13056212;
srom_1(84160) <= 12568245;
srom_1(84161) <= 12060678;
srom_1(84162) <= 11535891;
srom_1(84163) <= 10996345;
srom_1(84164) <= 10444571;
srom_1(84165) <= 9883156;
srom_1(84166) <= 9314732;
srom_1(84167) <= 8741965;
srom_1(84168) <= 8167541;
srom_1(84169) <= 7594154;
srom_1(84170) <= 7024493;
srom_1(84171) <= 6461228;
srom_1(84172) <= 5907001;
srom_1(84173) <= 5364412;
srom_1(84174) <= 4836004;
srom_1(84175) <= 4324255;
srom_1(84176) <= 3831565;
srom_1(84177) <= 3360245;
srom_1(84178) <= 2912505;
srom_1(84179) <= 2490444;
srom_1(84180) <= 2096042;
srom_1(84181) <= 1731147;
srom_1(84182) <= 1397472;
srom_1(84183) <= 1096580;
srom_1(84184) <= 829883;
srom_1(84185) <= 598632;
srom_1(84186) <= 403911;
srom_1(84187) <= 246632;
srom_1(84188) <= 127534;
srom_1(84189) <= 47176;
srom_1(84190) <= 5932;
srom_1(84191) <= 3999;
srom_1(84192) <= 41383;
srom_1(84193) <= 117911;
srom_1(84194) <= 233222;
srom_1(84195) <= 386777;
srom_1(84196) <= 577856;
srom_1(84197) <= 805561;
srom_1(84198) <= 1068826;
srom_1(84199) <= 1366416;
srom_1(84200) <= 1696936;
srom_1(84201) <= 2058835;
srom_1(84202) <= 2450417;
srom_1(84203) <= 2869844;
srom_1(84204) <= 3315152;
srom_1(84205) <= 3784250;
srom_1(84206) <= 4274940;
srom_1(84207) <= 4784920;
srom_1(84208) <= 5311799;
srom_1(84209) <= 5853106;
srom_1(84210) <= 6406303;
srom_1(84211) <= 6968796;
srom_1(84212) <= 7537947;
srom_1(84213) <= 8111087;
srom_1(84214) <= 8685528;
srom_1(84215) <= 9258577;
srom_1(84216) <= 9827546;
srom_1(84217) <= 10389768;
srom_1(84218) <= 10942605;
srom_1(84219) <= 11483466;
srom_1(84220) <= 12009814;
srom_1(84221) <= 12519181;
srom_1(84222) <= 13009178;
srom_1(84223) <= 13477508;
srom_1(84224) <= 13921974;
srom_1(84225) <= 14340492;
srom_1(84226) <= 14731100;
srom_1(84227) <= 15091966;
srom_1(84228) <= 15421397;
srom_1(84229) <= 15717849;
srom_1(84230) <= 15979932;
srom_1(84231) <= 16206417;
srom_1(84232) <= 16396241;
srom_1(84233) <= 16548515;
srom_1(84234) <= 16662524;
srom_1(84235) <= 16737733;
srom_1(84236) <= 16773791;
srom_1(84237) <= 16770528;
srom_1(84238) <= 16727959;
srom_1(84239) <= 16646284;
srom_1(84240) <= 16525886;
srom_1(84241) <= 16367330;
srom_1(84242) <= 16171358;
srom_1(84243) <= 15938890;
srom_1(84244) <= 15671017;
srom_1(84245) <= 15368994;
srom_1(84246) <= 15034237;
srom_1(84247) <= 14668317;
srom_1(84248) <= 14272949;
srom_1(84249) <= 13849987;
srom_1(84250) <= 13401416;
srom_1(84251) <= 12929337;
srom_1(84252) <= 12435965;
srom_1(84253) <= 11923614;
srom_1(84254) <= 11394686;
srom_1(84255) <= 10851661;
srom_1(84256) <= 10297086;
srom_1(84257) <= 9733562;
srom_1(84258) <= 9163731;
srom_1(84259) <= 8590265;
srom_1(84260) <= 8015853;
srom_1(84261) <= 7443189;
srom_1(84262) <= 6874959;
srom_1(84263) <= 6313827;
srom_1(84264) <= 5762424;
srom_1(84265) <= 5223336;
srom_1(84266) <= 4699091;
srom_1(84267) <= 4192148;
srom_1(84268) <= 3704883;
srom_1(84269) <= 3239582;
srom_1(84270) <= 2798426;
srom_1(84271) <= 2383485;
srom_1(84272) <= 1996703;
srom_1(84273) <= 1639896;
srom_1(84274) <= 1314735;
srom_1(84275) <= 1022747;
srom_1(84276) <= 765299;
srom_1(84277) <= 543600;
srom_1(84278) <= 358688;
srom_1(84279) <= 211432;
srom_1(84280) <= 102521;
srom_1(84281) <= 32467;
srom_1(84282) <= 1597;
srom_1(84283) <= 10057;
srom_1(84284) <= 57807;
srom_1(84285) <= 144623;
srom_1(84286) <= 270098;
srom_1(84287) <= 433643;
srom_1(84288) <= 634492;
srom_1(84289) <= 871702;
srom_1(84290) <= 1144162;
srom_1(84291) <= 1450593;
srom_1(84292) <= 1789559;
srom_1(84293) <= 2159471;
srom_1(84294) <= 2558593;
srom_1(84295) <= 2985054;
srom_1(84296) <= 3436854;
srom_1(84297) <= 3911874;
srom_1(84298) <= 4407888;
srom_1(84299) <= 4922568;
srom_1(84300) <= 5453502;
srom_1(84301) <= 5998199;
srom_1(84302) <= 6554106;
srom_1(84303) <= 7118616;
srom_1(84304) <= 7689081;
srom_1(84305) <= 8262826;
srom_1(84306) <= 8837161;
srom_1(84307) <= 9409393;
srom_1(84308) <= 9976838;
srom_1(84309) <= 10536835;
srom_1(84310) <= 11086758;
srom_1(84311) <= 11624029;
srom_1(84312) <= 12146128;
srom_1(84313) <= 12650606;
srom_1(84314) <= 13135099;
srom_1(84315) <= 13597333;
srom_1(84316) <= 14035143;
srom_1(84317) <= 14446473;
srom_1(84318) <= 14829396;
srom_1(84319) <= 15182116;
srom_1(84320) <= 15502979;
srom_1(84321) <= 15790480;
srom_1(84322) <= 16043271;
srom_1(84323) <= 16260167;
srom_1(84324) <= 16440151;
srom_1(84325) <= 16582378;
srom_1(84326) <= 16686181;
srom_1(84327) <= 16751075;
srom_1(84328) <= 16776754;
srom_1(84329) <= 16763098;
srom_1(84330) <= 16710171;
srom_1(84331) <= 16618221;
srom_1(84332) <= 16487680;
srom_1(84333) <= 16319160;
srom_1(84334) <= 16113450;
srom_1(84335) <= 15871516;
srom_1(84336) <= 15594493;
srom_1(84337) <= 15283678;
srom_1(84338) <= 14940530;
srom_1(84339) <= 14566658;
srom_1(84340) <= 14163814;
srom_1(84341) <= 13733889;
srom_1(84342) <= 13278898;
srom_1(84343) <= 12800975;
srom_1(84344) <= 12302360;
srom_1(84345) <= 11785393;
srom_1(84346) <= 11252497;
srom_1(84347) <= 10706171;
srom_1(84348) <= 10148977;
srom_1(84349) <= 9583528;
srom_1(84350) <= 9012476;
srom_1(84351) <= 8438499;
srom_1(84352) <= 7864287;
srom_1(84353) <= 7292534;
srom_1(84354) <= 6725921;
srom_1(84355) <= 6167105;
srom_1(84356) <= 5618706;
srom_1(84357) <= 5083296;
srom_1(84358) <= 4563386;
srom_1(84359) <= 4061414;
srom_1(84360) <= 3579734;
srom_1(84361) <= 3120604;
srom_1(84362) <= 2686177;
srom_1(84363) <= 2278491;
srom_1(84364) <= 1899458;
srom_1(84365) <= 1550854;
srom_1(84366) <= 1234315;
srom_1(84367) <= 951325;
srom_1(84368) <= 703211;
srom_1(84369) <= 491136;
srom_1(84370) <= 316095;
srom_1(84371) <= 178909;
srom_1(84372) <= 80221;
srom_1(84373) <= 20494;
srom_1(84374) <= 8;
srom_1(84375) <= 18859;
srom_1(84376) <= 76959;
srom_1(84377) <= 174034;
srom_1(84378) <= 309631;
srom_1(84379) <= 483113;
srom_1(84380) <= 693666;
srom_1(84381) <= 940304;
srom_1(84382) <= 1221869;
srom_1(84383) <= 1537041;
srom_1(84384) <= 1884343;
srom_1(84385) <= 2262146;
srom_1(84386) <= 2668678;
srom_1(84387) <= 3102032;
srom_1(84388) <= 3560177;
srom_1(84389) <= 4040964;
srom_1(84390) <= 4542139;
srom_1(84391) <= 5061351;
srom_1(84392) <= 5596166;
srom_1(84393) <= 6144075;
srom_1(84394) <= 6702510;
srom_1(84395) <= 7268851;
srom_1(84396) <= 7840444;
srom_1(84397) <= 8414607;
srom_1(84398) <= 8988648;
srom_1(84399) <= 9559875;
srom_1(84400) <= 10125610;
srom_1(84401) <= 10683199;
srom_1(84402) <= 11230028;
srom_1(84403) <= 11763533;
srom_1(84404) <= 12281212;
srom_1(84405) <= 12780637;
srom_1(84406) <= 13259466;
srom_1(84407) <= 13715454;
srom_1(84408) <= 14146463;
srom_1(84409) <= 14550471;
srom_1(84410) <= 14925583;
srom_1(84411) <= 15270042;
srom_1(84412) <= 15582232;
srom_1(84413) <= 15860688;
srom_1(84414) <= 16104104;
srom_1(84415) <= 16311341;
srom_1(84416) <= 16481424;
srom_1(84417) <= 16613558;
srom_1(84418) <= 16707122;
srom_1(84419) <= 16761678;
srom_1(84420) <= 16776970;
srom_1(84421) <= 16752925;
srom_1(84422) <= 16689658;
srom_1(84423) <= 16587464;
srom_1(84424) <= 16446823;
srom_1(84425) <= 16268394;
srom_1(84426) <= 16053014;
srom_1(84427) <= 15801693;
srom_1(84428) <= 15515609;
srom_1(84429) <= 15196105;
srom_1(84430) <= 14844677;
srom_1(84431) <= 14462975;
srom_1(84432) <= 14052789;
srom_1(84433) <= 13616040;
srom_1(84434) <= 13154779;
srom_1(84435) <= 12671168;
srom_1(84436) <= 12167474;
srom_1(84437) <= 11646059;
srom_1(84438) <= 11109370;
srom_1(84439) <= 10559922;
srom_1(84440) <= 10000291;
srom_1(84441) <= 9433103;
srom_1(84442) <= 8861017;
srom_1(84443) <= 8286716;
srom_1(84444) <= 7712892;
srom_1(84445) <= 7142238;
srom_1(84446) <= 6577427;
srom_1(84447) <= 6021110;
srom_1(84448) <= 5475895;
srom_1(84449) <= 4944339;
srom_1(84450) <= 4428934;
srom_1(84451) <= 3932098;
srom_1(84452) <= 3456159;
srom_1(84453) <= 3003350;
srom_1(84454) <= 2575795;
srom_1(84455) <= 2175498;
srom_1(84456) <= 1804336;
srom_1(84457) <= 1464051;
srom_1(84458) <= 1156237;
srom_1(84459) <= 882338;
srom_1(84460) <= 643638;
srom_1(84461) <= 441257;
srom_1(84462) <= 276144;
srom_1(84463) <= 149074;
srom_1(84464) <= 60641;
srom_1(84465) <= 11261;
srom_1(84466) <= 1165;
srom_1(84467) <= 30401;
srom_1(84468) <= 98831;
srom_1(84469) <= 206135;
srom_1(84470) <= 351809;
srom_1(84471) <= 535171;
srom_1(84472) <= 755360;
srom_1(84473) <= 1011344;
srom_1(84474) <= 1301922;
srom_1(84475) <= 1625733;
srom_1(84476) <= 1981257;
srom_1(84477) <= 2366827;
srom_1(84478) <= 2780635;
srom_1(84479) <= 3220741;
srom_1(84480) <= 3685081;
srom_1(84481) <= 4171477;
srom_1(84482) <= 4677649;
srom_1(84483) <= 5201223;
srom_1(84484) <= 5739744;
srom_1(84485) <= 6290686;
srom_1(84486) <= 6851465;
srom_1(84487) <= 7419454;
srom_1(84488) <= 7991986;
srom_1(84489) <= 8566379;
srom_1(84490) <= 9139938;
srom_1(84491) <= 9709974;
srom_1(84492) <= 10273813;
srom_1(84493) <= 10828812;
srom_1(84494) <= 11372368;
srom_1(84495) <= 11901933;
srom_1(84496) <= 12415022;
srom_1(84497) <= 12909229;
srom_1(84498) <= 13382238;
srom_1(84499) <= 13831830;
srom_1(84500) <= 14255897;
srom_1(84501) <= 14652451;
srom_1(84502) <= 15019631;
srom_1(84503) <= 15355715;
srom_1(84504) <= 15659129;
srom_1(84505) <= 15928449;
srom_1(84506) <= 16162411;
srom_1(84507) <= 16359920;
srom_1(84508) <= 16520049;
srom_1(84509) <= 16642046;
srom_1(84510) <= 16725340;
srom_1(84511) <= 16769540;
srom_1(84512) <= 16774440;
srom_1(84513) <= 16740015;
srom_1(84514) <= 16666427;
srom_1(84515) <= 16554022;
srom_1(84516) <= 16403327;
srom_1(84517) <= 16215048;
srom_1(84518) <= 15990068;
srom_1(84519) <= 15729442;
srom_1(84520) <= 15434392;
srom_1(84521) <= 15106302;
srom_1(84522) <= 14746711;
srom_1(84523) <= 14357304;
srom_1(84524) <= 13939908;
srom_1(84525) <= 13496481;
srom_1(84526) <= 13029100;
srom_1(84527) <= 12539959;
srom_1(84528) <= 12031350;
srom_1(84529) <= 11505660;
srom_1(84530) <= 10965352;
srom_1(84531) <= 10412962;
srom_1(84532) <= 9851078;
srom_1(84533) <= 9282336;
srom_1(84534) <= 8709404;
srom_1(84535) <= 8134967;
srom_1(84536) <= 7561719;
srom_1(84537) <= 6992349;
srom_1(84538) <= 6429527;
srom_1(84539) <= 5875891;
srom_1(84540) <= 5334038;
srom_1(84541) <= 4806509;
srom_1(84542) <= 4295778;
srom_1(84543) <= 3804240;
srom_1(84544) <= 3334199;
srom_1(84545) <= 2887860;
srom_1(84546) <= 2467316;
srom_1(84547) <= 2074539;
srom_1(84548) <= 1711371;
srom_1(84549) <= 1379515;
srom_1(84550) <= 1080526;
srom_1(84551) <= 815808;
srom_1(84552) <= 586601;
srom_1(84553) <= 393981;
srom_1(84554) <= 238850;
srom_1(84555) <= 121936;
srom_1(84556) <= 43787;
srom_1(84557) <= 4770;
srom_1(84558) <= 5068;
srom_1(84559) <= 44679;
srom_1(84560) <= 123418;
srom_1(84561) <= 240915;
srom_1(84562) <= 396619;
srom_1(84563) <= 589800;
srom_1(84564) <= 819553;
srom_1(84565) <= 1084799;
srom_1(84566) <= 1384296;
srom_1(84567) <= 1716638;
srom_1(84568) <= 2080268;
srom_1(84569) <= 2473479;
srom_1(84570) <= 2894428;
srom_1(84571) <= 3341142;
srom_1(84572) <= 3811525;
srom_1(84573) <= 4303371;
srom_1(84574) <= 4814374;
srom_1(84575) <= 5342139;
srom_1(84576) <= 5884189;
srom_1(84577) <= 6437983;
srom_1(84578) <= 7000924;
srom_1(84579) <= 7570373;
srom_1(84580) <= 8143659;
srom_1(84581) <= 8718093;
srom_1(84582) <= 9290982;
srom_1(84583) <= 9859640;
srom_1(84584) <= 10421399;
srom_1(84585) <= 10973626;
srom_1(84586) <= 11513731;
srom_1(84587) <= 12039181;
srom_1(84588) <= 12547513;
srom_1(84589) <= 13036342;
srom_1(84590) <= 13503376;
srom_1(84591) <= 13946425;
srom_1(84592) <= 14363411;
srom_1(84593) <= 14752380;
srom_1(84594) <= 15111507;
srom_1(84595) <= 15439108;
srom_1(84596) <= 15733646;
srom_1(84597) <= 15993741;
srom_1(84598) <= 16218173;
srom_1(84599) <= 16405890;
srom_1(84600) <= 16556011;
srom_1(84601) <= 16667832;
srom_1(84602) <= 16740828;
srom_1(84603) <= 16774659;
srom_1(84604) <= 16769164;
srom_1(84605) <= 16724370;
srom_1(84606) <= 16640487;
srom_1(84607) <= 16517908;
srom_1(84608) <= 16357207;
srom_1(84609) <= 16159140;
srom_1(84610) <= 15924633;
srom_1(84611) <= 15654788;
srom_1(84612) <= 15350869;
srom_1(84613) <= 15014301;
srom_1(84614) <= 14646663;
srom_1(84615) <= 14249679;
srom_1(84616) <= 13825211;
srom_1(84617) <= 13375248;
srom_1(84618) <= 12901902;
srom_1(84619) <= 12407391;
srom_1(84620) <= 11894034;
srom_1(84621) <= 11364240;
srom_1(84622) <= 10820491;
srom_1(84623) <= 10265339;
srom_1(84624) <= 9701386;
srom_1(84625) <= 9131277;
srom_1(84626) <= 8557685;
srom_1(84627) <= 7983300;
srom_1(84628) <= 7410816;
srom_1(84629) <= 6842918;
srom_1(84630) <= 6282267;
srom_1(84631) <= 5731494;
srom_1(84632) <= 5193181;
srom_1(84633) <= 4669852;
srom_1(84634) <= 4163962;
srom_1(84635) <= 3677883;
srom_1(84636) <= 3213894;
srom_1(84637) <= 2774171;
srom_1(84638) <= 2360776;
srom_1(84639) <= 1975647;
srom_1(84640) <= 1620592;
srom_1(84641) <= 1297273;
srom_1(84642) <= 1007209;
srom_1(84643) <= 751758;
srom_1(84644) <= 532119;
srom_1(84645) <= 349322;
srom_1(84646) <= 204223;
srom_1(84647) <= 97505;
srom_1(84648) <= 29666;
srom_1(84649) <= 1025;
srom_1(84650) <= 11716;
srom_1(84651) <= 61689;
srom_1(84652) <= 150710;
srom_1(84653) <= 278362;
srom_1(84654) <= 444045;
srom_1(84655) <= 646983;
srom_1(84656) <= 886224;
srom_1(84657) <= 1160646;
srom_1(84658) <= 1468963;
srom_1(84659) <= 1809728;
srom_1(84660) <= 2181344;
srom_1(84661) <= 2582068;
srom_1(84662) <= 3010021;
srom_1(84663) <= 3463195;
srom_1(84664) <= 3939467;
srom_1(84665) <= 4436602;
srom_1(84666) <= 4952270;
srom_1(84667) <= 5484052;
srom_1(84668) <= 6029454;
srom_1(84669) <= 6585919;
srom_1(84670) <= 7150838;
srom_1(84671) <= 7721560;
srom_1(84672) <= 8295411;
srom_1(84673) <= 8869699;
srom_1(84674) <= 9441731;
srom_1(84675) <= 10008824;
srom_1(84676) <= 10568320;
srom_1(84677) <= 11117594;
srom_1(84678) <= 11654071;
srom_1(84679) <= 12175235;
srom_1(84680) <= 12678643;
srom_1(84681) <= 13161933;
srom_1(84682) <= 13622839;
srom_1(84683) <= 14059200;
srom_1(84684) <= 14468969;
srom_1(84685) <= 14850226;
srom_1(84686) <= 15201182;
srom_1(84687) <= 15520192;
srom_1(84688) <= 15805759;
srom_1(84689) <= 16056544;
srom_1(84690) <= 16271372;
srom_1(84691) <= 16449235;
srom_1(84692) <= 16589299;
srom_1(84693) <= 16690907;
srom_1(84694) <= 16753582;
srom_1(84695) <= 16777032;
srom_1(84696) <= 16761145;
srom_1(84697) <= 16705996;
srom_1(84698) <= 16611845;
srom_1(84699) <= 16479131;
srom_1(84700) <= 16308479;
srom_1(84701) <= 16100687;
srom_1(84702) <= 15856731;
srom_1(84703) <= 15577755;
srom_1(84704) <= 15265066;
srom_1(84705) <= 14920130;
srom_1(84706) <= 14544567;
srom_1(84707) <= 14140136;
srom_1(84708) <= 13708734;
srom_1(84709) <= 13252384;
srom_1(84710) <= 12773226;
srom_1(84711) <= 12273507;
srom_1(84712) <= 11755570;
srom_1(84713) <= 11221845;
srom_1(84714) <= 10674834;
srom_1(84715) <= 10117102;
srom_1(84716) <= 9551264;
srom_1(84717) <= 8979974;
srom_1(84718) <= 8405911;
srom_1(84719) <= 7831767;
srom_1(84720) <= 7260234;
srom_1(84721) <= 6693992;
srom_1(84722) <= 6135697;
srom_1(84723) <= 5587967;
srom_1(84724) <= 5053370;
srom_1(84725) <= 4534413;
srom_1(84726) <= 4033530;
srom_1(84727) <= 3553069;
srom_1(84728) <= 3095283;
srom_1(84729) <= 2662320;
srom_1(84730) <= 2256209;
srom_1(84731) <= 1878855;
srom_1(84732) <= 1532028;
srom_1(84733) <= 1217353;
srom_1(84734) <= 936307;
srom_1(84735) <= 690208;
srom_1(84736) <= 480209;
srom_1(84737) <= 307295;
srom_1(84738) <= 172277;
srom_1(84739) <= 75788;
srom_1(84740) <= 18281;
srom_1(84741) <= 25;
srom_1(84742) <= 21106;
srom_1(84743) <= 81425;
srom_1(84744) <= 180700;
srom_1(84745) <= 318464;
srom_1(84746) <= 494072;
srom_1(84747) <= 706700;
srom_1(84748) <= 955351;
srom_1(84749) <= 1238859;
srom_1(84750) <= 1555895;
srom_1(84751) <= 1904972;
srom_1(84752) <= 2284453;
srom_1(84753) <= 2692558;
srom_1(84754) <= 3127374;
srom_1(84755) <= 3586861;
srom_1(84756) <= 4068866;
srom_1(84757) <= 4571128;
srom_1(84758) <= 5091291;
srom_1(84759) <= 5626916;
srom_1(84760) <= 6175491;
srom_1(84761) <= 6734445;
srom_1(84762) <= 7301156;
srom_1(84763) <= 7872966;
srom_1(84764) <= 8447194;
srom_1(84765) <= 9021148;
srom_1(84766) <= 9592135;
srom_1(84767) <= 10157478;
srom_1(84768) <= 10714527;
srom_1(84769) <= 11260668;
srom_1(84770) <= 11793342;
srom_1(84771) <= 12310049;
srom_1(84772) <= 12808368;
srom_1(84773) <= 13285961;
srom_1(84774) <= 13740588;
srom_1(84775) <= 14170118;
srom_1(84776) <= 14572537;
srom_1(84777) <= 14945957;
srom_1(84778) <= 15288627;
srom_1(84779) <= 15598941;
srom_1(84780) <= 15875443;
srom_1(84781) <= 16116836;
srom_1(84782) <= 16321990;
srom_1(84783) <= 16489941;
srom_1(84784) <= 16619902;
srom_1(84785) <= 16711263;
srom_1(84786) <= 16763597;
srom_1(84787) <= 16776658;
srom_1(84788) <= 16750384;
srom_1(84789) <= 16684899;
srom_1(84790) <= 16580510;
srom_1(84791) <= 16437706;
srom_1(84792) <= 16257157;
srom_1(84793) <= 16039710;
srom_1(84794) <= 15786384;
srom_1(84795) <= 15498368;
srom_1(84796) <= 15177011;
srom_1(84797) <= 14823821;
srom_1(84798) <= 14440455;
srom_1(84799) <= 14028709;
srom_1(84800) <= 13590514;
srom_1(84801) <= 13127926;
srom_1(84802) <= 12643114;
srom_1(84803) <= 12138351;
srom_1(84804) <= 11616004;
srom_1(84805) <= 11078523;
srom_1(84806) <= 10528428;
srom_1(84807) <= 9968299;
srom_1(84808) <= 9400761;
srom_1(84809) <= 8828478;
srom_1(84810) <= 8254131;
srom_1(84811) <= 7680416;
srom_1(84812) <= 7110021;
srom_1(84813) <= 6545622;
srom_1(84814) <= 5989865;
srom_1(84815) <= 5445357;
srom_1(84816) <= 4914651;
srom_1(84817) <= 4400235;
srom_1(84818) <= 3904523;
srom_1(84819) <= 3429837;
srom_1(84820) <= 2978405;
srom_1(84821) <= 2552343;
srom_1(84822) <= 2153650;
srom_1(84823) <= 1784194;
srom_1(84824) <= 1445709;
srom_1(84825) <= 1139781;
srom_1(84826) <= 867846;
srom_1(84827) <= 631178;
srom_1(84828) <= 430887;
srom_1(84829) <= 267913;
srom_1(84830) <= 143020;
srom_1(84831) <= 56792;
srom_1(84832) <= 9636;
srom_1(84833) <= 1772;
srom_1(84834) <= 33236;
srom_1(84835) <= 103881;
srom_1(84836) <= 213377;
srom_1(84837) <= 361208;
srom_1(84838) <= 546683;
srom_1(84839) <= 768932;
srom_1(84840) <= 1026912;
srom_1(84841) <= 1319413;
srom_1(84842) <= 1645064;
srom_1(84843) <= 2002338;
srom_1(84844) <= 2389560;
srom_1(84845) <= 2804913;
srom_1(84846) <= 3246449;
srom_1(84847) <= 3712100;
srom_1(84848) <= 4199679;
srom_1(84849) <= 4706903;
srom_1(84850) <= 5231391;
srom_1(84851) <= 5770684;
srom_1(84852) <= 6322254;
srom_1(84853) <= 6883513;
srom_1(84854) <= 7451830;
srom_1(84855) <= 8024541;
srom_1(84856) <= 8598958;
srom_1(84857) <= 9172389;
srom_1(84858) <= 9742145;
srom_1(84859) <= 10305553;
srom_1(84860) <= 10859972;
srom_1(84861) <= 11402802;
srom_1(84862) <= 11931498;
srom_1(84863) <= 12443580;
srom_1(84864) <= 12936646;
srom_1(84865) <= 13408385;
srom_1(84866) <= 13856585;
srom_1(84867) <= 14279143;
srom_1(84868) <= 14674079;
srom_1(84869) <= 15039540;
srom_1(84870) <= 15373813;
srom_1(84871) <= 15675329;
srom_1(84872) <= 15942676;
srom_1(84873) <= 16174599;
srom_1(84874) <= 16370010;
srom_1(84875) <= 16527994;
srom_1(84876) <= 16647810;
srom_1(84877) <= 16728896;
srom_1(84878) <= 16770871;
srom_1(84879) <= 16773538;
srom_1(84880) <= 16736886;
srom_1(84881) <= 16661086;
srom_1(84882) <= 16546494;
srom_1(84883) <= 16393646;
srom_1(84884) <= 16203260;
srom_1(84885) <= 15976228;
srom_1(84886) <= 15713616;
srom_1(84887) <= 15416653;
srom_1(84888) <= 15086734;
srom_1(84889) <= 14725406;
srom_1(84890) <= 14334361;
srom_1(84891) <= 13915435;
srom_1(84892) <= 13470592;
srom_1(84893) <= 13001918;
srom_1(84894) <= 12511610;
srom_1(84895) <= 12001968;
srom_1(84896) <= 11475382;
srom_1(84897) <= 10934321;
srom_1(84898) <= 10381322;
srom_1(84899) <= 9818978;
srom_1(84900) <= 9249927;
srom_1(84901) <= 8676837;
srom_1(84902) <= 8102396;
srom_1(84903) <= 7529296;
srom_1(84904) <= 6960226;
srom_1(84905) <= 6397855;
srom_1(84906) <= 5844818;
srom_1(84907) <= 5303711;
srom_1(84908) <= 4777069;
srom_1(84909) <= 4267363;
srom_1(84910) <= 3776984;
srom_1(84911) <= 3308229;
srom_1(84912) <= 2863298;
srom_1(84913) <= 2444278;
srom_1(84914) <= 2053132;
srom_1(84915) <= 1691696;
srom_1(84916) <= 1361663;
srom_1(84917) <= 1064583;
srom_1(84918) <= 801847;
srom_1(84919) <= 574688;
srom_1(84920) <= 384171;
srom_1(84921) <= 231190;
srom_1(84922) <= 116462;
srom_1(84923) <= 40525;
srom_1(84924) <= 3735;
srom_1(84925) <= 6264;
srom_1(84926) <= 48101;
srom_1(84927) <= 129049;
srom_1(84928) <= 248730;
srom_1(84929) <= 406581;
srom_1(84930) <= 601862;
srom_1(84931) <= 833659;
srom_1(84932) <= 1100883;
srom_1(84933) <= 1402281;
srom_1(84934) <= 1736441;
srom_1(84935) <= 2101795;
srom_1(84936) <= 2496631;
srom_1(84937) <= 2919095;
srom_1(84938) <= 3367208;
srom_1(84939) <= 3838869;
srom_1(84940) <= 4331864;
srom_1(84941) <= 4843883;
srom_1(84942) <= 5372524;
srom_1(84943) <= 5915309;
srom_1(84944) <= 6469692;
srom_1(84945) <= 7033074;
srom_1(84946) <= 7602812;
srom_1(84947) <= 8176234;
srom_1(84948) <= 8750653;
srom_1(84949) <= 9323374;
srom_1(84950) <= 9891711;
srom_1(84951) <= 10453000;
srom_1(84952) <= 11004609;
srom_1(84953) <= 11543950;
srom_1(84954) <= 12068494;
srom_1(84955) <= 12575782;
srom_1(84956) <= 13063435;
srom_1(84957) <= 13529167;
srom_1(84958) <= 13970792;
srom_1(84959) <= 14386240;
srom_1(84960) <= 14773564;
srom_1(84961) <= 15130946;
srom_1(84962) <= 15456712;
srom_1(84963) <= 15749332;
srom_1(84964) <= 16007435;
srom_1(84965) <= 16229812;
srom_1(84966) <= 16415418;
srom_1(84967) <= 16563383;
srom_1(84968) <= 16673014;
srom_1(84969) <= 16743797;
srom_1(84970) <= 16775400;
srom_1(84971) <= 16767674;
srom_1(84972) <= 16720655;
srom_1(84973) <= 16634565;
srom_1(84974) <= 16509806;
srom_1(84975) <= 16346965;
srom_1(84976) <= 16146804;
srom_1(84977) <= 15910262;
srom_1(84978) <= 15638449;
srom_1(84979) <= 15332638;
srom_1(84980) <= 14994265;
srom_1(84981) <= 14624915;
srom_1(84982) <= 14226321;
srom_1(84983) <= 13800352;
srom_1(84984) <= 13349006;
srom_1(84985) <= 12874399;
srom_1(84986) <= 12378756;
srom_1(84987) <= 11864402;
srom_1(84988) <= 11333748;
srom_1(84989) <= 10789285;
srom_1(84990) <= 10233563;
srom_1(84991) <= 9669190;
srom_1(84992) <= 9098811;
srom_1(84993) <= 8525103;
srom_1(84994) <= 7950754;
srom_1(84995) <= 7378458;
srom_1(84996) <= 6810900;
srom_1(84997) <= 6250739;
srom_1(84998) <= 5700604;
srom_1(84999) <= 5163074;
srom_1(85000) <= 4640670;
srom_1(85001) <= 4135841;
srom_1(85002) <= 3650954;
srom_1(85003) <= 3188285;
srom_1(85004) <= 2750001;
srom_1(85005) <= 2338158;
srom_1(85006) <= 1954688;
srom_1(85007) <= 1601389;
srom_1(85008) <= 1279918;
srom_1(85009) <= 991782;
srom_1(85010) <= 738332;
srom_1(85011) <= 520756;
srom_1(85012) <= 340076;
srom_1(85013) <= 197138;
srom_1(85014) <= 92613;
srom_1(85015) <= 26990;
srom_1(85016) <= 578;
srom_1(85017) <= 13501;
srom_1(85018) <= 65697;
srom_1(85019) <= 156922;
srom_1(85020) <= 286748;
srom_1(85021) <= 454567;
srom_1(85022) <= 659591;
srom_1(85023) <= 900859;
srom_1(85024) <= 1177240;
srom_1(85025) <= 1487437;
srom_1(85026) <= 1829996;
srom_1(85027) <= 2203311;
srom_1(85028) <= 2605631;
srom_1(85029) <= 3035069;
srom_1(85030) <= 3489612;
srom_1(85031) <= 3967127;
srom_1(85032) <= 4465377;
srom_1(85033) <= 4982024;
srom_1(85034) <= 5514646;
srom_1(85035) <= 6060744;
srom_1(85036) <= 6617759;
srom_1(85037) <= 7183078;
srom_1(85038) <= 7754050;
srom_1(85039) <= 8327998;
srom_1(85040) <= 8902230;
srom_1(85041) <= 9474053;
srom_1(85042) <= 10040786;
srom_1(85043) <= 10599772;
srom_1(85044) <= 11148389;
srom_1(85045) <= 11684064;
srom_1(85046) <= 12204285;
srom_1(85047) <= 12706614;
srom_1(85048) <= 13188694;
srom_1(85049) <= 13648265;
srom_1(85050) <= 14083171;
srom_1(85051) <= 14491374;
srom_1(85052) <= 14870959;
srom_1(85053) <= 15220145;
srom_1(85054) <= 15537296;
srom_1(85055) <= 15820925;
srom_1(85056) <= 16069701;
srom_1(85057) <= 16282458;
srom_1(85058) <= 16458197;
srom_1(85059) <= 16596096;
srom_1(85060) <= 16695507;
srom_1(85061) <= 16755963;
srom_1(85062) <= 16777183;
srom_1(85063) <= 16759065;
srom_1(85064) <= 16701696;
srom_1(85065) <= 16605344;
srom_1(85066) <= 16470460;
srom_1(85067) <= 16297678;
srom_1(85068) <= 16087808;
srom_1(85069) <= 15841833;
srom_1(85070) <= 15560908;
srom_1(85071) <= 15246349;
srom_1(85072) <= 14899632;
srom_1(85073) <= 14522383;
srom_1(85074) <= 14116370;
srom_1(85075) <= 13683498;
srom_1(85076) <= 13225796;
srom_1(85077) <= 12745411;
srom_1(85078) <= 12244595;
srom_1(85079) <= 11725697;
srom_1(85080) <= 11191151;
srom_1(85081) <= 10643462;
srom_1(85082) <= 10085200;
srom_1(85083) <= 9518982;
srom_1(85084) <= 8947463;
srom_1(85085) <= 8373323;
srom_1(85086) <= 7799255;
srom_1(85087) <= 7227951;
srom_1(85088) <= 6662089;
srom_1(85089) <= 6104324;
srom_1(85090) <= 5557270;
srom_1(85091) <= 5023494;
srom_1(85092) <= 4505498;
srom_1(85093) <= 4005711;
srom_1(85094) <= 3526476;
srom_1(85095) <= 3070042;
srom_1(85096) <= 2638549;
srom_1(85097) <= 2234020;
srom_1(85098) <= 1858351;
srom_1(85099) <= 1513305;
srom_1(85100) <= 1200500;
srom_1(85101) <= 921402;
srom_1(85102) <= 677321;
srom_1(85103) <= 469401;
srom_1(85104) <= 298616;
srom_1(85105) <= 165768;
srom_1(85106) <= 71480;
srom_1(85107) <= 16194;
srom_1(85108) <= 168;
srom_1(85109) <= 23479;
srom_1(85110) <= 86017;
srom_1(85111) <= 187489;
srom_1(85112) <= 327419;
srom_1(85113) <= 505150;
srom_1(85114) <= 719850;
srom_1(85115) <= 970510;
srom_1(85116) <= 1255957;
srom_1(85117) <= 1574852;
srom_1(85118) <= 1925698;
srom_1(85119) <= 2306851;
srom_1(85120) <= 2716524;
srom_1(85121) <= 3152795;
srom_1(85122) <= 3613619;
srom_1(85123) <= 4096834;
srom_1(85124) <= 4600174;
srom_1(85125) <= 5121280;
srom_1(85126) <= 5657708;
srom_1(85127) <= 6206941;
srom_1(85128) <= 6766406;
srom_1(85129) <= 7333477;
srom_1(85130) <= 7905496;
srom_1(85131) <= 8479781;
srom_1(85132) <= 9053638;
srom_1(85133) <= 9624376;
srom_1(85134) <= 10189320;
srom_1(85135) <= 10745819;
srom_1(85136) <= 11291265;
srom_1(85137) <= 11823099;
srom_1(85138) <= 12338828;
srom_1(85139) <= 12836032;
srom_1(85140) <= 13312381;
srom_1(85141) <= 13765641;
srom_1(85142) <= 14193686;
srom_1(85143) <= 14594509;
srom_1(85144) <= 14966231;
srom_1(85145) <= 15307107;
srom_1(85146) <= 15615541;
srom_1(85147) <= 15890085;
srom_1(85148) <= 16129452;
srom_1(85149) <= 16332519;
srom_1(85150) <= 16498335;
srom_1(85151) <= 16626121;
srom_1(85152) <= 16715279;
srom_1(85153) <= 16765390;
srom_1(85154) <= 16776220;
srom_1(85155) <= 16747717;
srom_1(85156) <= 16680015;
srom_1(85157) <= 16573433;
srom_1(85158) <= 16428468;
srom_1(85159) <= 16245802;
srom_1(85160) <= 16026291;
srom_1(85161) <= 15770965;
srom_1(85162) <= 15481019;
srom_1(85163) <= 15157815;
srom_1(85164) <= 14802868;
srom_1(85165) <= 14417843;
srom_1(85166) <= 14004544;
srom_1(85167) <= 13564910;
srom_1(85168) <= 13101002;
srom_1(85169) <= 12614997;
srom_1(85170) <= 12109172;
srom_1(85171) <= 11585901;
srom_1(85172) <= 11047636;
srom_1(85173) <= 10496902;
srom_1(85174) <= 9936282;
srom_1(85175) <= 9368404;
srom_1(85176) <= 8795931;
srom_1(85177) <= 8221549;
srom_1(85178) <= 7647950;
srom_1(85179) <= 7077824;
srom_1(85180) <= 6513844;
srom_1(85181) <= 5958656;
srom_1(85182) <= 5414863;
srom_1(85183) <= 4885015;
srom_1(85184) <= 4371597;
srom_1(85185) <= 3877015;
srom_1(85186) <= 3403590;
srom_1(85187) <= 2953541;
srom_1(85188) <= 2528980;
srom_1(85189) <= 2131896;
srom_1(85190) <= 1764152;
srom_1(85191) <= 1427472;
srom_1(85192) <= 1123436;
srom_1(85193) <= 853468;
srom_1(85194) <= 618835;
srom_1(85195) <= 420637;
srom_1(85196) <= 259804;
srom_1(85197) <= 137090;
srom_1(85198) <= 53070;
srom_1(85199) <= 8138;
srom_1(85200) <= 2505;
srom_1(85201) <= 36197;
srom_1(85202) <= 109056;
srom_1(85203) <= 220742;
srom_1(85204) <= 370729;
srom_1(85205) <= 558314;
srom_1(85206) <= 782619;
srom_1(85207) <= 1042591;
srom_1(85208) <= 1337010;
srom_1(85209) <= 1664497;
srom_1(85210) <= 2023516;
srom_1(85211) <= 2412383;
srom_1(85212) <= 2829274;
srom_1(85213) <= 3272235;
srom_1(85214) <= 3739189;
srom_1(85215) <= 4227945;
srom_1(85216) <= 4736212;
srom_1(85217) <= 5261606;
srom_1(85218) <= 5801664;
srom_1(85219) <= 6353853;
srom_1(85220) <= 6915583;
srom_1(85221) <= 7484221;
srom_1(85222) <= 8057100;
srom_1(85223) <= 8631534;
srom_1(85224) <= 9204828;
srom_1(85225) <= 9774295;
srom_1(85226) <= 10337264;
srom_1(85227) <= 10891095;
srom_1(85228) <= 11433191;
srom_1(85229) <= 11961010;
srom_1(85230) <= 12472076;
srom_1(85231) <= 12963994;
srom_1(85232) <= 13434457;
srom_1(85233) <= 13881257;
srom_1(85234) <= 14302301;
srom_1(85235) <= 14695613;
srom_1(85236) <= 15059349;
srom_1(85237) <= 15391805;
srom_1(85238) <= 15691419;
srom_1(85239) <= 15956789;
srom_1(85240) <= 16186668;
srom_1(85241) <= 16379980;
srom_1(85242) <= 16535817;
srom_1(85243) <= 16653450;
srom_1(85244) <= 16732325;
srom_1(85245) <= 16772074;
srom_1(85246) <= 16772511;
srom_1(85247) <= 16733632;
srom_1(85248) <= 16655620;
srom_1(85249) <= 16538842;
srom_1(85250) <= 16383844;
srom_1(85251) <= 16191354;
srom_1(85252) <= 15962274;
srom_1(85253) <= 15697679;
srom_1(85254) <= 15398809;
srom_1(85255) <= 15067065;
srom_1(85256) <= 14704004;
srom_1(85257) <= 14311328;
srom_1(85258) <= 13890879;
srom_1(85259) <= 13444627;
srom_1(85260) <= 12974666;
srom_1(85261) <= 12483199;
srom_1(85262) <= 11972531;
srom_1(85263) <= 11445057;
srom_1(85264) <= 10903250;
srom_1(85265) <= 10349652;
srom_1(85266) <= 9786857;
srom_1(85267) <= 9217505;
srom_1(85268) <= 8644267;
srom_1(85269) <= 8069829;
srom_1(85270) <= 7496886;
srom_1(85271) <= 6928125;
srom_1(85272) <= 6366213;
srom_1(85273) <= 5813784;
srom_1(85274) <= 5273430;
srom_1(85275) <= 4747684;
srom_1(85276) <= 4239011;
srom_1(85277) <= 3749797;
srom_1(85278) <= 3282336;
srom_1(85279) <= 2838820;
srom_1(85280) <= 2421329;
srom_1(85281) <= 2031821;
srom_1(85282) <= 1672121;
srom_1(85283) <= 1343918;
srom_1(85284) <= 1048750;
srom_1(85285) <= 788000;
srom_1(85286) <= 562893;
srom_1(85287) <= 374483;
srom_1(85288) <= 223654;
srom_1(85289) <= 111113;
srom_1(85290) <= 37389;
srom_1(85291) <= 2826;
srom_1(85292) <= 7586;
srom_1(85293) <= 51649;
srom_1(85294) <= 134806;
srom_1(85295) <= 256668;
srom_1(85296) <= 416664;
srom_1(85297) <= 614042;
srom_1(85298) <= 847879;
srom_1(85299) <= 1117076;
srom_1(85300) <= 1420372;
srom_1(85301) <= 1756345;
srom_1(85302) <= 2123418;
srom_1(85303) <= 2519871;
srom_1(85304) <= 2943845;
srom_1(85305) <= 3393351;
srom_1(85306) <= 3866281;
srom_1(85307) <= 4360418;
srom_1(85308) <= 4873445;
srom_1(85309) <= 5402956;
srom_1(85310) <= 5946467;
srom_1(85311) <= 6501430;
srom_1(85312) <= 7065243;
srom_1(85313) <= 7635262;
srom_1(85314) <= 8208813;
srom_1(85315) <= 8783208;
srom_1(85316) <= 9355752;
srom_1(85317) <= 9923760;
srom_1(85318) <= 10484570;
srom_1(85319) <= 11035552;
srom_1(85320) <= 11574120;
srom_1(85321) <= 12097751;
srom_1(85322) <= 12603988;
srom_1(85323) <= 13090458;
srom_1(85324) <= 13554880;
srom_1(85325) <= 13995075;
srom_1(85326) <= 14408979;
srom_1(85327) <= 14794652;
srom_1(85328) <= 15150284;
srom_1(85329) <= 15474209;
srom_1(85330) <= 15764907;
srom_1(85331) <= 16021015;
srom_1(85332) <= 16241332;
srom_1(85333) <= 16424824;
srom_1(85334) <= 16570632;
srom_1(85335) <= 16678072;
srom_1(85336) <= 16746640;
srom_1(85337) <= 16776014;
srom_1(85338) <= 16766057;
srom_1(85339) <= 16716814;
srom_1(85340) <= 16628518;
srom_1(85341) <= 16501583;
srom_1(85342) <= 16336602;
srom_1(85343) <= 16134351;
srom_1(85344) <= 15895777;
srom_1(85345) <= 15622000;
srom_1(85346) <= 15314303;
srom_1(85347) <= 14974129;
srom_1(85348) <= 14603073;
srom_1(85349) <= 14202875;
srom_1(85350) <= 13775412;
srom_1(85351) <= 13322689;
srom_1(85352) <= 12846828;
srom_1(85353) <= 12350061;
srom_1(85354) <= 11834717;
srom_1(85355) <= 11303213;
srom_1(85356) <= 10758042;
srom_1(85357) <= 10201759;
srom_1(85358) <= 9636974;
srom_1(85359) <= 9066335;
srom_1(85360) <= 8492518;
srom_1(85361) <= 7918214;
srom_1(85362) <= 7346115;
srom_1(85363) <= 6778905;
srom_1(85364) <= 6219244;
srom_1(85365) <= 5669755;
srom_1(85366) <= 5133016;
srom_1(85367) <= 4611544;
srom_1(85368) <= 4107783;
srom_1(85369) <= 3624097;
srom_1(85370) <= 3162753;
srom_1(85371) <= 2725915;
srom_1(85372) <= 2315632;
srom_1(85373) <= 1933826;
srom_1(85374) <= 1582290;
srom_1(85375) <= 1262670;
srom_1(85376) <= 976467;
srom_1(85377) <= 725021;
srom_1(85378) <= 509513;
srom_1(85379) <= 330952;
srom_1(85380) <= 190177;
srom_1(85381) <= 87847;
srom_1(85382) <= 24442;
srom_1(85383) <= 259;
srom_1(85384) <= 15412;
srom_1(85385) <= 69830;
srom_1(85386) <= 163258;
srom_1(85387) <= 295257;
srom_1(85388) <= 465208;
srom_1(85389) <= 672315;
srom_1(85390) <= 915607;
srom_1(85391) <= 1193942;
srom_1(85392) <= 1506015;
srom_1(85393) <= 1850363;
srom_1(85394) <= 2225371;
srom_1(85395) <= 2629281;
srom_1(85396) <= 3060198;
srom_1(85397) <= 3516102;
srom_1(85398) <= 3994854;
srom_1(85399) <= 4494211;
srom_1(85400) <= 5011829;
srom_1(85401) <= 5545283;
srom_1(85402) <= 6092070;
srom_1(85403) <= 6649626;
srom_1(85404) <= 7215336;
srom_1(85405) <= 7786549;
srom_1(85406) <= 8360585;
srom_1(85407) <= 8934752;
srom_1(85408) <= 9506358;
srom_1(85409) <= 10072723;
srom_1(85410) <= 10631190;
srom_1(85411) <= 11179141;
srom_1(85412) <= 11714007;
srom_1(85413) <= 12233278;
srom_1(85414) <= 12734520;
srom_1(85415) <= 13215383;
srom_1(85416) <= 13673612;
srom_1(85417) <= 14107057;
srom_1(85418) <= 14513686;
srom_1(85419) <= 14891593;
srom_1(85420) <= 15239005;
srom_1(85421) <= 15554293;
srom_1(85422) <= 15835979;
srom_1(85423) <= 16082742;
srom_1(85424) <= 16293424;
srom_1(85425) <= 16467038;
srom_1(85426) <= 16602769;
srom_1(85427) <= 16699981;
srom_1(85428) <= 16758218;
srom_1(85429) <= 16777208;
srom_1(85430) <= 16756860;
srom_1(85431) <= 16697271;
srom_1(85432) <= 16598719;
srom_1(85433) <= 16461667;
srom_1(85434) <= 16286758;
srom_1(85435) <= 16074812;
srom_1(85436) <= 15826823;
srom_1(85437) <= 15543953;
srom_1(85438) <= 15227530;
srom_1(85439) <= 14879036;
srom_1(85440) <= 14500107;
srom_1(85441) <= 14092518;
srom_1(85442) <= 13658182;
srom_1(85443) <= 13199135;
srom_1(85444) <= 12717530;
srom_1(85445) <= 12215625;
srom_1(85446) <= 11695774;
srom_1(85447) <= 11160415;
srom_1(85448) <= 10612057;
srom_1(85449) <= 10053273;
srom_1(85450) <= 9486683;
srom_1(85451) <= 8914943;
srom_1(85452) <= 8340736;
srom_1(85453) <= 7766752;
srom_1(85454) <= 7195685;
srom_1(85455) <= 6630212;
srom_1(85456) <= 6072985;
srom_1(85457) <= 5526616;
srom_1(85458) <= 4993669;
srom_1(85459) <= 4476641;
srom_1(85460) <= 3977958;
srom_1(85461) <= 3499957;
srom_1(85462) <= 3044882;
srom_1(85463) <= 2614865;
srom_1(85464) <= 2211923;
srom_1(85465) <= 1837946;
srom_1(85466) <= 1494687;
srom_1(85467) <= 1183755;
srom_1(85468) <= 906610;
srom_1(85469) <= 664551;
srom_1(85470) <= 458712;
srom_1(85471) <= 290060;
srom_1(85472) <= 159384;
srom_1(85473) <= 67298;
srom_1(85474) <= 14233;
srom_1(85475) <= 438;
srom_1(85476) <= 25979;
srom_1(85477) <= 90735;
srom_1(85478) <= 194402;
srom_1(85479) <= 336495;
srom_1(85480) <= 516347;
srom_1(85481) <= 733115;
srom_1(85482) <= 985782;
srom_1(85483) <= 1273163;
srom_1(85484) <= 1593911;
srom_1(85485) <= 1946522;
srom_1(85486) <= 2329342;
srom_1(85487) <= 2740576;
srom_1(85488) <= 3178295;
srom_1(85489) <= 3640448;
srom_1(85490) <= 4124866;
srom_1(85491) <= 4629278;
srom_1(85492) <= 5151319;
srom_1(85493) <= 5688541;
srom_1(85494) <= 6238424;
srom_1(85495) <= 6798390;
srom_1(85496) <= 7365814;
srom_1(85497) <= 7938033;
srom_1(85498) <= 8512366;
srom_1(85499) <= 9086118;
srom_1(85500) <= 9656599;
srom_1(85501) <= 10221134;
srom_1(85502) <= 10777076;
srom_1(85503) <= 11321818;
srom_1(85504) <= 11852804;
srom_1(85505) <= 12367546;
srom_1(85506) <= 12863629;
srom_1(85507) <= 13338728;
srom_1(85508) <= 13790613;
srom_1(85509) <= 14217167;
srom_1(85510) <= 14616388;
srom_1(85511) <= 14986406;
srom_1(85512) <= 15325484;
srom_1(85513) <= 15632032;
srom_1(85514) <= 15904614;
srom_1(85515) <= 16141950;
srom_1(85516) <= 16342929;
srom_1(85517) <= 16506606;
srom_1(85518) <= 16632216;
srom_1(85519) <= 16719169;
srom_1(85520) <= 16767057;
srom_1(85521) <= 16775655;
srom_1(85522) <= 16744923;
srom_1(85523) <= 16675006;
srom_1(85524) <= 16566232;
srom_1(85525) <= 16419109;
srom_1(85526) <= 16234329;
srom_1(85527) <= 16012757;
srom_1(85528) <= 15755433;
srom_1(85529) <= 15463564;
srom_1(85530) <= 15138517;
srom_1(85531) <= 14781818;
srom_1(85532) <= 14395140;
srom_1(85533) <= 13980294;
srom_1(85534) <= 13539227;
srom_1(85535) <= 13074007;
srom_1(85536) <= 12586815;
srom_1(85537) <= 12079937;
srom_1(85538) <= 11555749;
srom_1(85539) <= 11016709;
srom_1(85540) <= 10465345;
srom_1(85541) <= 9904242;
srom_1(85542) <= 9336032;
srom_1(85543) <= 8763379;
srom_1(85544) <= 8188969;
srom_1(85545) <= 7615495;
srom_1(85546) <= 7045646;
srom_1(85547) <= 6482095;
srom_1(85548) <= 5927484;
srom_1(85549) <= 5384414;
srom_1(85550) <= 4855432;
srom_1(85551) <= 4343018;
srom_1(85552) <= 3849576;
srom_1(85553) <= 3377418;
srom_1(85554) <= 2928760;
srom_1(85555) <= 2505705;
srom_1(85556) <= 2110236;
srom_1(85557) <= 1744209;
srom_1(85558) <= 1409340;
srom_1(85559) <= 1107199;
srom_1(85560) <= 839204;
srom_1(85561) <= 606609;
srom_1(85562) <= 410508;
srom_1(85563) <= 251818;
srom_1(85564) <= 131285;
srom_1(85565) <= 49473;
srom_1(85566) <= 6766;
srom_1(85567) <= 3364;
srom_1(85568) <= 39284;
srom_1(85569) <= 114356;
srom_1(85570) <= 228230;
srom_1(85571) <= 380370;
srom_1(85572) <= 570063;
srom_1(85573) <= 796421;
srom_1(85574) <= 1058381;
srom_1(85575) <= 1354714;
srom_1(85576) <= 1684032;
srom_1(85577) <= 2044790;
srom_1(85578) <= 2435297;
srom_1(85579) <= 2853720;
srom_1(85580) <= 3298099;
srom_1(85581) <= 3766348;
srom_1(85582) <= 4256273;
srom_1(85583) <= 4765576;
srom_1(85584) <= 5291869;
srom_1(85585) <= 5832683;
srom_1(85586) <= 6385483;
srom_1(85587) <= 6947676;
srom_1(85588) <= 7516626;
srom_1(85589) <= 8089665;
srom_1(85590) <= 8664106;
srom_1(85591) <= 9237255;
srom_1(85592) <= 9806425;
srom_1(85593) <= 10368946;
srom_1(85594) <= 10922180;
srom_1(85595) <= 11463534;
srom_1(85596) <= 11990468;
srom_1(85597) <= 12500512;
srom_1(85598) <= 12991273;
srom_1(85599) <= 13460452;
srom_1(85600) <= 13905846;
srom_1(85601) <= 14325369;
srom_1(85602) <= 14717051;
srom_1(85603) <= 15079058;
srom_1(85604) <= 15409691;
srom_1(85605) <= 15707399;
srom_1(85606) <= 15970787;
srom_1(85607) <= 16198620;
srom_1(85608) <= 16389829;
srom_1(85609) <= 16543517;
srom_1(85610) <= 16658964;
srom_1(85611) <= 16735629;
srom_1(85612) <= 16773152;
srom_1(85613) <= 16771356;
srom_1(85614) <= 16730251;
srom_1(85615) <= 16650029;
srom_1(85616) <= 16531067;
srom_1(85617) <= 16373922;
srom_1(85618) <= 16179330;
srom_1(85619) <= 15948206;
srom_1(85620) <= 15681632;
srom_1(85621) <= 15380858;
srom_1(85622) <= 15047295;
srom_1(85623) <= 14682508;
srom_1(85624) <= 14288206;
srom_1(85625) <= 13866239;
srom_1(85626) <= 13418585;
srom_1(85627) <= 12947344;
srom_1(85628) <= 12454726;
srom_1(85629) <= 11943040;
srom_1(85630) <= 11414686;
srom_1(85631) <= 10872142;
srom_1(85632) <= 10317952;
srom_1(85633) <= 9754715;
srom_1(85634) <= 9185071;
srom_1(85635) <= 8611692;
srom_1(85636) <= 8037267;
srom_1(85637) <= 7464490;
srom_1(85638) <= 6896046;
srom_1(85639) <= 6334602;
srom_1(85640) <= 5782789;
srom_1(85641) <= 5243196;
srom_1(85642) <= 4718353;
srom_1(85643) <= 4210721;
srom_1(85644) <= 3722680;
srom_1(85645) <= 3256520;
srom_1(85646) <= 2814425;
srom_1(85647) <= 2398470;
srom_1(85648) <= 2010605;
srom_1(85649) <= 1652648;
srom_1(85650) <= 1326279;
srom_1(85651) <= 1033027;
srom_1(85652) <= 774268;
srom_1(85653) <= 551216;
srom_1(85654) <= 364915;
srom_1(85655) <= 216241;
srom_1(85656) <= 105889;
srom_1(85657) <= 34378;
srom_1(85658) <= 2043;
srom_1(85659) <= 9035;
srom_1(85660) <= 55322;
srom_1(85661) <= 140687;
srom_1(85662) <= 264729;
srom_1(85663) <= 426866;
srom_1(85664) <= 626339;
srom_1(85665) <= 862212;
srom_1(85666) <= 1133379;
srom_1(85667) <= 1438568;
srom_1(85668) <= 1776348;
srom_1(85669) <= 2145135;
srom_1(85670) <= 2543200;
srom_1(85671) <= 2968676;
srom_1(85672) <= 3419568;
srom_1(85673) <= 3893762;
srom_1(85674) <= 4389034;
srom_1(85675) <= 4903060;
srom_1(85676) <= 5433432;
srom_1(85677) <= 5977662;
srom_1(85678) <= 6533197;
srom_1(85679) <= 7097433;
srom_1(85680) <= 7667724;
srom_1(85681) <= 8241395;
srom_1(85682) <= 8815756;
srom_1(85683) <= 9388115;
srom_1(85684) <= 9955786;
srom_1(85685) <= 10516109;
srom_1(85686) <= 11066454;
srom_1(85687) <= 11604243;
srom_1(85688) <= 12126952;
srom_1(85689) <= 12632131;
srom_1(85690) <= 13117411;
srom_1(85691) <= 13580515;
srom_1(85692) <= 14019273;
srom_1(85693) <= 14431627;
srom_1(85694) <= 14815643;
srom_1(85695) <= 15169520;
srom_1(85696) <= 15491599;
srom_1(85697) <= 15780370;
srom_1(85698) <= 16034479;
srom_1(85699) <= 16252733;
srom_1(85700) <= 16434110;
srom_1(85701) <= 16577758;
srom_1(85702) <= 16683005;
srom_1(85703) <= 16749357;
srom_1(85704) <= 16776502;
srom_1(85705) <= 16764313;
srom_1(85706) <= 16712848;
srom_1(85707) <= 16622348;
srom_1(85708) <= 16493236;
srom_1(85709) <= 16326120;
srom_1(85710) <= 16121781;
srom_1(85711) <= 15881180;
srom_1(85712) <= 15605442;
srom_1(85713) <= 15295863;
srom_1(85714) <= 14953893;
srom_1(85715) <= 14581137;
srom_1(85716) <= 14179341;
srom_1(85717) <= 13750391;
srom_1(85718) <= 13296297;
srom_1(85719) <= 12819190;
srom_1(85720) <= 12321306;
srom_1(85721) <= 11804980;
srom_1(85722) <= 11272633;
srom_1(85723) <= 10726763;
srom_1(85724) <= 10169928;
srom_1(85725) <= 9604740;
srom_1(85726) <= 9033849;
srom_1(85727) <= 8459932;
srom_1(85728) <= 7885681;
srom_1(85729) <= 7313788;
srom_1(85730) <= 6746935;
srom_1(85731) <= 6187781;
srom_1(85732) <= 5638947;
srom_1(85733) <= 5103007;
srom_1(85734) <= 4582475;
srom_1(85735) <= 4079791;
srom_1(85736) <= 3597312;
srom_1(85737) <= 3137301;
srom_1(85738) <= 2701916;
srom_1(85739) <= 2293197;
srom_1(85740) <= 1913062;
srom_1(85741) <= 1563293;
srom_1(85742) <= 1245530;
srom_1(85743) <= 961263;
srom_1(85744) <= 711826;
srom_1(85745) <= 498388;
srom_1(85746) <= 321950;
srom_1(85747) <= 183339;
srom_1(85748) <= 83205;
srom_1(85749) <= 22019;
srom_1(85750) <= 66;
srom_1(85751) <= 17450;
srom_1(85752) <= 74089;
srom_1(85753) <= 169718;
srom_1(85754) <= 303888;
srom_1(85755) <= 475970;
srom_1(85756) <= 685157;
srom_1(85757) <= 930468;
srom_1(85758) <= 1210753;
srom_1(85759) <= 1524697;
srom_1(85760) <= 1870829;
srom_1(85761) <= 2247524;
srom_1(85762) <= 2653018;
srom_1(85763) <= 3085407;
srom_1(85764) <= 3542665;
srom_1(85765) <= 4022647;
srom_1(85766) <= 4523103;
srom_1(85767) <= 5041686;
srom_1(85768) <= 5575963;
srom_1(85769) <= 6123430;
srom_1(85770) <= 6681519;
srom_1(85771) <= 7247613;
srom_1(85772) <= 7819057;
srom_1(85773) <= 8393173;
srom_1(85774) <= 8967267;
srom_1(85775) <= 9538647;
srom_1(85776) <= 10104635;
srom_1(85777) <= 10662575;
srom_1(85778) <= 11209852;
srom_1(85779) <= 11743899;
srom_1(85780) <= 12262213;
srom_1(85781) <= 12762361;
srom_1(85782) <= 13241999;
srom_1(85783) <= 13698879;
srom_1(85784) <= 14130856;
srom_1(85785) <= 14535906;
srom_1(85786) <= 14912130;
srom_1(85787) <= 15257762;
srom_1(85788) <= 15571182;
srom_1(85789) <= 15850921;
srom_1(85790) <= 16095667;
srom_1(85791) <= 16304271;
srom_1(85792) <= 16475756;
srom_1(85793) <= 16609318;
srom_1(85794) <= 16704330;
srom_1(85795) <= 16760347;
srom_1(85796) <= 16777106;
srom_1(85797) <= 16754528;
srom_1(85798) <= 16692720;
srom_1(85799) <= 16591970;
srom_1(85800) <= 16452753;
srom_1(85801) <= 16275719;
srom_1(85802) <= 16061701;
srom_1(85803) <= 15811700;
srom_1(85804) <= 15526891;
srom_1(85805) <= 15208607;
srom_1(85806) <= 14858342;
srom_1(85807) <= 14477738;
srom_1(85808) <= 14068580;
srom_1(85809) <= 13632787;
srom_1(85810) <= 13172402;
srom_1(85811) <= 12689584;
srom_1(85812) <= 12186598;
srom_1(85813) <= 11665801;
srom_1(85814) <= 11129636;
srom_1(85815) <= 10580618;
srom_1(85816) <= 10021321;
srom_1(85817) <= 9454367;
srom_1(85818) <= 8882416;
srom_1(85819) <= 8308149;
srom_1(85820) <= 7734259;
srom_1(85821) <= 7163438;
srom_1(85822) <= 6598362;
srom_1(85823) <= 6041681;
srom_1(85824) <= 5496005;
srom_1(85825) <= 4963894;
srom_1(85826) <= 4447843;
srom_1(85827) <= 3950271;
srom_1(85828) <= 3473512;
srom_1(85829) <= 3019802;
srom_1(85830) <= 2591268;
srom_1(85831) <= 2189920;
srom_1(85832) <= 1817639;
srom_1(85833) <= 1476172;
srom_1(85834) <= 1167119;
srom_1(85835) <= 891931;
srom_1(85836) <= 651897;
srom_1(85837) <= 448143;
srom_1(85838) <= 281625;
srom_1(85839) <= 153123;
srom_1(85840) <= 63241;
srom_1(85841) <= 12398;
srom_1(85842) <= 835;
srom_1(85843) <= 28605;
srom_1(85844) <= 95578;
srom_1(85845) <= 201439;
srom_1(85846) <= 345693;
srom_1(85847) <= 527663;
srom_1(85848) <= 746496;
srom_1(85849) <= 1001165;
srom_1(85850) <= 1290476;
srom_1(85851) <= 1613073;
srom_1(85852) <= 1967443;
srom_1(85853) <= 2351924;
srom_1(85854) <= 2764713;
srom_1(85855) <= 3203874;
srom_1(85856) <= 3667348;
srom_1(85857) <= 4152962;
srom_1(85858) <= 4658439;
srom_1(85859) <= 5181407;
srom_1(85860) <= 5719415;
srom_1(85861) <= 6269939;
srom_1(85862) <= 6830399;
srom_1(85863) <= 7398166;
srom_1(85864) <= 7970577;
srom_1(85865) <= 8544949;
srom_1(85866) <= 9118588;
srom_1(85867) <= 9688803;
srom_1(85868) <= 10252921;
srom_1(85869) <= 10808297;
srom_1(85870) <= 11352326;
srom_1(85871) <= 11882457;
srom_1(85872) <= 12396205;
srom_1(85873) <= 12891159;
srom_1(85874) <= 13364999;
srom_1(85875) <= 13815504;
srom_1(85876) <= 14240559;
srom_1(85877) <= 14638173;
srom_1(85878) <= 15006481;
srom_1(85879) <= 15343755;
srom_1(85880) <= 15648414;
srom_1(85881) <= 15919029;
srom_1(85882) <= 16154332;
srom_1(85883) <= 16353218;
srom_1(85884) <= 16514756;
srom_1(85885) <= 16638187;
srom_1(85886) <= 16722933;
srom_1(85887) <= 16768596;
srom_1(85888) <= 16774963;
srom_1(85889) <= 16742004;
srom_1(85890) <= 16669872;
srom_1(85891) <= 16558907;
srom_1(85892) <= 16409629;
srom_1(85893) <= 16222737;
srom_1(85894) <= 15999108;
srom_1(85895) <= 15739791;
srom_1(85896) <= 15446002;
srom_1(85897) <= 15119118;
srom_1(85898) <= 14760672;
srom_1(85899) <= 14372346;
srom_1(85900) <= 13955960;
srom_1(85901) <= 13513466;
srom_1(85902) <= 13046941;
srom_1(85903) <= 12558571;
srom_1(85904) <= 12050646;
srom_1(85905) <= 11525549;
srom_1(85906) <= 10985742;
srom_1(85907) <= 10433756;
srom_1(85908) <= 9872179;
srom_1(85909) <= 9303645;
srom_1(85910) <= 8730821;
srom_1(85911) <= 8156392;
srom_1(85912) <= 7583051;
srom_1(85913) <= 7013489;
srom_1(85914) <= 6450374;
srom_1(85915) <= 5896349;
srom_1(85916) <= 5354011;
srom_1(85917) <= 4825903;
srom_1(85918) <= 4314501;
srom_1(85919) <= 3822205;
srom_1(85920) <= 3351322;
srom_1(85921) <= 2904061;
srom_1(85922) <= 2482518;
srom_1(85923) <= 2088671;
srom_1(85924) <= 1724367;
srom_1(85925) <= 1391314;
srom_1(85926) <= 1091073;
srom_1(85927) <= 825053;
srom_1(85928) <= 594501;
srom_1(85929) <= 400499;
srom_1(85930) <= 243955;
srom_1(85931) <= 125604;
srom_1(85932) <= 46002;
srom_1(85933) <= 5520;
srom_1(85934) <= 4350;
srom_1(85935) <= 42497;
srom_1(85936) <= 119781;
srom_1(85937) <= 235841;
srom_1(85938) <= 390132;
srom_1(85939) <= 581931;
srom_1(85940) <= 810337;
srom_1(85941) <= 1074281;
srom_1(85942) <= 1372524;
srom_1(85943) <= 1703668;
srom_1(85944) <= 2066160;
srom_1(85945) <= 2458300;
srom_1(85946) <= 2878249;
srom_1(85947) <= 3324039;
srom_1(85948) <= 3793577;
srom_1(85949) <= 4284664;
srom_1(85950) <= 4794995;
srom_1(85951) <= 5322178;
srom_1(85952) <= 5863740;
srom_1(85953) <= 6417143;
srom_1(85954) <= 6979790;
srom_1(85955) <= 7549044;
srom_1(85956) <= 8122235;
srom_1(85957) <= 8696674;
srom_1(85958) <= 9269669;
srom_1(85959) <= 9838533;
srom_1(85960) <= 10400597;
srom_1(85961) <= 10953227;
srom_1(85962) <= 11493830;
srom_1(85963) <= 12019872;
srom_1(85964) <= 12528885;
srom_1(85965) <= 13018483;
srom_1(85966) <= 13486370;
srom_1(85967) <= 13930352;
srom_1(85968) <= 14348347;
srom_1(85969) <= 14738394;
srom_1(85970) <= 15098666;
srom_1(85971) <= 15427471;
srom_1(85972) <= 15723269;
srom_1(85973) <= 15984672;
srom_1(85974) <= 16210454;
srom_1(85975) <= 16399557;
srom_1(85976) <= 16551094;
srom_1(85977) <= 16664354;
srom_1(85978) <= 16738807;
srom_1(85979) <= 16774102;
srom_1(85980) <= 16770075;
srom_1(85981) <= 16726745;
srom_1(85982) <= 16644314;
srom_1(85983) <= 16523169;
srom_1(85984) <= 16363879;
srom_1(85985) <= 16167189;
srom_1(85986) <= 15934023;
srom_1(85987) <= 15665475;
srom_1(85988) <= 15362802;
srom_1(85989) <= 15027425;
srom_1(85990) <= 14660916;
srom_1(85991) <= 14264995;
srom_1(85992) <= 13841517;
srom_1(85993) <= 13392468;
srom_1(85994) <= 12919954;
srom_1(85995) <= 12426192;
srom_1(85996) <= 11913496;
srom_1(85997) <= 11384270;
srom_1(85998) <= 10840997;
srom_1(85999) <= 10286223;
srom_1(86000) <= 9722551;
srom_1(86001) <= 9152624;
srom_1(86002) <= 8579114;
srom_1(86003) <= 8004711;
srom_1(86004) <= 7432108;
srom_1(86005) <= 6863990;
srom_1(86006) <= 6303021;
srom_1(86007) <= 5751833;
srom_1(86008) <= 5213010;
srom_1(86009) <= 4689077;
srom_1(86010) <= 4182494;
srom_1(86011) <= 3695634;
srom_1(86012) <= 3230781;
srom_1(86013) <= 2790115;
srom_1(86014) <= 2375702;
srom_1(86015) <= 1989486;
srom_1(86016) <= 1633277;
srom_1(86017) <= 1308747;
srom_1(86018) <= 1017416;
srom_1(86019) <= 760651;
srom_1(86020) <= 539657;
srom_1(86021) <= 355469;
srom_1(86022) <= 208951;
srom_1(86023) <= 100790;
srom_1(86024) <= 31494;
srom_1(86025) <= 1387;
srom_1(86026) <= 10611;
srom_1(86027) <= 59122;
srom_1(86028) <= 146692;
srom_1(86029) <= 272912;
srom_1(86030) <= 437190;
srom_1(86031) <= 638754;
srom_1(86032) <= 876660;
srom_1(86033) <= 1149791;
srom_1(86034) <= 1456869;
srom_1(86035) <= 1796451;
srom_1(86036) <= 2166947;
srom_1(86037) <= 2566618;
srom_1(86038) <= 2993590;
srom_1(86039) <= 3445861;
srom_1(86040) <= 3921311;
srom_1(86041) <= 4417709;
srom_1(86042) <= 4932728;
srom_1(86043) <= 5463953;
srom_1(86044) <= 6008893;
srom_1(86045) <= 6564992;
srom_1(86046) <= 7129642;
srom_1(86047) <= 7700196;
srom_1(86048) <= 8273979;
srom_1(86049) <= 8848299;
srom_1(86050) <= 9420463;
srom_1(86051) <= 9987788;
srom_1(86052) <= 10547615;
srom_1(86053) <= 11097317;
srom_1(86054) <= 11634317;
srom_1(86055) <= 12156097;
srom_1(86056) <= 12660210;
srom_1(86057) <= 13144291;
srom_1(86058) <= 13606072;
srom_1(86059) <= 14043386;
srom_1(86060) <= 14454183;
srom_1(86061) <= 14836536;
srom_1(86062) <= 15188653;
srom_1(86063) <= 15508882;
srom_1(86064) <= 15795722;
srom_1(86065) <= 16047827;
srom_1(86066) <= 16264016;
srom_1(86067) <= 16443274;
srom_1(86068) <= 16584760;
srom_1(86069) <= 16687813;
srom_1(86070) <= 16751947;
srom_1(86071) <= 16776863;
srom_1(86072) <= 16762443;
srom_1(86073) <= 16708756;
srom_1(86074) <= 16616053;
srom_1(86075) <= 16484768;
srom_1(86076) <= 16315518;
srom_1(86077) <= 16109095;
srom_1(86078) <= 15866469;
srom_1(86079) <= 15588776;
srom_1(86080) <= 15277319;
srom_1(86081) <= 14933559;
srom_1(86082) <= 14559107;
srom_1(86083) <= 14155720;
srom_1(86084) <= 13725288;
srom_1(86085) <= 13269831;
srom_1(86086) <= 12791485;
srom_1(86087) <= 12292491;
srom_1(86088) <= 11775191;
srom_1(86089) <= 11242010;
srom_1(86090) <= 10695449;
srom_1(86091) <= 10138070;
srom_1(86092) <= 9572487;
srom_1(86093) <= 9001353;
srom_1(86094) <= 8427345;
srom_1(86095) <= 7853156;
srom_1(86096) <= 7281477;
srom_1(86097) <= 6714990;
srom_1(86098) <= 6156351;
srom_1(86099) <= 5608181;
srom_1(86100) <= 5073048;
srom_1(86101) <= 4553463;
srom_1(86102) <= 4051863;
srom_1(86103) <= 3570599;
srom_1(86104) <= 3111928;
srom_1(86105) <= 2678002;
srom_1(86106) <= 2270854;
srom_1(86107) <= 1892395;
srom_1(86108) <= 1544399;
srom_1(86109) <= 1228497;
srom_1(86110) <= 946172;
srom_1(86111) <= 698747;
srom_1(86112) <= 487382;
srom_1(86113) <= 313069;
srom_1(86114) <= 176625;
srom_1(86115) <= 78690;
srom_1(86116) <= 19722;
srom_1(86117) <= 0;
srom_1(86118) <= 19614;
srom_1(86119) <= 78473;
srom_1(86120) <= 176302;
srom_1(86121) <= 312640;
srom_1(86122) <= 486850;
srom_1(86123) <= 698114;
srom_1(86124) <= 945441;
srom_1(86125) <= 1227672;
srom_1(86126) <= 1543483;
srom_1(86127) <= 1891393;
srom_1(86128) <= 2269770;
srom_1(86129) <= 2676841;
srom_1(86130) <= 3110697;
srom_1(86131) <= 3569302;
srom_1(86132) <= 4050507;
srom_1(86133) <= 4552054;
srom_1(86134) <= 5071593;
srom_1(86135) <= 5606686;
srom_1(86136) <= 6154824;
srom_1(86137) <= 6713437;
srom_1(86138) <= 7279906;
srom_1(86139) <= 7851574;
srom_1(86140) <= 8425760;
srom_1(86141) <= 8999772;
srom_1(86142) <= 9570919;
srom_1(86143) <= 10136520;
srom_1(86144) <= 10693926;
srom_1(86145) <= 11240520;
srom_1(86146) <= 11773742;
srom_1(86147) <= 12291089;
srom_1(86148) <= 12790136;
srom_1(86149) <= 13268542;
srom_1(86150) <= 13724066;
srom_1(86151) <= 14154569;
srom_1(86152) <= 14558033;
srom_1(86153) <= 14932568;
srom_1(86154) <= 15276415;
srom_1(86155) <= 15587963;
srom_1(86156) <= 15865750;
srom_1(86157) <= 16108475;
srom_1(86158) <= 16314999;
srom_1(86159) <= 16484353;
srom_1(86160) <= 16615743;
srom_1(86161) <= 16708554;
srom_1(86162) <= 16762349;
srom_1(86163) <= 16776877;
srom_1(86164) <= 16752070;
srom_1(86165) <= 16688043;
srom_1(86166) <= 16585098;
srom_1(86167) <= 16443716;
srom_1(86168) <= 16264561;
srom_1(86169) <= 16048473;
srom_1(86170) <= 15796466;
srom_1(86171) <= 15509720;
srom_1(86172) <= 15189581;
srom_1(86173) <= 14837550;
srom_1(86174) <= 14455278;
srom_1(86175) <= 14044556;
srom_1(86176) <= 13607313;
srom_1(86177) <= 13145596;
srom_1(86178) <= 12661573;
srom_1(86179) <= 12157513;
srom_1(86180) <= 11635778;
srom_1(86181) <= 11098817;
srom_1(86182) <= 10549146;
srom_1(86183) <= 9989344;
srom_1(86184) <= 9422035;
srom_1(86185) <= 8849881;
srom_1(86186) <= 8275563;
srom_1(86187) <= 7701776;
srom_1(86188) <= 7131209;
srom_1(86189) <= 6566538;
srom_1(86190) <= 6010412;
srom_1(86191) <= 5465438;
srom_1(86192) <= 4934172;
srom_1(86193) <= 4419105;
srom_1(86194) <= 3922652;
srom_1(86195) <= 3447142;
srom_1(86196) <= 2994803;
srom_1(86197) <= 2567759;
srom_1(86198) <= 2168010;
srom_1(86199) <= 1797431;
srom_1(86200) <= 1457761;
srom_1(86201) <= 1150592;
srom_1(86202) <= 877365;
srom_1(86203) <= 639360;
srom_1(86204) <= 437695;
srom_1(86205) <= 273313;
srom_1(86206) <= 146988;
srom_1(86207) <= 59310;
srom_1(86208) <= 10691;
srom_1(86209) <= 1358;
srom_1(86210) <= 31357;
srom_1(86211) <= 100546;
srom_1(86212) <= 208600;
srom_1(86213) <= 355013;
srom_1(86214) <= 539098;
srom_1(86215) <= 759992;
srom_1(86216) <= 1016660;
srom_1(86217) <= 1307897;
srom_1(86218) <= 1632338;
srom_1(86219) <= 1988461;
srom_1(86220) <= 2374597;
srom_1(86221) <= 2788935;
srom_1(86222) <= 3229531;
srom_1(86223) <= 3694320;
srom_1(86224) <= 4181123;
srom_1(86225) <= 4687655;
srom_1(86226) <= 5211543;
srom_1(86227) <= 5750329;
srom_1(86228) <= 6301487;
srom_1(86229) <= 6862432;
srom_1(86230) <= 7430533;
srom_1(86231) <= 8003128;
srom_1(86232) <= 8577530;
srom_1(86233) <= 9151046;
srom_1(86234) <= 9720987;
srom_1(86235) <= 10284680;
srom_1(86236) <= 10839481;
srom_1(86237) <= 11382790;
srom_1(86238) <= 11912058;
srom_1(86239) <= 12424803;
srom_1(86240) <= 12918621;
srom_1(86241) <= 13391196;
srom_1(86242) <= 13840312;
srom_1(86243) <= 14263864;
srom_1(86244) <= 14659864;
srom_1(86245) <= 15026456;
srom_1(86246) <= 15361921;
srom_1(86247) <= 15664686;
srom_1(86248) <= 15933331;
srom_1(86249) <= 16166596;
srom_1(86250) <= 16363387;
srom_1(86251) <= 16522782;
srom_1(86252) <= 16644033;
srom_1(86253) <= 16726571;
srom_1(86254) <= 16770010;
srom_1(86255) <= 16774145;
srom_1(86256) <= 16738958;
srom_1(86257) <= 16664613;
srom_1(86258) <= 16551459;
srom_1(86259) <= 16400027;
srom_1(86260) <= 16211026;
srom_1(86261) <= 15985344;
srom_1(86262) <= 15724037;
srom_1(86263) <= 15428333;
srom_1(86264) <= 15099616;
srom_1(86265) <= 14739430;
srom_1(86266) <= 14349462;
srom_1(86267) <= 13931542;
srom_1(86268) <= 13487628;
srom_1(86269) <= 13019804;
srom_1(86270) <= 12530263;
srom_1(86271) <= 12021300;
srom_1(86272) <= 11495302;
srom_1(86273) <= 10954736;
srom_1(86274) <= 10402136;
srom_1(86275) <= 9840094;
srom_1(86276) <= 9271245;
srom_1(86277) <= 8698258;
srom_1(86278) <= 8123818;
srom_1(86279) <= 7550620;
srom_1(86280) <= 6981352;
srom_1(86281) <= 6418683;
srom_1(86282) <= 5865252;
srom_1(86283) <= 5323653;
srom_1(86284) <= 4796427;
srom_1(86285) <= 4286046;
srom_1(86286) <= 3794903;
srom_1(86287) <= 3325302;
srom_1(86288) <= 2879444;
srom_1(86289) <= 2459421;
srom_1(86290) <= 2067202;
srom_1(86291) <= 1704625;
srom_1(86292) <= 1373393;
srom_1(86293) <= 1075057;
srom_1(86294) <= 811017;
srom_1(86295) <= 582511;
srom_1(86296) <= 390610;
srom_1(86297) <= 236214;
srom_1(86298) <= 120048;
srom_1(86299) <= 42657;
srom_1(86300) <= 4402;
srom_1(86301) <= 5463;
srom_1(86302) <= 45836;
srom_1(86303) <= 125331;
srom_1(86304) <= 243576;
srom_1(86305) <= 400015;
srom_1(86306) <= 593915;
srom_1(86307) <= 824368;
srom_1(86308) <= 1090292;
srom_1(86309) <= 1390440;
srom_1(86310) <= 1723405;
srom_1(86311) <= 2087625;
srom_1(86312) <= 2481393;
srom_1(86313) <= 2902862;
srom_1(86314) <= 3350055;
srom_1(86315) <= 3820876;
srom_1(86316) <= 4313116;
srom_1(86317) <= 4824468;
srom_1(86318) <= 5352534;
srom_1(86319) <= 5894836;
srom_1(86320) <= 6448833;
srom_1(86321) <= 7011926;
srom_1(86322) <= 7581474;
srom_1(86323) <= 8154808;
srom_1(86324) <= 8729238;
srom_1(86325) <= 9302070;
srom_1(86326) <= 9870619;
srom_1(86327) <= 10432219;
srom_1(86328) <= 10984235;
srom_1(86329) <= 11524079;
srom_1(86330) <= 12049220;
srom_1(86331) <= 12557196;
srom_1(86332) <= 13045623;
srom_1(86333) <= 13512212;
srom_1(86334) <= 13954774;
srom_1(86335) <= 14371235;
srom_1(86336) <= 14759641;
srom_1(86337) <= 15118172;
srom_1(86338) <= 15445145;
srom_1(86339) <= 15739027;
srom_1(86340) <= 15998441;
srom_1(86341) <= 16222170;
srom_1(86342) <= 16409165;
srom_1(86343) <= 16558548;
srom_1(86344) <= 16669620;
srom_1(86345) <= 16741859;
srom_1(86346) <= 16774927;
srom_1(86347) <= 16768668;
srom_1(86348) <= 16723113;
srom_1(86349) <= 16638474;
srom_1(86350) <= 16515149;
srom_1(86351) <= 16353715;
srom_1(86352) <= 16154931;
srom_1(86353) <= 15919727;
srom_1(86354) <= 15649208;
srom_1(86355) <= 15344641;
srom_1(86356) <= 15007454;
srom_1(86357) <= 14639230;
srom_1(86358) <= 14241695;
srom_1(86359) <= 13816712;
srom_1(86360) <= 13366275;
srom_1(86361) <= 12892496;
srom_1(86362) <= 12397597;
srom_1(86363) <= 11883898;
srom_1(86364) <= 11353809;
srom_1(86365) <= 10809814;
srom_1(86366) <= 10254466;
srom_1(86367) <= 9690368;
srom_1(86368) <= 9120166;
srom_1(86369) <= 8546533;
srom_1(86370) <= 7972160;
srom_1(86371) <= 7399740;
srom_1(86372) <= 6831956;
srom_1(86373) <= 6271473;
srom_1(86374) <= 5720917;
srom_1(86375) <= 5182871;
srom_1(86376) <= 4659858;
srom_1(86377) <= 4154330;
srom_1(86378) <= 3668658;
srom_1(86379) <= 3205120;
srom_1(86380) <= 2765889;
srom_1(86381) <= 2353024;
srom_1(86382) <= 1968463;
srom_1(86383) <= 1614008;
srom_1(86384) <= 1291321;
srom_1(86385) <= 1001916;
srom_1(86386) <= 747150;
srom_1(86387) <= 528217;
srom_1(86388) <= 346144;
srom_1(86389) <= 201785;
srom_1(86390) <= 95816;
srom_1(86391) <= 28736;
srom_1(86392) <= 858;
srom_1(86393) <= 12313;
srom_1(86394) <= 63047;
srom_1(86395) <= 152822;
srom_1(86396) <= 281218;
srom_1(86397) <= 447633;
srom_1(86398) <= 651285;
srom_1(86399) <= 891220;
srom_1(86400) <= 1166313;
srom_1(86401) <= 1475274;
srom_1(86402) <= 1816654;
srom_1(86403) <= 2188852;
srom_1(86404) <= 2590123;
srom_1(86405) <= 3018585;
srom_1(86406) <= 3472228;
srom_1(86407) <= 3948927;
srom_1(86408) <= 4446444;
srom_1(86409) <= 4962448;
srom_1(86410) <= 5494518;
srom_1(86411) <= 6040160;
srom_1(86412) <= 6596814;
srom_1(86413) <= 7161870;
srom_1(86414) <= 7732679;
srom_1(86415) <= 8306564;
srom_1(86416) <= 8880834;
srom_1(86417) <= 9452795;
srom_1(86418) <= 10019767;
srom_1(86419) <= 10579089;
srom_1(86420) <= 11128139;
srom_1(86421) <= 11664342;
srom_1(86422) <= 12185185;
srom_1(86423) <= 12688224;
srom_1(86424) <= 13171100;
srom_1(86425) <= 13631550;
srom_1(86426) <= 14067414;
srom_1(86427) <= 14476648;
srom_1(86428) <= 14857333;
srom_1(86429) <= 15207684;
srom_1(86430) <= 15526058;
srom_1(86431) <= 15810962;
srom_1(86432) <= 16061060;
srom_1(86433) <= 16275180;
srom_1(86434) <= 16452316;
srom_1(86435) <= 16591639;
srom_1(86436) <= 16692495;
srom_1(86437) <= 16754411;
srom_1(86438) <= 16777098;
srom_1(86439) <= 16760447;
srom_1(86440) <= 16704539;
srom_1(86441) <= 16609633;
srom_1(86442) <= 16476177;
srom_1(86443) <= 16304796;
srom_1(86444) <= 16096292;
srom_1(86445) <= 15851645;
srom_1(86446) <= 15572001;
srom_1(86447) <= 15258671;
srom_1(86448) <= 14913126;
srom_1(86449) <= 14536984;
srom_1(86450) <= 14132011;
srom_1(86451) <= 13700105;
srom_1(86452) <= 13243292;
srom_1(86453) <= 12763713;
srom_1(86454) <= 12263618;
srom_1(86455) <= 11745352;
srom_1(86456) <= 11211344;
srom_1(86457) <= 10664100;
srom_1(86458) <= 10106186;
srom_1(86459) <= 9540217;
srom_1(86460) <= 8968848;
srom_1(86461) <= 8394757;
srom_1(86462) <= 7820638;
srom_1(86463) <= 7249183;
srom_1(86464) <= 6683070;
srom_1(86465) <= 6124955;
srom_1(86466) <= 5577456;
srom_1(86467) <= 5043139;
srom_1(86468) <= 4524510;
srom_1(86469) <= 4024001;
srom_1(86470) <= 3543959;
srom_1(86471) <= 3086635;
srom_1(86472) <= 2654174;
srom_1(86473) <= 2248604;
srom_1(86474) <= 1871826;
srom_1(86475) <= 1525608;
srom_1(86476) <= 1211573;
srom_1(86477) <= 931193;
srom_1(86478) <= 685784;
srom_1(86479) <= 476496;
srom_1(86480) <= 304310;
srom_1(86481) <= 170035;
srom_1(86482) <= 74299;
srom_1(86483) <= 17552;
srom_1(86484) <= 60;
srom_1(86485) <= 21904;
srom_1(86486) <= 82983;
srom_1(86487) <= 183010;
srom_1(86488) <= 321515;
srom_1(86489) <= 497850;
srom_1(86490) <= 711188;
srom_1(86491) <= 960527;
srom_1(86492) <= 1244699;
srom_1(86493) <= 1562372;
srom_1(86494) <= 1912055;
srom_1(86495) <= 2292109;
srom_1(86496) <= 2700751;
srom_1(86497) <= 3136066;
srom_1(86498) <= 3596011;
srom_1(86499) <= 4078431;
srom_1(86500) <= 4581063;
srom_1(86501) <= 5101549;
srom_1(86502) <= 5637450;
srom_1(86503) <= 6186252;
srom_1(86504) <= 6745381;
srom_1(86505) <= 7312217;
srom_1(86506) <= 7884099;
srom_1(86507) <= 8458348;
srom_1(86508) <= 9032269;
srom_1(86509) <= 9603172;
srom_1(86510) <= 10168380;
srom_1(86511) <= 10725241;
srom_1(86512) <= 11271145;
srom_1(86513) <= 11803533;
srom_1(86514) <= 12319906;
srom_1(86515) <= 12817844;
srom_1(86516) <= 13295012;
srom_1(86517) <= 13749172;
srom_1(86518) <= 14178194;
srom_1(86519) <= 14580068;
srom_1(86520) <= 14952907;
srom_1(86521) <= 15294964;
srom_1(86522) <= 15604635;
srom_1(86523) <= 15880467;
srom_1(86524) <= 16121167;
srom_1(86525) <= 16325607;
srom_1(86526) <= 16492827;
srom_1(86527) <= 16622044;
srom_1(86528) <= 16712652;
srom_1(86529) <= 16764225;
srom_1(86530) <= 16776522;
srom_1(86531) <= 16749486;
srom_1(86532) <= 16683242;
srom_1(86533) <= 16578102;
srom_1(86534) <= 16434558;
srom_1(86535) <= 16253284;
srom_1(86536) <= 16035130;
srom_1(86537) <= 15781119;
srom_1(86538) <= 15492442;
srom_1(86539) <= 15170453;
srom_1(86540) <= 14816661;
srom_1(86541) <= 14432726;
srom_1(86542) <= 14020447;
srom_1(86543) <= 13581760;
srom_1(86544) <= 13118719;
srom_1(86545) <= 12633498;
srom_1(86546) <= 12128371;
srom_1(86547) <= 11605706;
srom_1(86548) <= 11067956;
srom_1(86549) <= 10517641;
srom_1(86550) <= 9957343;
srom_1(86551) <= 9389688;
srom_1(86552) <= 8817339;
srom_1(86553) <= 8242979;
srom_1(86554) <= 7669302;
srom_1(86555) <= 7098999;
srom_1(86556) <= 6534742;
srom_1(86557) <= 5979179;
srom_1(86558) <= 5434915;
srom_1(86559) <= 4904502;
srom_1(86560) <= 4390426;
srom_1(86561) <= 3895100;
srom_1(86562) <= 3420845;
srom_1(86563) <= 2969886;
srom_1(86564) <= 2544337;
srom_1(86565) <= 2146194;
srom_1(86566) <= 1777323;
srom_1(86567) <= 1439455;
srom_1(86568) <= 1134174;
srom_1(86569) <= 862912;
srom_1(86570) <= 626940;
srom_1(86571) <= 427366;
srom_1(86572) <= 265124;
srom_1(86573) <= 140976;
srom_1(86574) <= 55504;
srom_1(86575) <= 9109;
srom_1(86576) <= 2008;
srom_1(86577) <= 34235;
srom_1(86578) <= 105638;
srom_1(86579) <= 215883;
srom_1(86580) <= 364453;
srom_1(86581) <= 550651;
srom_1(86582) <= 773604;
srom_1(86583) <= 1032266;
srom_1(86584) <= 1325424;
srom_1(86585) <= 1651704;
srom_1(86586) <= 2009576;
srom_1(86587) <= 2397361;
srom_1(86588) <= 2813241;
srom_1(86589) <= 3255266;
srom_1(86590) <= 3721363;
srom_1(86591) <= 4209347;
srom_1(86592) <= 4716928;
srom_1(86593) <= 5241727;
srom_1(86594) <= 5781283;
srom_1(86595) <= 6333065;
srom_1(86596) <= 6894487;
srom_1(86597) <= 7462915;
srom_1(86598) <= 8035684;
srom_1(86599) <= 8610108;
srom_1(86600) <= 9183493;
srom_1(86601) <= 9753151;
srom_1(86602) <= 10316410;
srom_1(86603) <= 10870629;
srom_1(86604) <= 11413209;
srom_1(86605) <= 11941605;
srom_1(86606) <= 12453340;
srom_1(86607) <= 12946014;
srom_1(86608) <= 13417317;
srom_1(86609) <= 13865039;
srom_1(86610) <= 14287079;
srom_1(86611) <= 14681460;
srom_1(86612) <= 15046332;
srom_1(86613) <= 15379983;
srom_1(86614) <= 15680849;
srom_1(86615) <= 15947519;
srom_1(86616) <= 16178743;
srom_1(86617) <= 16373436;
srom_1(86618) <= 16530686;
srom_1(86619) <= 16649754;
srom_1(86620) <= 16730084;
srom_1(86621) <= 16771297;
srom_1(86622) <= 16773201;
srom_1(86623) <= 16735787;
srom_1(86624) <= 16659229;
srom_1(86625) <= 16543889;
srom_1(86626) <= 16390305;
srom_1(86627) <= 16199198;
srom_1(86628) <= 15971465;
srom_1(86629) <= 15708173;
srom_1(86630) <= 15410558;
srom_1(86631) <= 15080014;
srom_1(86632) <= 14718091;
srom_1(86633) <= 14326488;
srom_1(86634) <= 13907040;
srom_1(86635) <= 13461714;
srom_1(86636) <= 12992598;
srom_1(86637) <= 12501893;
srom_1(86638) <= 11991899;
srom_1(86639) <= 11465008;
srom_1(86640) <= 10923691;
srom_1(86641) <= 10370485;
srom_1(86642) <= 9807987;
srom_1(86643) <= 9238832;
srom_1(86644) <= 8665690;
srom_1(86645) <= 8091249;
srom_1(86646) <= 7518202;
srom_1(86647) <= 6949237;
srom_1(86648) <= 6387021;
srom_1(86649) <= 5834192;
srom_1(86650) <= 5293341;
srom_1(86651) <= 4767005;
srom_1(86652) <= 4257652;
srom_1(86653) <= 3767671;
srom_1(86654) <= 3299358;
srom_1(86655) <= 2854911;
srom_1(86656) <= 2436413;
srom_1(86657) <= 2045827;
srom_1(86658) <= 1684985;
srom_1(86659) <= 1355578;
srom_1(86660) <= 1059151;
srom_1(86661) <= 797095;
srom_1(86662) <= 570638;
srom_1(86663) <= 380842;
srom_1(86664) <= 228597;
srom_1(86665) <= 114617;
srom_1(86666) <= 39437;
srom_1(86667) <= 3409;
srom_1(86668) <= 6702;
srom_1(86669) <= 49301;
srom_1(86670) <= 131006;
srom_1(86671) <= 251433;
srom_1(86672) <= 410018;
srom_1(86673) <= 606018;
srom_1(86674) <= 838513;
srom_1(86675) <= 1106413;
srom_1(86676) <= 1408461;
srom_1(86677) <= 1743242;
srom_1(86678) <= 2109185;
srom_1(86679) <= 2504575;
srom_1(86680) <= 2927557;
srom_1(86681) <= 3376148;
srom_1(86682) <= 3848243;
srom_1(86683) <= 4341630;
srom_1(86684) <= 4853995;
srom_1(86685) <= 5382935;
srom_1(86686) <= 5925969;
srom_1(86687) <= 6480552;
srom_1(86688) <= 7044082;
srom_1(86689) <= 7613917;
srom_1(86690) <= 8187385;
srom_1(86691) <= 8761796;
srom_1(86692) <= 9334457;
srom_1(86693) <= 9902683;
srom_1(86694) <= 10463809;
srom_1(86695) <= 11015204;
srom_1(86696) <= 11554281;
srom_1(86697) <= 12078514;
srom_1(86698) <= 12585443;
srom_1(86699) <= 13072692;
srom_1(86700) <= 13537976;
srom_1(86701) <= 13979113;
srom_1(86702) <= 14394033;
srom_1(86703) <= 14780792;
srom_1(86704) <= 15137577;
srom_1(86705) <= 15462712;
srom_1(86706) <= 15754675;
srom_1(86707) <= 16012096;
srom_1(86708) <= 16233768;
srom_1(86709) <= 16418651;
srom_1(86710) <= 16565878;
srom_1(86711) <= 16674760;
srom_1(86712) <= 16744784;
srom_1(86713) <= 16775624;
srom_1(86714) <= 16767134;
srom_1(86715) <= 16719355;
srom_1(86716) <= 16632509;
srom_1(86717) <= 16507005;
srom_1(86718) <= 16343432;
srom_1(86719) <= 16142555;
srom_1(86720) <= 15905317;
srom_1(86721) <= 15632831;
srom_1(86722) <= 15326374;
srom_1(86723) <= 14987384;
srom_1(86724) <= 14617450;
srom_1(86725) <= 14218306;
srom_1(86726) <= 13791825;
srom_1(86727) <= 13340007;
srom_1(86728) <= 12864970;
srom_1(86729) <= 12368941;
srom_1(86730) <= 11854247;
srom_1(86731) <= 11323302;
srom_1(86732) <= 10778595;
srom_1(86733) <= 10222681;
srom_1(86734) <= 9658166;
srom_1(86735) <= 9087697;
srom_1(86736) <= 8513950;
srom_1(86737) <= 7939616;
srom_1(86738) <= 7367387;
srom_1(86739) <= 6799946;
srom_1(86740) <= 6239956;
srom_1(86741) <= 5690041;
srom_1(86742) <= 5152781;
srom_1(86743) <= 4630695;
srom_1(86744) <= 4126230;
srom_1(86745) <= 3641754;
srom_1(86746) <= 3179537;
srom_1(86747) <= 2741748;
srom_1(86748) <= 2330438;
srom_1(86749) <= 1947537;
srom_1(86750) <= 1594841;
srom_1(86751) <= 1274003;
srom_1(86752) <= 986527;
srom_1(86753) <= 733763;
srom_1(86754) <= 516895;
srom_1(86755) <= 336940;
srom_1(86756) <= 194742;
srom_1(86757) <= 90968;
srom_1(86758) <= 26104;
srom_1(86759) <= 455;
srom_1(86760) <= 14141;
srom_1(86761) <= 67097;
srom_1(86762) <= 159076;
srom_1(86763) <= 289647;
srom_1(86764) <= 458196;
srom_1(86765) <= 663933;
srom_1(86766) <= 905894;
srom_1(86767) <= 1182944;
srom_1(86768) <= 1493784;
srom_1(86769) <= 1836956;
srom_1(86770) <= 2210851;
srom_1(86771) <= 2613715;
srom_1(86772) <= 3043661;
srom_1(86773) <= 3498670;
srom_1(86774) <= 3976610;
srom_1(86775) <= 4475239;
srom_1(86776) <= 4992220;
srom_1(86777) <= 5525127;
srom_1(86778) <= 6071462;
srom_1(86779) <= 6628663;
srom_1(86780) <= 7194117;
srom_1(86781) <= 7765172;
srom_1(86782) <= 8339151;
srom_1(86783) <= 8913362;
srom_1(86784) <= 9485112;
srom_1(86785) <= 10051720;
srom_1(86786) <= 10610529;
srom_1(86787) <= 11158919;
srom_1(86788) <= 11694318;
srom_1(86789) <= 12214215;
srom_1(86790) <= 12716173;
srom_1(86791) <= 13197837;
srom_1(86792) <= 13656949;
srom_1(86793) <= 14091356;
srom_1(86794) <= 14499021;
srom_1(86795) <= 14878032;
srom_1(86796) <= 15226612;
srom_1(86797) <= 15543126;
srom_1(86798) <= 15826090;
srom_1(86799) <= 16074177;
srom_1(86800) <= 16286224;
srom_1(86801) <= 16461237;
srom_1(86802) <= 16598394;
srom_1(86803) <= 16697052;
srom_1(86804) <= 16756749;
srom_1(86805) <= 16777206;
srom_1(86806) <= 16758325;
srom_1(86807) <= 16700195;
srom_1(86808) <= 16603090;
srom_1(86809) <= 16467465;
srom_1(86810) <= 16293954;
srom_1(86811) <= 16083373;
srom_1(86812) <= 15836708;
srom_1(86813) <= 15555117;
srom_1(86814) <= 15239920;
srom_1(86815) <= 14892594;
srom_1(86816) <= 14514769;
srom_1(86817) <= 14108216;
srom_1(86818) <= 13674842;
srom_1(86819) <= 13216679;
srom_1(86820) <= 12735876;
srom_1(86821) <= 12234686;
srom_1(86822) <= 11715461;
srom_1(86823) <= 11180636;
srom_1(86824) <= 10632717;
srom_1(86825) <= 10074275;
srom_1(86826) <= 9507929;
srom_1(86827) <= 8936333;
srom_1(86828) <= 8362170;
srom_1(86829) <= 7788130;
srom_1(86830) <= 7216905;
srom_1(86831) <= 6651176;
srom_1(86832) <= 6093594;
srom_1(86833) <= 5546774;
srom_1(86834) <= 5013280;
srom_1(86835) <= 4495614;
srom_1(86836) <= 3996204;
srom_1(86837) <= 3517392;
srom_1(86838) <= 3061422;
srom_1(86839) <= 2630433;
srom_1(86840) <= 2226446;
srom_1(86841) <= 1851356;
srom_1(86842) <= 1506921;
srom_1(86843) <= 1194757;
srom_1(86844) <= 916327;
srom_1(86845) <= 672937;
srom_1(86846) <= 465729;
srom_1(86847) <= 295674;
srom_1(86848) <= 163569;
srom_1(86849) <= 70034;
srom_1(86850) <= 15508;
srom_1(86851) <= 247;
srom_1(86852) <= 24321;
srom_1(86853) <= 87618;
srom_1(86854) <= 189841;
srom_1(86855) <= 330512;
srom_1(86856) <= 508969;
srom_1(86857) <= 724377;
srom_1(86858) <= 975725;
srom_1(86859) <= 1261834;
srom_1(86860) <= 1581364;
srom_1(86861) <= 1932815;
srom_1(86862) <= 2314539;
srom_1(86863) <= 2724747;
srom_1(86864) <= 3161514;
srom_1(86865) <= 3622793;
srom_1(86866) <= 4106421;
srom_1(86867) <= 4610129;
srom_1(86868) <= 5131556;
srom_1(86869) <= 5668256;
srom_1(86870) <= 6217713;
srom_1(86871) <= 6777350;
srom_1(86872) <= 7344543;
srom_1(86873) <= 7916632;
srom_1(86874) <= 8490934;
srom_1(86875) <= 9064756;
srom_1(86876) <= 9635407;
srom_1(86877) <= 10200212;
srom_1(86878) <= 10756522;
srom_1(86879) <= 11301727;
srom_1(86880) <= 11833272;
srom_1(86881) <= 12348664;
srom_1(86882) <= 12845485;
srom_1(86883) <= 13321407;
srom_1(86884) <= 13774197;
srom_1(86885) <= 14201733;
srom_1(86886) <= 14602008;
srom_1(86887) <= 14973147;
srom_1(86888) <= 15313409;
srom_1(86889) <= 15621198;
srom_1(86890) <= 15895070;
srom_1(86891) <= 16133743;
srom_1(86892) <= 16336095;
srom_1(86893) <= 16501180;
srom_1(86894) <= 16628221;
srom_1(86895) <= 16716624;
srom_1(86896) <= 16765975;
srom_1(86897) <= 16776041;
srom_1(86898) <= 16746775;
srom_1(86899) <= 16678315;
srom_1(86900) <= 16570982;
srom_1(86901) <= 16425279;
srom_1(86902) <= 16241889;
srom_1(86903) <= 16021672;
srom_1(86904) <= 15765661;
srom_1(86905) <= 15475057;
srom_1(86906) <= 15151222;
srom_1(86907) <= 14795675;
srom_1(86908) <= 14410082;
srom_1(86909) <= 13996253;
srom_1(86910) <= 13556128;
srom_1(86911) <= 13091771;
srom_1(86912) <= 12605358;
srom_1(86913) <= 12099172;
srom_1(86914) <= 11575586;
srom_1(86915) <= 11037055;
srom_1(86916) <= 10486105;
srom_1(86917) <= 9925318;
srom_1(86918) <= 9357326;
srom_1(86919) <= 8784791;
srom_1(86920) <= 8210397;
srom_1(86921) <= 7636840;
srom_1(86922) <= 7066808;
srom_1(86923) <= 6502974;
srom_1(86924) <= 5947983;
srom_1(86925) <= 5404437;
srom_1(86926) <= 4874884;
srom_1(86927) <= 4361808;
srom_1(86928) <= 3867616;
srom_1(86929) <= 3394624;
srom_1(86930) <= 2945050;
srom_1(86931) <= 2521003;
srom_1(86932) <= 2124472;
srom_1(86933) <= 1757315;
srom_1(86934) <= 1421254;
srom_1(86935) <= 1117866;
srom_1(86936) <= 848573;
srom_1(86937) <= 614637;
srom_1(86938) <= 417157;
srom_1(86939) <= 257057;
srom_1(86940) <= 135089;
srom_1(86941) <= 51824;
srom_1(86942) <= 7654;
srom_1(86943) <= 2785;
srom_1(86944) <= 37239;
srom_1(86945) <= 110856;
srom_1(86946) <= 223291;
srom_1(86947) <= 374015;
srom_1(86948) <= 562322;
srom_1(86949) <= 787330;
srom_1(86950) <= 1047983;
srom_1(86951) <= 1343058;
srom_1(86952) <= 1671172;
srom_1(86953) <= 2030787;
srom_1(86954) <= 2420215;
srom_1(86955) <= 2837632;
srom_1(86956) <= 3281079;
srom_1(86957) <= 3748477;
srom_1(86958) <= 4237634;
srom_1(86959) <= 4746256;
srom_1(86960) <= 5271959;
srom_1(86961) <= 5812276;
srom_1(86962) <= 6364675;
srom_1(86963) <= 6926565;
srom_1(86964) <= 7495311;
srom_1(86965) <= 8068246;
srom_1(86966) <= 8642683;
srom_1(86967) <= 9215928;
srom_1(86968) <= 9785295;
srom_1(86969) <= 10348111;
srom_1(86970) <= 10901739;
srom_1(86971) <= 11443581;
srom_1(86972) <= 11971098;
srom_1(86973) <= 12481816;
srom_1(86974) <= 12973339;
srom_1(86975) <= 13443362;
srom_1(86976) <= 13889682;
srom_1(86977) <= 14310206;
srom_1(86978) <= 14702961;
srom_1(86979) <= 15066106;
srom_1(86980) <= 15397938;
srom_1(86981) <= 15696901;
srom_1(86982) <= 15961593;
srom_1(86983) <= 16190772;
srom_1(86984) <= 16383364;
srom_1(86985) <= 16538467;
srom_1(86986) <= 16655351;
srom_1(86987) <= 16733470;
srom_1(86988) <= 16772457;
srom_1(86989) <= 16772130;
srom_1(86990) <= 16732489;
srom_1(86991) <= 16653721;
srom_1(86992) <= 16536195;
srom_1(86993) <= 16380462;
srom_1(86994) <= 16187252;
srom_1(86995) <= 15957472;
srom_1(86996) <= 15692199;
srom_1(86997) <= 15392677;
srom_1(86998) <= 15060310;
srom_1(86999) <= 14696658;
srom_1(87000) <= 14303424;
srom_1(87001) <= 13882455;
srom_1(87002) <= 13435722;
srom_1(87003) <= 12965322;
srom_1(87004) <= 12473461;
srom_1(87005) <= 11962443;
srom_1(87006) <= 11434667;
srom_1(87007) <= 10892607;
srom_1(87008) <= 10338805;
srom_1(87009) <= 9775858;
srom_1(87010) <= 9206405;
srom_1(87011) <= 8633118;
srom_1(87012) <= 8058684;
srom_1(87013) <= 7485797;
srom_1(87014) <= 6917143;
srom_1(87015) <= 6355390;
srom_1(87016) <= 5803171;
srom_1(87017) <= 5263076;
srom_1(87018) <= 4737638;
srom_1(87019) <= 4229321;
srom_1(87020) <= 3740508;
srom_1(87021) <= 3273491;
srom_1(87022) <= 2830461;
srom_1(87023) <= 2413495;
srom_1(87024) <= 2024548;
srom_1(87025) <= 1665445;
srom_1(87026) <= 1337869;
srom_1(87027) <= 1043356;
srom_1(87028) <= 783287;
srom_1(87029) <= 558883;
srom_1(87030) <= 371195;
srom_1(87031) <= 221103;
srom_1(87032) <= 109311;
srom_1(87033) <= 36344;
srom_1(87034) <= 2544;
srom_1(87035) <= 8068;
srom_1(87036) <= 52892;
srom_1(87037) <= 136805;
srom_1(87038) <= 259413;
srom_1(87039) <= 420142;
srom_1(87040) <= 618238;
srom_1(87041) <= 852772;
srom_1(87042) <= 1122644;
srom_1(87043) <= 1426588;
srom_1(87044) <= 1763180;
srom_1(87045) <= 2130841;
srom_1(87046) <= 2527846;
srom_1(87047) <= 2952335;
srom_1(87048) <= 3402316;
srom_1(87049) <= 3875679;
srom_1(87050) <= 4370206;
srom_1(87051) <= 4883576;
srom_1(87052) <= 5413382;
srom_1(87053) <= 5957140;
srom_1(87054) <= 6512300;
srom_1(87055) <= 7076258;
srom_1(87056) <= 7646371;
srom_1(87057) <= 8219965;
srom_1(87058) <= 8794349;
srom_1(87059) <= 9366830;
srom_1(87060) <= 9934724;
srom_1(87061) <= 10495368;
srom_1(87062) <= 11046133;
srom_1(87063) <= 11584436;
srom_1(87064) <= 12107752;
srom_1(87065) <= 12613628;
srom_1(87066) <= 13099691;
srom_1(87067) <= 13563663;
srom_1(87068) <= 14003366;
srom_1(87069) <= 14416741;
srom_1(87070) <= 14801847;
srom_1(87071) <= 15156879;
srom_1(87072) <= 15480173;
srom_1(87073) <= 15770212;
srom_1(87074) <= 16025636;
srom_1(87075) <= 16245247;
srom_1(87076) <= 16428016;
srom_1(87077) <= 16573085;
srom_1(87078) <= 16679775;
srom_1(87079) <= 16747584;
srom_1(87080) <= 16776195;
srom_1(87081) <= 16765474;
srom_1(87082) <= 16715471;
srom_1(87083) <= 16626420;
srom_1(87084) <= 16498740;
srom_1(87085) <= 16333028;
srom_1(87086) <= 16130062;
srom_1(87087) <= 15890794;
srom_1(87088) <= 15616345;
srom_1(87089) <= 15308003;
srom_1(87090) <= 14967214;
srom_1(87091) <= 14595575;
srom_1(87092) <= 14194830;
srom_1(87093) <= 13766857;
srom_1(87094) <= 13313664;
srom_1(87095) <= 12837376;
srom_1(87096) <= 12340225;
srom_1(87097) <= 11824545;
srom_1(87098) <= 11292752;
srom_1(87099) <= 10747340;
srom_1(87100) <= 10190868;
srom_1(87101) <= 9625944;
srom_1(87102) <= 9055217;
srom_1(87103) <= 8481365;
srom_1(87104) <= 7907078;
srom_1(87105) <= 7335049;
srom_1(87106) <= 6767960;
srom_1(87107) <= 6208471;
srom_1(87108) <= 5659206;
srom_1(87109) <= 5122740;
srom_1(87110) <= 4601588;
srom_1(87111) <= 4098195;
srom_1(87112) <= 3614921;
srom_1(87113) <= 3154033;
srom_1(87114) <= 2717692;
srom_1(87115) <= 2307943;
srom_1(87116) <= 1926708;
srom_1(87117) <= 1575776;
srom_1(87118) <= 1256792;
srom_1(87119) <= 971250;
srom_1(87120) <= 720492;
srom_1(87121) <= 505692;
srom_1(87122) <= 327857;
srom_1(87123) <= 187822;
srom_1(87124) <= 86244;
srom_1(87125) <= 23598;
srom_1(87126) <= 179;
srom_1(87127) <= 16095;
srom_1(87128) <= 71274;
srom_1(87129) <= 165455;
srom_1(87130) <= 298197;
srom_1(87131) <= 468878;
srom_1(87132) <= 676697;
srom_1(87133) <= 920681;
srom_1(87134) <= 1199683;
srom_1(87135) <= 1512398;
srom_1(87136) <= 1857357;
srom_1(87137) <= 2232943;
srom_1(87138) <= 2637395;
srom_1(87139) <= 3068817;
srom_1(87140) <= 3525185;
srom_1(87141) <= 4004360;
srom_1(87142) <= 4504093;
srom_1(87143) <= 5022042;
srom_1(87144) <= 5555779;
srom_1(87145) <= 6102799;
srom_1(87146) <= 6660539;
srom_1(87147) <= 7226382;
srom_1(87148) <= 7797675;
srom_1(87149) <= 8371739;
srom_1(87150) <= 8945882;
srom_1(87151) <= 9517412;
srom_1(87152) <= 10083648;
srom_1(87153) <= 10641936;
srom_1(87154) <= 11189657;
srom_1(87155) <= 11724244;
srom_1(87156) <= 12243188;
srom_1(87157) <= 12744057;
srom_1(87158) <= 13224501;
srom_1(87159) <= 13682269;
srom_1(87160) <= 14115212;
srom_1(87161) <= 14521302;
srom_1(87162) <= 14898633;
srom_1(87163) <= 15245437;
srom_1(87164) <= 15560086;
srom_1(87165) <= 15841106;
srom_1(87166) <= 16087179;
srom_1(87167) <= 16297150;
srom_1(87168) <= 16470036;
srom_1(87169) <= 16605024;
srom_1(87170) <= 16701484;
srom_1(87171) <= 16758961;
srom_1(87172) <= 16777187;
srom_1(87173) <= 16756076;
srom_1(87174) <= 16695727;
srom_1(87175) <= 16596423;
srom_1(87176) <= 16458630;
srom_1(87177) <= 16282994;
srom_1(87178) <= 16070338;
srom_1(87179) <= 15821660;
srom_1(87180) <= 15538125;
srom_1(87181) <= 15221065;
srom_1(87182) <= 14871964;
srom_1(87183) <= 14492461;
srom_1(87184) <= 14084335;
srom_1(87185) <= 13649499;
srom_1(87186) <= 13189993;
srom_1(87187) <= 12707972;
srom_1(87188) <= 12205697;
srom_1(87189) <= 11685521;
srom_1(87190) <= 11149885;
srom_1(87191) <= 10601300;
srom_1(87192) <= 10042340;
srom_1(87193) <= 9475624;
srom_1(87194) <= 8903811;
srom_1(87195) <= 8329582;
srom_1(87196) <= 7755630;
srom_1(87197) <= 7184646;
srom_1(87198) <= 6619308;
srom_1(87199) <= 6062267;
srom_1(87200) <= 5516134;
srom_1(87201) <= 4983472;
srom_1(87202) <= 4466778;
srom_1(87203) <= 3968474;
srom_1(87204) <= 3490898;
srom_1(87205) <= 3036289;
srom_1(87206) <= 2606779;
srom_1(87207) <= 2204381;
srom_1(87208) <= 1830984;
srom_1(87209) <= 1488338;
srom_1(87210) <= 1178049;
srom_1(87211) <= 901573;
srom_1(87212) <= 660207;
srom_1(87213) <= 455081;
srom_1(87214) <= 287159;
srom_1(87215) <= 157227;
srom_1(87216) <= 65895;
srom_1(87217) <= 13591;
srom_1(87218) <= 560;
srom_1(87219) <= 26864;
srom_1(87220) <= 92378;
srom_1(87221) <= 196797;
srom_1(87222) <= 339630;
srom_1(87223) <= 520207;
srom_1(87224) <= 737682;
srom_1(87225) <= 991034;
srom_1(87226) <= 1279077;
srom_1(87227) <= 1600458;
srom_1(87228) <= 1953672;
srom_1(87229) <= 2337061;
srom_1(87230) <= 2748828;
srom_1(87231) <= 3187041;
srom_1(87232) <= 3649647;
srom_1(87233) <= 4134475;
srom_1(87234) <= 4639252;
srom_1(87235) <= 5161612;
srom_1(87236) <= 5699103;
srom_1(87237) <= 6249207;
srom_1(87238) <= 6809343;
srom_1(87239) <= 7376885;
srom_1(87240) <= 7949171;
srom_1(87241) <= 8523518;
srom_1(87242) <= 9097232;
srom_1(87243) <= 9667624;
srom_1(87244) <= 10232017;
srom_1(87245) <= 10787766;
srom_1(87246) <= 11332265;
srom_1(87247) <= 11862960;
srom_1(87248) <= 12377362;
srom_1(87249) <= 12873060;
srom_1(87250) <= 13347728;
srom_1(87251) <= 13799142;
srom_1(87252) <= 14225183;
srom_1(87253) <= 14623855;
srom_1(87254) <= 14993288;
srom_1(87255) <= 15331749;
srom_1(87256) <= 15637651;
srom_1(87257) <= 15909560;
srom_1(87258) <= 16146201;
srom_1(87259) <= 16346464;
srom_1(87260) <= 16509409;
srom_1(87261) <= 16634274;
srom_1(87262) <= 16720471;
srom_1(87263) <= 16767598;
srom_1(87264) <= 16775432;
srom_1(87265) <= 16743938;
srom_1(87266) <= 16673263;
srom_1(87267) <= 16563739;
srom_1(87268) <= 16415878;
srom_1(87269) <= 16230374;
srom_1(87270) <= 16008098;
srom_1(87271) <= 15750092;
srom_1(87272) <= 15457565;
srom_1(87273) <= 15131889;
srom_1(87274) <= 14774592;
srom_1(87275) <= 14387348;
srom_1(87276) <= 13971975;
srom_1(87277) <= 13530419;
srom_1(87278) <= 13064751;
srom_1(87279) <= 12577155;
srom_1(87280) <= 12069918;
srom_1(87281) <= 11545418;
srom_1(87282) <= 11006114;
srom_1(87283) <= 10454536;
srom_1(87284) <= 9893270;
srom_1(87285) <= 9324949;
srom_1(87286) <= 8752236;
srom_1(87287) <= 8177818;
srom_1(87288) <= 7604389;
srom_1(87289) <= 7034637;
srom_1(87290) <= 6471235;
srom_1(87291) <= 5916823;
srom_1(87292) <= 5374003;
srom_1(87293) <= 4845319;
srom_1(87294) <= 4333251;
srom_1(87295) <= 3840200;
srom_1(87296) <= 3368478;
srom_1(87297) <= 2920297;
srom_1(87298) <= 2497759;
srom_1(87299) <= 2102845;
srom_1(87300) <= 1737407;
srom_1(87301) <= 1403159;
srom_1(87302) <= 1101668;
srom_1(87303) <= 834347;
srom_1(87304) <= 602452;
srom_1(87305) <= 407068;
srom_1(87306) <= 249113;
srom_1(87307) <= 129326;
srom_1(87308) <= 48271;
srom_1(87309) <= 6325;
srom_1(87310) <= 3688;
srom_1(87311) <= 40370;
srom_1(87312) <= 116199;
srom_1(87313) <= 230821;
srom_1(87314) <= 383698;
srom_1(87315) <= 574112;
srom_1(87316) <= 801171;
srom_1(87317) <= 1063810;
srom_1(87318) <= 1360798;
srom_1(87319) <= 1690741;
srom_1(87320) <= 2052094;
srom_1(87321) <= 2443160;
srom_1(87322) <= 2862106;
srom_1(87323) <= 3306968;
srom_1(87324) <= 3775660;
srom_1(87325) <= 4265983;
srom_1(87326) <= 4775639;
srom_1(87327) <= 5302237;
srom_1(87328) <= 5843308;
srom_1(87329) <= 6396316;
srom_1(87330) <= 6958665;
srom_1(87331) <= 7527720;
srom_1(87332) <= 8100812;
srom_1(87333) <= 8675254;
srom_1(87334) <= 9248351;
srom_1(87335) <= 9817417;
srom_1(87336) <= 10379782;
srom_1(87337) <= 10932811;
srom_1(87338) <= 11473908;
srom_1(87339) <= 12000538;
srom_1(87340) <= 12510230;
srom_1(87341) <= 13000594;
srom_1(87342) <= 13469331;
srom_1(87343) <= 13914243;
srom_1(87344) <= 14333243;
srom_1(87345) <= 14724367;
srom_1(87346) <= 15085780;
srom_1(87347) <= 15415788;
srom_1(87348) <= 15712843;
srom_1(87349) <= 15975552;
srom_1(87350) <= 16202684;
srom_1(87351) <= 16393172;
srom_1(87352) <= 16546124;
srom_1(87353) <= 16660823;
srom_1(87354) <= 16736731;
srom_1(87355) <= 16773491;
srom_1(87356) <= 16770932;
srom_1(87357) <= 16729065;
srom_1(87358) <= 16648087;
srom_1(87359) <= 16528378;
srom_1(87360) <= 16370498;
srom_1(87361) <= 16175188;
srom_1(87362) <= 15943365;
srom_1(87363) <= 15676114;
srom_1(87364) <= 15374690;
srom_1(87365) <= 15040506;
srom_1(87366) <= 14675128;
srom_1(87367) <= 14280272;
srom_1(87368) <= 13857787;
srom_1(87369) <= 13409655;
srom_1(87370) <= 12937977;
srom_1(87371) <= 12444967;
srom_1(87372) <= 11932934;
srom_1(87373) <= 11404281;
srom_1(87374) <= 10861487;
srom_1(87375) <= 10307096;
srom_1(87376) <= 9743708;
srom_1(87377) <= 9173967;
srom_1(87378) <= 8600542;
srom_1(87379) <= 8026124;
srom_1(87380) <= 7453405;
srom_1(87381) <= 6885072;
srom_1(87382) <= 6323789;
srom_1(87383) <= 5772189;
srom_1(87384) <= 5232859;
srom_1(87385) <= 4708327;
srom_1(87386) <= 4201052;
srom_1(87387) <= 3713415;
srom_1(87388) <= 3247701;
srom_1(87389) <= 2806095;
srom_1(87390) <= 2390667;
srom_1(87391) <= 2003366;
srom_1(87392) <= 1646007;
srom_1(87393) <= 1320266;
srom_1(87394) <= 1027672;
srom_1(87395) <= 769595;
srom_1(87396) <= 547246;
srom_1(87397) <= 361669;
srom_1(87398) <= 213732;
srom_1(87399) <= 104130;
srom_1(87400) <= 33377;
srom_1(87401) <= 1804;
srom_1(87402) <= 9560;
srom_1(87403) <= 56609;
srom_1(87404) <= 142728;
srom_1(87405) <= 267516;
srom_1(87406) <= 430386;
srom_1(87407) <= 630575;
srom_1(87408) <= 867144;
srom_1(87409) <= 1138984;
srom_1(87410) <= 1444820;
srom_1(87411) <= 1783217;
srom_1(87412) <= 2152590;
srom_1(87413) <= 2551205;
srom_1(87414) <= 2977194;
srom_1(87415) <= 3428559;
srom_1(87416) <= 3903183;
srom_1(87417) <= 4398841;
srom_1(87418) <= 4913209;
srom_1(87419) <= 5443873;
srom_1(87420) <= 5988347;
srom_1(87421) <= 6544076;
srom_1(87422) <= 7108455;
srom_1(87423) <= 7678837;
srom_1(87424) <= 8252547;
srom_1(87425) <= 8826895;
srom_1(87426) <= 9399188;
srom_1(87427) <= 9966742;
srom_1(87428) <= 10526896;
srom_1(87429) <= 11077022;
srom_1(87430) <= 11614542;
srom_1(87431) <= 12136934;
srom_1(87432) <= 12641749;
srom_1(87433) <= 13126619;
srom_1(87434) <= 13589271;
srom_1(87435) <= 14027536;
srom_1(87436) <= 14439357;
srom_1(87437) <= 14822805;
srom_1(87438) <= 15176080;
srom_1(87439) <= 15497527;
srom_1(87440) <= 15785637;
srom_1(87441) <= 16039060;
srom_1(87442) <= 16256608;
srom_1(87443) <= 16437260;
srom_1(87444) <= 16580169;
srom_1(87445) <= 16684665;
srom_1(87446) <= 16750258;
srom_1(87447) <= 16776640;
srom_1(87448) <= 16763687;
srom_1(87449) <= 16711462;
srom_1(87450) <= 16620207;
srom_1(87451) <= 16490352;
srom_1(87452) <= 16322504;
srom_1(87453) <= 16117452;
srom_1(87454) <= 15876157;
srom_1(87455) <= 15599750;
srom_1(87456) <= 15289528;
srom_1(87457) <= 14946945;
srom_1(87458) <= 14573607;
srom_1(87459) <= 14171266;
srom_1(87460) <= 13741808;
srom_1(87461) <= 13287247;
srom_1(87462) <= 12809715;
srom_1(87463) <= 12311450;
srom_1(87464) <= 11794790;
srom_1(87465) <= 11262157;
srom_1(87466) <= 10716049;
srom_1(87467) <= 10159027;
srom_1(87468) <= 9593703;
srom_1(87469) <= 9022728;
srom_1(87470) <= 8448779;
srom_1(87471) <= 7874548;
srom_1(87472) <= 7302727;
srom_1(87473) <= 6735999;
srom_1(87474) <= 6177020;
srom_1(87475) <= 5628412;
srom_1(87476) <= 5092748;
srom_1(87477) <= 4572539;
srom_1(87478) <= 4070225;
srom_1(87479) <= 3588161;
srom_1(87480) <= 3128608;
srom_1(87481) <= 2693721;
srom_1(87482) <= 2285540;
srom_1(87483) <= 1905977;
srom_1(87484) <= 1556814;
srom_1(87485) <= 1239688;
srom_1(87486) <= 956085;
srom_1(87487) <= 707337;
srom_1(87488) <= 494608;
srom_1(87489) <= 318897;
srom_1(87490) <= 181027;
srom_1(87491) <= 81646;
srom_1(87492) <= 21219;
srom_1(87493) <= 29;
srom_1(87494) <= 18176;
srom_1(87495) <= 75575;
srom_1(87496) <= 171957;
srom_1(87497) <= 306870;
srom_1(87498) <= 479680;
srom_1(87499) <= 689578;
srom_1(87500) <= 935580;
srom_1(87501) <= 1216531;
srom_1(87502) <= 1531115;
srom_1(87503) <= 1877856;
srom_1(87504) <= 2255128;
srom_1(87505) <= 2661162;
srom_1(87506) <= 3094054;
srom_1(87507) <= 3551774;
srom_1(87508) <= 4032175;
srom_1(87509) <= 4533006;
srom_1(87510) <= 5051916;
srom_1(87511) <= 5586474;
srom_1(87512) <= 6134171;
srom_1(87513) <= 6692441;
srom_1(87514) <= 7258664;
srom_1(87515) <= 7830186;
srom_1(87516) <= 8404326;
srom_1(87517) <= 8978393;
srom_1(87518) <= 9549695;
srom_1(87519) <= 10115551;
srom_1(87520) <= 10673309;
srom_1(87521) <= 11220354;
srom_1(87522) <= 11754119;
srom_1(87523) <= 12272102;
srom_1(87524) <= 12771875;
srom_1(87525) <= 13251092;
srom_1(87526) <= 13707508;
srom_1(87527) <= 14138982;
srom_1(87528) <= 14543490;
srom_1(87529) <= 14919136;
srom_1(87530) <= 15264158;
srom_1(87531) <= 15576938;
srom_1(87532) <= 15856009;
srom_1(87533) <= 16100064;
srom_1(87534) <= 16307956;
srom_1(87535) <= 16478712;
srom_1(87536) <= 16611531;
srom_1(87537) <= 16705790;
srom_1(87538) <= 16761047;
srom_1(87539) <= 16777042;
srom_1(87540) <= 16753701;
srom_1(87541) <= 16691133;
srom_1(87542) <= 16589632;
srom_1(87543) <= 16449673;
srom_1(87544) <= 16271914;
srom_1(87545) <= 16057186;
srom_1(87546) <= 15806499;
srom_1(87547) <= 15521026;
srom_1(87548) <= 15202107;
srom_1(87549) <= 14851236;
srom_1(87550) <= 14470061;
srom_1(87551) <= 14060367;
srom_1(87552) <= 13624077;
srom_1(87553) <= 13163235;
srom_1(87554) <= 12680004;
srom_1(87555) <= 12176649;
srom_1(87556) <= 11655531;
srom_1(87557) <= 11119092;
srom_1(87558) <= 10569850;
srom_1(87559) <= 10010379;
srom_1(87560) <= 9443303;
srom_1(87561) <= 8871281;
srom_1(87562) <= 8296996;
srom_1(87563) <= 7723140;
srom_1(87564) <= 7152405;
srom_1(87565) <= 6587467;
srom_1(87566) <= 6030975;
srom_1(87567) <= 5485538;
srom_1(87568) <= 4953716;
srom_1(87569) <= 4438000;
srom_1(87570) <= 3940811;
srom_1(87571) <= 3464478;
srom_1(87572) <= 3011237;
srom_1(87573) <= 2583212;
srom_1(87574) <= 2182410;
srom_1(87575) <= 1810711;
srom_1(87576) <= 1469859;
srom_1(87577) <= 1161450;
srom_1(87578) <= 886933;
srom_1(87579) <= 647593;
srom_1(87580) <= 444554;
srom_1(87581) <= 278767;
srom_1(87582) <= 151009;
srom_1(87583) <= 61881;
srom_1(87584) <= 11800;
srom_1(87585) <= 1000;
srom_1(87586) <= 29533;
srom_1(87587) <= 97264;
srom_1(87588) <= 203876;
srom_1(87589) <= 348869;
srom_1(87590) <= 531564;
srom_1(87591) <= 751102;
srom_1(87592) <= 1006456;
srom_1(87593) <= 1296427;
srom_1(87594) <= 1619655;
srom_1(87595) <= 1974626;
srom_1(87596) <= 2359674;
srom_1(87597) <= 2772994;
srom_1(87598) <= 3212647;
srom_1(87599) <= 3676572;
srom_1(87600) <= 4162593;
srom_1(87601) <= 4668432;
srom_1(87602) <= 5191716;
srom_1(87603) <= 5729991;
srom_1(87604) <= 6280733;
srom_1(87605) <= 6841360;
srom_1(87606) <= 7409243;
srom_1(87607) <= 7981718;
srom_1(87608) <= 8556101;
srom_1(87609) <= 9129698;
srom_1(87610) <= 9699821;
srom_1(87611) <= 10263794;
srom_1(87612) <= 10818975;
srom_1(87613) <= 11362758;
srom_1(87614) <= 11892595;
srom_1(87615) <= 12406000;
srom_1(87616) <= 12900566;
srom_1(87617) <= 13373974;
srom_1(87618) <= 13824004;
srom_1(87619) <= 14248546;
srom_1(87620) <= 14645608;
srom_1(87621) <= 15013329;
srom_1(87622) <= 15349985;
srom_1(87623) <= 15653996;
srom_1(87624) <= 15923937;
srom_1(87625) <= 16158542;
srom_1(87626) <= 16356712;
srom_1(87627) <= 16517517;
srom_1(87628) <= 16640202;
srom_1(87629) <= 16724192;
srom_1(87630) <= 16769094;
srom_1(87631) <= 16774698;
srom_1(87632) <= 16740976;
srom_1(87633) <= 16668086;
srom_1(87634) <= 16556372;
srom_1(87635) <= 16406356;
srom_1(87636) <= 16218742;
srom_1(87637) <= 15994410;
srom_1(87638) <= 15734411;
srom_1(87639) <= 15439966;
srom_1(87640) <= 15112454;
srom_1(87641) <= 14753412;
srom_1(87642) <= 14364524;
srom_1(87643) <= 13947612;
srom_1(87644) <= 13504632;
srom_1(87645) <= 13037661;
srom_1(87646) <= 12548889;
srom_1(87647) <= 12040608;
srom_1(87648) <= 11515202;
srom_1(87649) <= 10975134;
srom_1(87650) <= 10422937;
srom_1(87651) <= 9861200;
srom_1(87652) <= 9292558;
srom_1(87653) <= 8719676;
srom_1(87654) <= 8145243;
srom_1(87655) <= 7571950;
srom_1(87656) <= 7002487;
srom_1(87657) <= 6439524;
srom_1(87658) <= 5885701;
srom_1(87659) <= 5343615;
srom_1(87660) <= 4815808;
srom_1(87661) <= 4304755;
srom_1(87662) <= 3812853;
srom_1(87663) <= 3342408;
srom_1(87664) <= 2895626;
srom_1(87665) <= 2474603;
srom_1(87666) <= 2081312;
srom_1(87667) <= 1717599;
srom_1(87668) <= 1385168;
srom_1(87669) <= 1085579;
srom_1(87670) <= 820236;
srom_1(87671) <= 590384;
srom_1(87672) <= 397100;
srom_1(87673) <= 241292;
srom_1(87674) <= 123689;
srom_1(87675) <= 44843;
srom_1(87676) <= 5123;
srom_1(87677) <= 4717;
srom_1(87678) <= 43626;
srom_1(87679) <= 121667;
srom_1(87680) <= 238475;
srom_1(87681) <= 393501;
srom_1(87682) <= 586019;
srom_1(87683) <= 815127;
srom_1(87684) <= 1079748;
srom_1(87685) <= 1378644;
srom_1(87686) <= 1710412;
srom_1(87687) <= 2073496;
srom_1(87688) <= 2466194;
srom_1(87689) <= 2886664;
srom_1(87690) <= 3332935;
srom_1(87691) <= 3802913;
srom_1(87692) <= 4294395;
srom_1(87693) <= 4805077;
srom_1(87694) <= 5332562;
srom_1(87695) <= 5874379;
srom_1(87696) <= 6427986;
srom_1(87697) <= 6990787;
srom_1(87698) <= 7560142;
srom_1(87699) <= 8133383;
srom_1(87700) <= 8707820;
srom_1(87701) <= 9280761;
srom_1(87702) <= 9849518;
srom_1(87703) <= 10411424;
srom_1(87704) <= 10963844;
srom_1(87705) <= 11504189;
srom_1(87706) <= 12029923;
srom_1(87707) <= 12538582;
srom_1(87708) <= 13027780;
srom_1(87709) <= 13495224;
srom_1(87710) <= 13938720;
srom_1(87711) <= 14356191;
srom_1(87712) <= 14745677;
srom_1(87713) <= 15105353;
srom_1(87714) <= 15433532;
srom_1(87715) <= 15728675;
srom_1(87716) <= 15989397;
srom_1(87717) <= 16214477;
srom_1(87718) <= 16402859;
srom_1(87719) <= 16553659;
srom_1(87720) <= 16666171;
srom_1(87721) <= 16739866;
srom_1(87722) <= 16774399;
srom_1(87723) <= 16769608;
srom_1(87724) <= 16725516;
srom_1(87725) <= 16642329;
srom_1(87726) <= 16520438;
srom_1(87727) <= 16360414;
srom_1(87728) <= 16163007;
srom_1(87729) <= 15929143;
srom_1(87730) <= 15659919;
srom_1(87731) <= 15356598;
srom_1(87732) <= 15020601;
srom_1(87733) <= 14653505;
srom_1(87734) <= 14257030;
srom_1(87735) <= 13833036;
srom_1(87736) <= 13383511;
srom_1(87737) <= 12910564;
srom_1(87738) <= 12416412;
srom_1(87739) <= 11903371;
srom_1(87740) <= 11373849;
srom_1(87741) <= 10830328;
srom_1(87742) <= 10275357;
srom_1(87743) <= 9711539;
srom_1(87744) <= 9141516;
srom_1(87745) <= 8567963;
srom_1(87746) <= 7993569;
srom_1(87747) <= 7421028;
srom_1(87748) <= 6853023;
srom_1(87749) <= 6292220;
srom_1(87750) <= 5741247;
srom_1(87751) <= 5202689;
srom_1(87752) <= 4679070;
srom_1(87753) <= 4172847;
srom_1(87754) <= 3686393;
srom_1(87755) <= 3221989;
srom_1(87756) <= 2781814;
srom_1(87757) <= 2367930;
srom_1(87758) <= 1982279;
srom_1(87759) <= 1626670;
srom_1(87760) <= 1302770;
srom_1(87761) <= 1012098;
srom_1(87762) <= 756017;
srom_1(87763) <= 535728;
srom_1(87764) <= 352263;
srom_1(87765) <= 206484;
srom_1(87766) <= 99074;
srom_1(87767) <= 30536;
srom_1(87768) <= 1192;
srom_1(87769) <= 11179;
srom_1(87770) <= 60451;
srom_1(87771) <= 148776;
srom_1(87772) <= 275741;
srom_1(87773) <= 440750;
srom_1(87774) <= 643030;
srom_1(87775) <= 881630;
srom_1(87776) <= 1155434;
srom_1(87777) <= 1463157;
srom_1(87778) <= 1803355;
srom_1(87779) <= 2174434;
srom_1(87780) <= 2574653;
srom_1(87781) <= 3002136;
srom_1(87782) <= 3454877;
srom_1(87783) <= 3930755;
srom_1(87784) <= 4427537;
srom_1(87785) <= 4942894;
srom_1(87786) <= 5474409;
srom_1(87787) <= 6019590;
srom_1(87788) <= 6575880;
srom_1(87789) <= 7140671;
srom_1(87790) <= 7711313;
srom_1(87791) <= 8285131;
srom_1(87792) <= 8859435;
srom_1(87793) <= 9431531;
srom_1(87794) <= 9998736;
srom_1(87795) <= 10558391;
srom_1(87796) <= 11107871;
srom_1(87797) <= 11644599;
srom_1(87798) <= 12166059;
srom_1(87799) <= 12669805;
srom_1(87800) <= 13153475;
srom_1(87801) <= 13614801;
srom_1(87802) <= 14051620;
srom_1(87803) <= 14461882;
srom_1(87804) <= 14843665;
srom_1(87805) <= 15195178;
srom_1(87806) <= 15514773;
srom_1(87807) <= 15800951;
srom_1(87808) <= 16052369;
srom_1(87809) <= 16267850;
srom_1(87810) <= 16446382;
srom_1(87811) <= 16587129;
srom_1(87812) <= 16689429;
srom_1(87813) <= 16752805;
srom_1(87814) <= 16776958;
srom_1(87815) <= 16761774;
srom_1(87816) <= 16707327;
srom_1(87817) <= 16613870;
srom_1(87818) <= 16481841;
srom_1(87819) <= 16311861;
srom_1(87820) <= 16104726;
srom_1(87821) <= 15861408;
srom_1(87822) <= 15583047;
srom_1(87823) <= 15270948;
srom_1(87824) <= 14926576;
srom_1(87825) <= 14551546;
srom_1(87826) <= 14147615;
srom_1(87827) <= 13716678;
srom_1(87828) <= 13260756;
srom_1(87829) <= 12781987;
srom_1(87830) <= 12282616;
srom_1(87831) <= 11764984;
srom_1(87832) <= 11231519;
srom_1(87833) <= 10684723;
srom_1(87834) <= 10127160;
srom_1(87835) <= 9561444;
srom_1(87836) <= 8990228;
srom_1(87837) <= 8416191;
srom_1(87838) <= 7842025;
srom_1(87839) <= 7270422;
srom_1(87840) <= 6704062;
srom_1(87841) <= 6145602;
srom_1(87842) <= 5597660;
srom_1(87843) <= 5062805;
srom_1(87844) <= 4543547;
srom_1(87845) <= 4042319;
srom_1(87846) <= 3561473;
srom_1(87847) <= 3103262;
srom_1(87848) <= 2669837;
srom_1(87849) <= 2263228;
srom_1(87850) <= 1885344;
srom_1(87851) <= 1537956;
srom_1(87852) <= 1222693;
srom_1(87853) <= 941033;
srom_1(87854) <= 694297;
srom_1(87855) <= 483643;
srom_1(87856) <= 310058;
srom_1(87857) <= 174355;
srom_1(87858) <= 77173;
srom_1(87859) <= 18965;
srom_1(87860) <= 6;
srom_1(87861) <= 20384;
srom_1(87862) <= 80003;
srom_1(87863) <= 178584;
srom_1(87864) <= 315664;
srom_1(87865) <= 490602;
srom_1(87866) <= 702576;
srom_1(87867) <= 950592;
srom_1(87868) <= 1233488;
srom_1(87869) <= 1549936;
srom_1(87870) <= 1898454;
srom_1(87871) <= 2277406;
srom_1(87872) <= 2685015;
srom_1(87873) <= 3119371;
srom_1(87874) <= 3578435;
srom_1(87875) <= 4060057;
srom_1(87876) <= 4561976;
srom_1(87877) <= 5081840;
srom_1(87878) <= 5617211;
srom_1(87879) <= 6165577;
srom_1(87880) <= 6724368;
srom_1(87881) <= 7290963;
srom_1(87882) <= 7862706;
srom_1(87883) <= 8436914;
srom_1(87884) <= 9010896;
srom_1(87885) <= 9581960;
srom_1(87886) <= 10147428;
srom_1(87887) <= 10704648;
srom_1(87888) <= 11251007;
srom_1(87889) <= 11783944;
srom_1(87890) <= 12300958;
srom_1(87891) <= 12799627;
srom_1(87892) <= 13277610;
srom_1(87893) <= 13732668;
srom_1(87894) <= 14162665;
srom_1(87895) <= 14565586;
srom_1(87896) <= 14939540;
srom_1(87897) <= 15282775;
srom_1(87898) <= 15593681;
srom_1(87899) <= 15870800;
srom_1(87900) <= 16112832;
srom_1(87901) <= 16318643;
srom_1(87902) <= 16487267;
srom_1(87903) <= 16617914;
srom_1(87904) <= 16709971;
srom_1(87905) <= 16763006;
srom_1(87906) <= 16776770;
srom_1(87907) <= 16751200;
srom_1(87908) <= 16686414;
srom_1(87909) <= 16582717;
srom_1(87910) <= 16440595;
srom_1(87911) <= 16260715;
srom_1(87912) <= 16043919;
srom_1(87913) <= 15791226;
srom_1(87914) <= 15503818;
srom_1(87915) <= 15183046;
srom_1(87916) <= 14830411;
srom_1(87917) <= 14447569;
srom_1(87918) <= 14036314;
srom_1(87919) <= 13598575;
srom_1(87920) <= 13136405;
srom_1(87921) <= 12651971;
srom_1(87922) <= 12147545;
srom_1(87923) <= 11625491;
srom_1(87924) <= 11088259;
srom_1(87925) <= 10538367;
srom_1(87926) <= 9978394;
srom_1(87927) <= 9410966;
srom_1(87928) <= 8838744;
srom_1(87929) <= 8264411;
srom_1(87930) <= 7690660;
srom_1(87931) <= 7120182;
srom_1(87932) <= 6555652;
srom_1(87933) <= 5999718;
srom_1(87934) <= 5454986;
srom_1(87935) <= 4924011;
srom_1(87936) <= 4409282;
srom_1(87937) <= 3913214;
srom_1(87938) <= 3438133;
srom_1(87939) <= 2986266;
srom_1(87940) <= 2559732;
srom_1(87941) <= 2160532;
srom_1(87942) <= 1790538;
srom_1(87943) <= 1451484;
srom_1(87944) <= 1144961;
srom_1(87945) <= 872405;
srom_1(87946) <= 635096;
srom_1(87947) <= 434146;
srom_1(87948) <= 270497;
srom_1(87949) <= 144916;
srom_1(87950) <= 57993;
srom_1(87951) <= 10135;
srom_1(87952) <= 1567;
srom_1(87953) <= 32328;
srom_1(87954) <= 102275;
srom_1(87955) <= 211079;
srom_1(87956) <= 358230;
srom_1(87957) <= 543039;
srom_1(87958) <= 764638;
srom_1(87959) <= 1021989;
srom_1(87960) <= 1313884;
srom_1(87961) <= 1638955;
srom_1(87962) <= 1995677;
srom_1(87963) <= 2382378;
srom_1(87964) <= 2797245;
srom_1(87965) <= 3238331;
srom_1(87966) <= 3703568;
srom_1(87967) <= 4190776;
srom_1(87968) <= 4697668;
srom_1(87969) <= 5221869;
srom_1(87970) <= 5760919;
srom_1(87971) <= 6312292;
srom_1(87972) <= 6873401;
srom_1(87973) <= 7441615;
srom_1(87974) <= 8014270;
srom_1(87975) <= 8588681;
srom_1(87976) <= 9162153;
srom_1(87977) <= 9731998;
srom_1(87978) <= 10295543;
srom_1(87979) <= 10850146;
srom_1(87980) <= 11393206;
srom_1(87981) <= 11922177;
srom_1(87982) <= 12434577;
srom_1(87983) <= 12928004;
srom_1(87984) <= 13400145;
srom_1(87985) <= 13848785;
srom_1(87986) <= 14271820;
srom_1(87987) <= 14667266;
srom_1(87988) <= 15033270;
srom_1(87989) <= 15368115;
srom_1(87990) <= 15670230;
srom_1(87991) <= 15938200;
srom_1(87992) <= 16170767;
srom_1(87993) <= 16366840;
srom_1(87994) <= 16525501;
srom_1(87995) <= 16646005;
srom_1(87996) <= 16727788;
srom_1(87997) <= 16770465;
srom_1(87998) <= 16773836;
srom_1(87999) <= 16737887;
srom_1(88000) <= 16662785;
srom_1(88001) <= 16548882;
srom_1(88002) <= 16396713;
srom_1(88003) <= 16206991;
srom_1(88004) <= 15980606;
srom_1(88005) <= 15718620;
srom_1(88006) <= 15422261;
srom_1(88007) <= 15092918;
srom_1(88008) <= 14732137;
srom_1(88009) <= 14341609;
srom_1(88010) <= 13923165;
srom_1(88011) <= 13478767;
srom_1(88012) <= 13010500;
srom_1(88013) <= 12520560;
srom_1(88014) <= 12011243;
srom_1(88015) <= 11484939;
srom_1(88016) <= 10944114;
srom_1(88017) <= 10391306;
srom_1(88018) <= 9829107;
srom_1(88019) <= 9260153;
srom_1(88020) <= 8687111;
srom_1(88021) <= 8112670;
srom_1(88022) <= 7539523;
srom_1(88023) <= 6970358;
srom_1(88024) <= 6407843;
srom_1(88025) <= 5854617;
srom_1(88026) <= 5313273;
srom_1(88027) <= 4786351;
srom_1(88028) <= 4276321;
srom_1(88029) <= 3785575;
srom_1(88030) <= 3316414;
srom_1(88031) <= 2871038;
srom_1(88032) <= 2451536;
srom_1(88033) <= 2059875;
srom_1(88034) <= 1697892;
srom_1(88035) <= 1367283;
srom_1(88036) <= 1069600;
srom_1(88037) <= 806239;
srom_1(88038) <= 578434;
srom_1(88039) <= 387253;
srom_1(88040) <= 233593;
srom_1(88041) <= 118176;
srom_1(88042) <= 41540;
srom_1(88043) <= 4048;
srom_1(88044) <= 5873;
srom_1(88045) <= 47008;
srom_1(88046) <= 127259;
srom_1(88047) <= 246251;
srom_1(88048) <= 403425;
srom_1(88049) <= 598044;
srom_1(88050) <= 829196;
srom_1(88051) <= 1095797;
srom_1(88052) <= 1396596;
srom_1(88053) <= 1730183;
srom_1(88054) <= 2094994;
srom_1(88055) <= 2489317;
srom_1(88056) <= 2911305;
srom_1(88057) <= 3358977;
srom_1(88058) <= 3830235;
srom_1(88059) <= 4322869;
srom_1(88060) <= 4834568;
srom_1(88061) <= 5362934;
srom_1(88062) <= 5905488;
srom_1(88063) <= 6459686;
srom_1(88064) <= 7022929;
srom_1(88065) <= 7592577;
srom_1(88066) <= 8165957;
srom_1(88067) <= 8740382;
srom_1(88068) <= 9313157;
srom_1(88069) <= 9881596;
srom_1(88070) <= 10443035;
srom_1(88071) <= 10994839;
srom_1(88072) <= 11534422;
srom_1(88073) <= 12059253;
srom_1(88074) <= 12566871;
srom_1(88075) <= 13054896;
srom_1(88076) <= 13521039;
srom_1(88077) <= 13963114;
srom_1(88078) <= 14379048;
srom_1(88079) <= 14766892;
srom_1(88080) <= 15124825;
srom_1(88081) <= 15451170;
srom_1(88082) <= 15744396;
srom_1(88083) <= 16003128;
srom_1(88084) <= 16226153;
srom_1(88085) <= 16412425;
srom_1(88086) <= 16561071;
srom_1(88087) <= 16671393;
srom_1(88088) <= 16742874;
srom_1(88089) <= 16775180;
srom_1(88090) <= 16768157;
srom_1(88091) <= 16721841;
srom_1(88092) <= 16636446;
srom_1(88093) <= 16512375;
srom_1(88094) <= 16350209;
srom_1(88095) <= 16150708;
srom_1(88096) <= 15914808;
srom_1(88097) <= 15643615;
srom_1(88098) <= 15338401;
srom_1(88099) <= 15000596;
srom_1(88100) <= 14631786;
srom_1(88101) <= 14233700;
srom_1(88102) <= 13808203;
srom_1(88103) <= 13357293;
srom_1(88104) <= 12883082;
srom_1(88105) <= 12387796;
srom_1(88106) <= 11873755;
srom_1(88107) <= 11343372;
srom_1(88108) <= 10799133;
srom_1(88109) <= 10243590;
srom_1(88110) <= 9679349;
srom_1(88111) <= 9109054;
srom_1(88112) <= 8535382;
srom_1(88113) <= 7961021;
srom_1(88114) <= 7388665;
srom_1(88115) <= 6820998;
srom_1(88116) <= 6260682;
srom_1(88117) <= 5710345;
srom_1(88118) <= 5172567;
srom_1(88119) <= 4649870;
srom_1(88120) <= 4144705;
srom_1(88121) <= 3659442;
srom_1(88122) <= 3196355;
srom_1(88123) <= 2757616;
srom_1(88124) <= 2345284;
srom_1(88125) <= 1961290;
srom_1(88126) <= 1607436;
srom_1(88127) <= 1285381;
srom_1(88128) <= 996636;
srom_1(88129) <= 742555;
srom_1(88130) <= 524328;
srom_1(88131) <= 342980;
srom_1(88132) <= 199360;
srom_1(88133) <= 94143;
srom_1(88134) <= 27821;
srom_1(88135) <= 706;
srom_1(88136) <= 12924;
srom_1(88137) <= 64419;
srom_1(88138) <= 154949;
srom_1(88139) <= 284089;
srom_1(88140) <= 451234;
srom_1(88141) <= 655601;
srom_1(88142) <= 896230;
srom_1(88143) <= 1171993;
srom_1(88144) <= 1481598;
srom_1(88145) <= 1823591;
srom_1(88146) <= 2196371;
srom_1(88147) <= 2598188;
srom_1(88148) <= 3027158;
srom_1(88149) <= 3481270;
srom_1(88150) <= 3958394;
srom_1(88151) <= 4456293;
srom_1(88152) <= 4972632;
srom_1(88153) <= 5504990;
srom_1(88154) <= 6050869;
srom_1(88155) <= 6607712;
srom_1(88156) <= 7172905;
srom_1(88157) <= 7743799;
srom_1(88158) <= 8317718;
srom_1(88159) <= 8891968;
srom_1(88160) <= 9463858;
srom_1(88161) <= 10030706;
srom_1(88162) <= 10589853;
srom_1(88163) <= 11138678;
srom_1(88164) <= 11674607;
srom_1(88165) <= 12195127;
srom_1(88166) <= 12697797;
srom_1(88167) <= 13180259;
srom_1(88168) <= 13640252;
srom_1(88169) <= 14075618;
srom_1(88170) <= 14484316;
srom_1(88171) <= 14864429;
srom_1(88172) <= 15214174;
srom_1(88173) <= 15531912;
srom_1(88174) <= 15816153;
srom_1(88175) <= 16065563;
srom_1(88176) <= 16278973;
srom_1(88177) <= 16455383;
srom_1(88178) <= 16593965;
srom_1(88179) <= 16694069;
srom_1(88180) <= 16755226;
srom_1(88181) <= 16777149;
srom_1(88182) <= 16759735;
srom_1(88183) <= 16703066;
srom_1(88184) <= 16607408;
srom_1(88185) <= 16473209;
srom_1(88186) <= 16301098;
srom_1(88187) <= 16091884;
srom_1(88188) <= 15846545;
srom_1(88189) <= 15566234;
srom_1(88190) <= 15252265;
srom_1(88191) <= 14906109;
srom_1(88192) <= 14529391;
srom_1(88193) <= 14123877;
srom_1(88194) <= 13691467;
srom_1(88195) <= 13234191;
srom_1(88196) <= 12754193;
srom_1(88197) <= 12253722;
srom_1(88198) <= 11735127;
srom_1(88199) <= 11200839;
srom_1(88200) <= 10653363;
srom_1(88201) <= 10095267;
srom_1(88202) <= 9529168;
srom_1(88203) <= 8957720;
srom_1(88204) <= 8383604;
srom_1(88205) <= 7809511;
srom_1(88206) <= 7238133;
srom_1(88207) <= 6672151;
srom_1(88208) <= 6114218;
srom_1(88209) <= 5566950;
srom_1(88210) <= 5032913;
srom_1(88211) <= 4514613;
srom_1(88212) <= 4014479;
srom_1(88213) <= 3534857;
srom_1(88214) <= 3077996;
srom_1(88215) <= 2646039;
srom_1(88216) <= 2241010;
srom_1(88217) <= 1864809;
srom_1(88218) <= 1519201;
srom_1(88219) <= 1205805;
srom_1(88220) <= 926092;
srom_1(88221) <= 681374;
srom_1(88222) <= 472797;
srom_1(88223) <= 301341;
srom_1(88224) <= 167808;
srom_1(88225) <= 72825;
srom_1(88226) <= 16838;
srom_1(88227) <= 109;
srom_1(88228) <= 22717;
srom_1(88229) <= 84555;
srom_1(88230) <= 185334;
srom_1(88231) <= 324581;
srom_1(88232) <= 501642;
srom_1(88233) <= 715689;
srom_1(88234) <= 965716;
srom_1(88235) <= 1250552;
srom_1(88236) <= 1568860;
srom_1(88237) <= 1919149;
srom_1(88238) <= 2299775;
srom_1(88239) <= 2708954;
srom_1(88240) <= 3144767;
srom_1(88241) <= 3605170;
srom_1(88242) <= 4088004;
srom_1(88243) <= 4591005;
srom_1(88244) <= 5111814;
srom_1(88245) <= 5647989;
srom_1(88246) <= 6197016;
srom_1(88247) <= 6756321;
srom_1(88248) <= 7323279;
srom_1(88249) <= 7895233;
srom_1(88250) <= 8469501;
srom_1(88251) <= 9043389;
srom_1(88252) <= 9614207;
srom_1(88253) <= 10179278;
srom_1(88254) <= 10735951;
srom_1(88255) <= 11281617;
srom_1(88256) <= 11813717;
srom_1(88257) <= 12329755;
srom_1(88258) <= 12827312;
srom_1(88259) <= 13304054;
srom_1(88260) <= 13757746;
srom_1(88261) <= 14186261;
srom_1(88262) <= 14587588;
srom_1(88263) <= 14959846;
srom_1(88264) <= 15301289;
srom_1(88265) <= 15610316;
srom_1(88266) <= 15885478;
srom_1(88267) <= 16125485;
srom_1(88268) <= 16329210;
srom_1(88269) <= 16495700;
srom_1(88270) <= 16624173;
srom_1(88271) <= 16714026;
srom_1(88272) <= 16764838;
srom_1(88273) <= 16776372;
srom_1(88274) <= 16748572;
srom_1(88275) <= 16681570;
srom_1(88276) <= 16575679;
srom_1(88277) <= 16431396;
srom_1(88278) <= 16249397;
srom_1(88279) <= 16030537;
srom_1(88280) <= 15775841;
srom_1(88281) <= 15486504;
srom_1(88282) <= 15163882;
srom_1(88283) <= 14809489;
srom_1(88284) <= 14424986;
srom_1(88285) <= 14012176;
srom_1(88286) <= 13572996;
srom_1(88287) <= 13109504;
srom_1(88288) <= 12623874;
srom_1(88289) <= 12118383;
srom_1(88290) <= 11595403;
srom_1(88291) <= 11057384;
srom_1(88292) <= 10506851;
srom_1(88293) <= 9946385;
srom_1(88294) <= 9378613;
srom_1(88295) <= 8806199;
srom_1(88296) <= 8231827;
srom_1(88297) <= 7658190;
srom_1(88298) <= 7087979;
srom_1(88299) <= 6523866;
srom_1(88300) <= 5968498;
srom_1(88301) <= 5424478;
srom_1(88302) <= 4894359;
srom_1(88303) <= 4380625;
srom_1(88304) <= 3885685;
srom_1(88305) <= 3411862;
srom_1(88306) <= 2961376;
srom_1(88307) <= 2536341;
srom_1(88308) <= 2138748;
srom_1(88309) <= 1770464;
srom_1(88310) <= 1433214;
srom_1(88311) <= 1128580;
srom_1(88312) <= 857991;
srom_1(88313) <= 622716;
srom_1(88314) <= 423858;
srom_1(88315) <= 262349;
srom_1(88316) <= 138947;
srom_1(88317) <= 54231;
srom_1(88318) <= 8597;
srom_1(88319) <= 2260;
srom_1(88320) <= 35249;
srom_1(88321) <= 107410;
srom_1(88322) <= 218405;
srom_1(88323) <= 367712;
srom_1(88324) <= 554632;
srom_1(88325) <= 778289;
srom_1(88326) <= 1037633;
srom_1(88327) <= 1331448;
srom_1(88328) <= 1658356;
srom_1(88329) <= 2016825;
srom_1(88330) <= 2405173;
srom_1(88331) <= 2821580;
srom_1(88332) <= 3264092;
srom_1(88333) <= 3730635;
srom_1(88334) <= 4219021;
srom_1(88335) <= 4726960;
srom_1(88336) <= 5252069;
srom_1(88337) <= 5791887;
srom_1(88338) <= 6343881;
srom_1(88339) <= 6905464;
srom_1(88340) <= 7474002;
srom_1(88341) <= 8046828;
srom_1(88342) <= 8621258;
srom_1(88343) <= 9194596;
srom_1(88344) <= 9764155;
srom_1(88345) <= 10327263;
srom_1(88346) <= 10881281;
srom_1(88347) <= 11423609;
srom_1(88348) <= 11951706;
srom_1(88349) <= 12463093;
srom_1(88350) <= 12955374;
srom_1(88351) <= 13426240;
srom_1(88352) <= 13873483;
srom_1(88353) <= 14295005;
srom_1(88354) <= 14688830;
srom_1(88355) <= 15053111;
srom_1(88356) <= 15386140;
srom_1(88357) <= 15686355;
srom_1(88358) <= 15952349;
srom_1(88359) <= 16182873;
srom_1(88360) <= 16376848;
srom_1(88361) <= 16533363;
srom_1(88362) <= 16651684;
srom_1(88363) <= 16731257;
srom_1(88364) <= 16771708;
srom_1(88365) <= 16772848;
srom_1(88366) <= 16734672;
srom_1(88367) <= 16657358;
srom_1(88368) <= 16541269;
srom_1(88369) <= 16386949;
srom_1(88370) <= 16195123;
srom_1(88371) <= 15966689;
srom_1(88372) <= 15702718;
srom_1(88373) <= 15404450;
srom_1(88374) <= 15073281;
srom_1(88375) <= 14710766;
srom_1(88376) <= 14318604;
srom_1(88377) <= 13898634;
srom_1(88378) <= 13452826;
srom_1(88379) <= 12983270;
srom_1(88380) <= 12492168;
srom_1(88381) <= 11981823;
srom_1(88382) <= 11454629;
srom_1(88383) <= 10913056;
srom_1(88384) <= 10359646;
srom_1(88385) <= 9796992;
srom_1(88386) <= 9227735;
srom_1(88387) <= 8654542;
srom_1(88388) <= 8080102;
srom_1(88389) <= 7507109;
srom_1(88390) <= 6938250;
srom_1(88391) <= 6376192;
srom_1(88392) <= 5823570;
srom_1(88393) <= 5282977;
srom_1(88394) <= 4756948;
srom_1(88395) <= 4247948;
srom_1(88396) <= 3758366;
srom_1(88397) <= 3290496;
srom_1(88398) <= 2846533;
srom_1(88399) <= 2428559;
srom_1(88400) <= 2038533;
srom_1(88401) <= 1678285;
srom_1(88402) <= 1349505;
srom_1(88403) <= 1053732;
srom_1(88404) <= 792356;
srom_1(88405) <= 566601;
srom_1(88406) <= 377526;
srom_1(88407) <= 226018;
srom_1(88408) <= 112787;
srom_1(88409) <= 38364;
srom_1(88410) <= 3099;
srom_1(88411) <= 7156;
srom_1(88412) <= 50516;
srom_1(88413) <= 132976;
srom_1(88414) <= 254151;
srom_1(88415) <= 413470;
srom_1(88416) <= 610187;
srom_1(88417) <= 843380;
srom_1(88418) <= 1111956;
srom_1(88419) <= 1414654;
srom_1(88420) <= 1750055;
srom_1(88421) <= 2116587;
srom_1(88422) <= 2512530;
srom_1(88423) <= 2936028;
srom_1(88424) <= 3385096;
srom_1(88425) <= 3857626;
srom_1(88426) <= 4351404;
srom_1(88427) <= 4864114;
srom_1(88428) <= 5393351;
srom_1(88429) <= 5936634;
srom_1(88430) <= 6491415;
srom_1(88431) <= 7055093;
srom_1(88432) <= 7625024;
srom_1(88433) <= 8198535;
srom_1(88434) <= 8772938;
srom_1(88435) <= 9345539;
srom_1(88436) <= 9913653;
srom_1(88437) <= 10474614;
srom_1(88438) <= 11025794;
srom_1(88439) <= 11564608;
srom_1(88440) <= 12088527;
srom_1(88441) <= 12595097;
srom_1(88442) <= 13081941;
srom_1(88443) <= 13546776;
srom_1(88444) <= 13987423;
srom_1(88445) <= 14401816;
srom_1(88446) <= 14788010;
srom_1(88447) <= 15144195;
srom_1(88448) <= 15468701;
srom_1(88449) <= 15760005;
srom_1(88450) <= 16016743;
srom_1(88451) <= 16237710;
srom_1(88452) <= 16421870;
srom_1(88453) <= 16568359;
srom_1(88454) <= 16676490;
srom_1(88455) <= 16745757;
srom_1(88456) <= 16775834;
srom_1(88457) <= 16766580;
srom_1(88458) <= 16718040;
srom_1(88459) <= 16630439;
srom_1(88460) <= 16504190;
srom_1(88461) <= 16339884;
srom_1(88462) <= 16138292;
srom_1(88463) <= 15900359;
srom_1(88464) <= 15627201;
srom_1(88465) <= 15320098;
srom_1(88466) <= 14980492;
srom_1(88467) <= 14609973;
srom_1(88468) <= 14210281;
srom_1(88469) <= 13783289;
srom_1(88470) <= 13330999;
srom_1(88471) <= 12855533;
srom_1(88472) <= 12359119;
srom_1(88473) <= 11844087;
srom_1(88474) <= 11312851;
srom_1(88475) <= 10767902;
srom_1(88476) <= 10211795;
srom_1(88477) <= 9647139;
srom_1(88478) <= 9076581;
srom_1(88479) <= 8502798;
srom_1(88480) <= 7928478;
srom_1(88481) <= 7356317;
srom_1(88482) <= 6788996;
srom_1(88483) <= 6229176;
srom_1(88484) <= 5679483;
srom_1(88485) <= 5142493;
srom_1(88486) <= 4620726;
srom_1(88487) <= 4116628;
srom_1(88488) <= 3632562;
srom_1(88489) <= 3170799;
srom_1(88490) <= 2733504;
srom_1(88491) <= 2322728;
srom_1(88492) <= 1940397;
srom_1(88493) <= 1588304;
srom_1(88494) <= 1268100;
srom_1(88495) <= 981286;
srom_1(88496) <= 729208;
srom_1(88497) <= 513047;
srom_1(88498) <= 333817;
srom_1(88499) <= 192360;
srom_1(88500) <= 89337;
srom_1(88501) <= 25232;
srom_1(88502) <= 346;
srom_1(88503) <= 14795;
srom_1(88504) <= 68513;
srom_1(88505) <= 161246;
srom_1(88506) <= 292559;
srom_1(88507) <= 461838;
srom_1(88508) <= 668289;
srom_1(88509) <= 910942;
srom_1(88510) <= 1188661;
srom_1(88511) <= 1500143;
srom_1(88512) <= 1843927;
srom_1(88513) <= 2218402;
srom_1(88514) <= 2621811;
srom_1(88515) <= 3052262;
srom_1(88516) <= 3507737;
srom_1(88517) <= 3986100;
srom_1(88518) <= 4485108;
srom_1(88519) <= 5002421;
srom_1(88520) <= 5535613;
srom_1(88521) <= 6082184;
srom_1(88522) <= 6639570;
srom_1(88523) <= 7205158;
srom_1(88524) <= 7776296;
srom_1(88525) <= 8350305;
srom_1(88526) <= 8924493;
srom_1(88527) <= 9496169;
srom_1(88528) <= 10062651;
srom_1(88529) <= 10621283;
srom_1(88530) <= 11169444;
srom_1(88531) <= 11704566;
srom_1(88532) <= 12224138;
srom_1(88533) <= 12725724;
srom_1(88534) <= 13206971;
srom_1(88535) <= 13665624;
srom_1(88536) <= 14099531;
srom_1(88537) <= 14506657;
srom_1(88538) <= 14885094;
srom_1(88539) <= 15233067;
srom_1(88540) <= 15548943;
srom_1(88541) <= 15831242;
srom_1(88542) <= 16078640;
srom_1(88543) <= 16289977;
srom_1(88544) <= 16464262;
srom_1(88545) <= 16600677;
srom_1(88546) <= 16698583;
srom_1(88547) <= 16757521;
srom_1(88548) <= 16777213;
srom_1(88549) <= 16757569;
srom_1(88550) <= 16698680;
srom_1(88551) <= 16600822;
srom_1(88552) <= 16464454;
srom_1(88553) <= 16290216;
srom_1(88554) <= 16078925;
srom_1(88555) <= 15831570;
srom_1(88556) <= 15549314;
srom_1(88557) <= 15233478;
srom_1(88558) <= 14885544;
srom_1(88559) <= 14507144;
srom_1(88560) <= 14100052;
srom_1(88561) <= 13666177;
srom_1(88562) <= 13207554;
srom_1(88563) <= 12726333;
srom_1(88564) <= 12224771;
srom_1(88565) <= 11705219;
srom_1(88566) <= 11170115;
srom_1(88567) <= 10621968;
srom_1(88568) <= 10063348;
srom_1(88569) <= 9496874;
srom_1(88570) <= 8925203;
srom_1(88571) <= 8351016;
srom_1(88572) <= 7777005;
srom_1(88573) <= 7205862;
srom_1(88574) <= 6640266;
srom_1(88575) <= 6082868;
srom_1(88576) <= 5536282;
srom_1(88577) <= 5003072;
srom_1(88578) <= 4485738;
srom_1(88579) <= 3986706;
srom_1(88580) <= 3508315;
srom_1(88581) <= 3052811;
srom_1(88582) <= 2622327;
srom_1(88583) <= 2218884;
srom_1(88584) <= 1844372;
srom_1(88585) <= 1500549;
srom_1(88586) <= 1189026;
srom_1(88587) <= 911265;
srom_1(88588) <= 668567;
srom_1(88589) <= 462071;
srom_1(88590) <= 292746;
srom_1(88591) <= 161384;
srom_1(88592) <= 68603;
srom_1(88593) <= 14838;
srom_1(88594) <= 340;
srom_1(88595) <= 25177;
srom_1(88596) <= 89233;
srom_1(88597) <= 192208;
srom_1(88598) <= 333619;
srom_1(88599) <= 512802;
srom_1(88600) <= 728918;
srom_1(88601) <= 980952;
srom_1(88602) <= 1267724;
srom_1(88603) <= 1587888;
srom_1(88604) <= 1939942;
srom_1(88605) <= 2322237;
srom_1(88606) <= 2732979;
srom_1(88607) <= 3170242;
srom_1(88608) <= 3631976;
srom_1(88609) <= 4116016;
srom_1(88610) <= 4620091;
srom_1(88611) <= 5141837;
srom_1(88612) <= 5678810;
srom_1(88613) <= 6228489;
srom_1(88614) <= 6788298;
srom_1(88615) <= 7355611;
srom_1(88616) <= 7927768;
srom_1(88617) <= 8502086;
srom_1(88618) <= 9075873;
srom_1(88619) <= 9646436;
srom_1(88620) <= 10211101;
srom_1(88621) <= 10767220;
srom_1(88622) <= 11312184;
srom_1(88623) <= 11843439;
srom_1(88624) <= 12358493;
srom_1(88625) <= 12854931;
srom_1(88626) <= 13330424;
srom_1(88627) <= 13782744;
srom_1(88628) <= 14209769;
srom_1(88629) <= 14609496;
srom_1(88630) <= 14980052;
srom_1(88631) <= 15319698;
srom_1(88632) <= 15626841;
srom_1(88633) <= 15900043;
srom_1(88634) <= 16138020;
srom_1(88635) <= 16339658;
srom_1(88636) <= 16504010;
srom_1(88637) <= 16630307;
srom_1(88638) <= 16717955;
srom_1(88639) <= 16766545;
srom_1(88640) <= 16775847;
srom_1(88641) <= 16745818;
srom_1(88642) <= 16676600;
srom_1(88643) <= 16568517;
srom_1(88644) <= 16422075;
srom_1(88645) <= 16237961;
srom_1(88646) <= 16017039;
srom_1(88647) <= 15760345;
srom_1(88648) <= 15469082;
srom_1(88649) <= 15144616;
srom_1(88650) <= 14788469;
srom_1(88651) <= 14402311;
srom_1(88652) <= 13987953;
srom_1(88653) <= 13547337;
srom_1(88654) <= 13082531;
srom_1(88655) <= 12595712;
srom_1(88656) <= 12089166;
srom_1(88657) <= 11565266;
srom_1(88658) <= 11026470;
srom_1(88659) <= 10475303;
srom_1(88660) <= 9914352;
srom_1(88661) <= 9346246;
srom_1(88662) <= 8773649;
srom_1(88663) <= 8199246;
srom_1(88664) <= 7625732;
srom_1(88665) <= 7055795;
srom_1(88666) <= 6492108;
srom_1(88667) <= 5937314;
srom_1(88668) <= 5394015;
srom_1(88669) <= 4864759;
srom_1(88670) <= 4352027;
srom_1(88671) <= 3858225;
srom_1(88672) <= 3385666;
srom_1(88673) <= 2936569;
srom_1(88674) <= 2513038;
srom_1(88675) <= 2117059;
srom_1(88676) <= 1750490;
srom_1(88677) <= 1415049;
srom_1(88678) <= 1112310;
srom_1(88679) <= 843691;
srom_1(88680) <= 610454;
srom_1(88681) <= 413690;
srom_1(88682) <= 254324;
srom_1(88683) <= 133103;
srom_1(88684) <= 50594;
srom_1(88685) <= 7185;
srom_1(88686) <= 3079;
srom_1(88687) <= 38296;
srom_1(88688) <= 112671;
srom_1(88689) <= 225854;
srom_1(88690) <= 377315;
srom_1(88691) <= 566344;
srom_1(88692) <= 792054;
srom_1(88693) <= 1053387;
srom_1(88694) <= 1349118;
srom_1(88695) <= 1677859;
srom_1(88696) <= 2038069;
srom_1(88697) <= 2428058;
srom_1(88698) <= 2845999;
srom_1(88699) <= 3289931;
srom_1(88700) <= 3757773;
srom_1(88701) <= 4247330;
srom_1(88702) <= 4756307;
srom_1(88703) <= 5282317;
srom_1(88704) <= 5822893;
srom_1(88705) <= 6375501;
srom_1(88706) <= 6937549;
srom_1(88707) <= 7506402;
srom_1(88708) <= 8079392;
srom_1(88709) <= 8653831;
srom_1(88710) <= 9227027;
srom_1(88711) <= 9796291;
srom_1(88712) <= 10358954;
srom_1(88713) <= 10912378;
srom_1(88714) <= 11453967;
srom_1(88715) <= 11981181;
srom_1(88716) <= 12491548;
srom_1(88717) <= 12982675;
srom_1(88718) <= 13452259;
srom_1(88719) <= 13898098;
srom_1(88720) <= 14318101;
srom_1(88721) <= 14710299;
srom_1(88722) <= 15072851;
srom_1(88723) <= 15404060;
srom_1(88724) <= 15702370;
srom_1(88725) <= 15966384;
srom_1(88726) <= 16194862;
srom_1(88727) <= 16386735;
srom_1(88728) <= 16541101;
srom_1(88729) <= 16657238;
srom_1(88730) <= 16734600;
srom_1(88731) <= 16772826;
srom_1(88732) <= 16771734;
srom_1(88733) <= 16731331;
srom_1(88734) <= 16651807;
srom_1(88735) <= 16533533;
srom_1(88736) <= 16377065;
srom_1(88737) <= 16183136;
srom_1(88738) <= 15952656;
srom_1(88739) <= 15686706;
srom_1(88740) <= 15386532;
srom_1(88741) <= 15053543;
srom_1(88742) <= 14689300;
srom_1(88743) <= 14295510;
srom_1(88744) <= 13874021;
srom_1(88745) <= 13426809;
srom_1(88746) <= 12955971;
srom_1(88747) <= 12463715;
srom_1(88748) <= 11952349;
srom_1(88749) <= 11424272;
srom_1(88750) <= 10881960;
srom_1(88751) <= 10327955;
srom_1(88752) <= 9764857;
srom_1(88753) <= 9195304;
srom_1(88754) <= 8621969;
srom_1(88755) <= 8047539;
srom_1(88756) <= 7474709;
srom_1(88757) <= 6906164;
srom_1(88758) <= 6344571;
srom_1(88759) <= 5792563;
srom_1(88760) <= 5252729;
srom_1(88761) <= 4727600;
srom_1(88762) <= 4219638;
srom_1(88763) <= 3731227;
srom_1(88764) <= 3264655;
srom_1(88765) <= 2822112;
srom_1(88766) <= 2405672;
srom_1(88767) <= 2017287;
srom_1(88768) <= 1658781;
srom_1(88769) <= 1331832;
srom_1(88770) <= 1037975;
srom_1(88771) <= 778588;
srom_1(88772) <= 554887;
srom_1(88773) <= 367921;
srom_1(88774) <= 218566;
srom_1(88775) <= 107524;
srom_1(88776) <= 35314;
srom_1(88777) <= 2276;
srom_1(88778) <= 8565;
srom_1(88779) <= 54150;
srom_1(88780) <= 138818;
srom_1(88781) <= 262173;
srom_1(88782) <= 423635;
srom_1(88783) <= 622447;
srom_1(88784) <= 857678;
srom_1(88785) <= 1128224;
srom_1(88786) <= 1432816;
srom_1(88787) <= 1770027;
srom_1(88788) <= 2138274;
srom_1(88789) <= 2535831;
srom_1(88790) <= 2960834;
srom_1(88791) <= 3411290;
srom_1(88792) <= 3885085;
srom_1(88793) <= 4380000;
srom_1(88794) <= 4893712;
srom_1(88795) <= 5423813;
srom_1(88796) <= 5967817;
srom_1(88797) <= 6523173;
srom_1(88798) <= 7087276;
srom_1(88799) <= 7657482;
srom_1(88800) <= 8231116;
srom_1(88801) <= 8805489;
srom_1(88802) <= 9377907;
srom_1(88803) <= 9945686;
srom_1(88804) <= 10506163;
srom_1(88805) <= 11056710;
srom_1(88806) <= 11594745;
srom_1(88807) <= 12117746;
srom_1(88808) <= 12623260;
srom_1(88809) <= 13108916;
srom_1(88810) <= 13572436;
srom_1(88811) <= 14011648;
srom_1(88812) <= 14424492;
srom_1(88813) <= 14809031;
srom_1(88814) <= 15163463;
srom_1(88815) <= 15486125;
srom_1(88816) <= 15775504;
srom_1(88817) <= 16030244;
srom_1(88818) <= 16249149;
srom_1(88819) <= 16431194;
srom_1(88820) <= 16575524;
srom_1(88821) <= 16681462;
srom_1(88822) <= 16748513;
srom_1(88823) <= 16776362;
srom_1(88824) <= 16764877;
srom_1(88825) <= 16714113;
srom_1(88826) <= 16624308;
srom_1(88827) <= 16495883;
srom_1(88828) <= 16329440;
srom_1(88829) <= 16125759;
srom_1(88830) <= 15885797;
srom_1(88831) <= 15610678;
srom_1(88832) <= 15301692;
srom_1(88833) <= 14960288;
srom_1(88834) <= 14588067;
srom_1(88835) <= 14186775;
srom_1(88836) <= 13758293;
srom_1(88837) <= 13304631;
srom_1(88838) <= 12827916;
srom_1(88839) <= 12330383;
srom_1(88840) <= 11814366;
srom_1(88841) <= 11282285;
srom_1(88842) <= 10736634;
srom_1(88843) <= 10179973;
srom_1(88844) <= 9614911;
srom_1(88845) <= 9044098;
srom_1(88846) <= 8470212;
srom_1(88847) <= 7895943;
srom_1(88848) <= 7323984;
srom_1(88849) <= 6757018;
srom_1(88850) <= 6197703;
srom_1(88851) <= 5648662;
srom_1(88852) <= 5112469;
srom_1(88853) <= 4591639;
srom_1(88854) <= 4088614;
srom_1(88855) <= 3605754;
srom_1(88856) <= 3145322;
srom_1(88857) <= 2709478;
srom_1(88858) <= 2300265;
srom_1(88859) <= 1919602;
srom_1(88860) <= 1569275;
srom_1(88861) <= 1250925;
srom_1(88862) <= 966047;
srom_1(88863) <= 715976;
srom_1(88864) <= 501885;
srom_1(88865) <= 324777;
srom_1(88866) <= 185483;
srom_1(88867) <= 84656;
srom_1(88868) <= 22769;
srom_1(88869) <= 113;
srom_1(88870) <= 16793;
srom_1(88871) <= 72732;
srom_1(88872) <= 167666;
srom_1(88873) <= 301152;
srom_1(88874) <= 472562;
srom_1(88875) <= 681093;
srom_1(88876) <= 925768;
srom_1(88877) <= 1205438;
srom_1(88878) <= 1518792;
srom_1(88879) <= 1864362;
srom_1(88880) <= 2240526;
srom_1(88881) <= 2645520;
srom_1(88882) <= 3077446;
srom_1(88883) <= 3534277;
srom_1(88884) <= 4013873;
srom_1(88885) <= 4513982;
srom_1(88886) <= 5032262;
srom_1(88887) <= 5566280;
srom_1(88888) <= 6113533;
srom_1(88889) <= 6671455;
srom_1(88890) <= 7237429;
srom_1(88891) <= 7808801;
srom_1(88892) <= 8382892;
srom_1(88893) <= 8957010;
srom_1(88894) <= 9528463;
srom_1(88895) <= 10094570;
srom_1(88896) <= 10652678;
srom_1(88897) <= 11200169;
srom_1(88898) <= 11734475;
srom_1(88899) <= 12253091;
srom_1(88900) <= 12753585;
srom_1(88901) <= 13233611;
srom_1(88902) <= 13690916;
srom_1(88903) <= 14123358;
srom_1(88904) <= 14528907;
srom_1(88905) <= 14905662;
srom_1(88906) <= 15251856;
srom_1(88907) <= 15565866;
srom_1(88908) <= 15846220;
srom_1(88909) <= 16091602;
srom_1(88910) <= 16300862;
srom_1(88911) <= 16473019;
srom_1(88912) <= 16607266;
srom_1(88913) <= 16702972;
srom_1(88914) <= 16759689;
srom_1(88915) <= 16777152;
srom_1(88916) <= 16755277;
srom_1(88917) <= 16694169;
srom_1(88918) <= 16594113;
srom_1(88919) <= 16455578;
srom_1(88920) <= 16279215;
srom_1(88921) <= 16065850;
srom_1(88922) <= 15816483;
srom_1(88923) <= 15532285;
srom_1(88924) <= 15214588;
srom_1(88925) <= 14864881;
srom_1(88926) <= 14484804;
srom_1(88927) <= 14076141;
srom_1(88928) <= 13640807;
srom_1(88929) <= 13180843;
srom_1(88930) <= 12698407;
srom_1(88931) <= 12195761;
srom_1(88932) <= 11675262;
srom_1(88933) <= 11139350;
srom_1(88934) <= 10590540;
srom_1(88935) <= 10031403;
srom_1(88936) <= 9464563;
srom_1(88937) <= 8892678;
srom_1(88938) <= 8318429;
srom_1(88939) <= 7744509;
srom_1(88940) <= 7173609;
srom_1(88941) <= 6608407;
srom_1(88942) <= 6051552;
srom_1(88943) <= 5505657;
srom_1(88944) <= 4973282;
srom_1(88945) <= 4456921;
srom_1(88946) <= 3958998;
srom_1(88947) <= 3481847;
srom_1(88948) <= 3027705;
srom_1(88949) <= 2598703;
srom_1(88950) <= 2196851;
srom_1(88951) <= 1824034;
srom_1(88952) <= 1482001;
srom_1(88953) <= 1172356;
srom_1(88954) <= 896550;
srom_1(88955) <= 655876;
srom_1(88956) <= 451465;
srom_1(88957) <= 284273;
srom_1(88958) <= 155085;
srom_1(88959) <= 64507;
srom_1(88960) <= 12964;
srom_1(88961) <= 696;
srom_1(88962) <= 27763;
srom_1(88963) <= 94036;
srom_1(88964) <= 199206;
srom_1(88965) <= 342778;
srom_1(88966) <= 524081;
srom_1(88967) <= 742262;
srom_1(88968) <= 996300;
srom_1(88969) <= 1285003;
srom_1(88970) <= 1607017;
srom_1(88971) <= 1960833;
srom_1(88972) <= 2344790;
srom_1(88973) <= 2757089;
srom_1(88974) <= 3195796;
srom_1(88975) <= 3658854;
srom_1(88976) <= 4144092;
srom_1(88977) <= 4649233;
srom_1(88978) <= 5171910;
srom_1(88979) <= 5709671;
srom_1(88980) <= 6259994;
srom_1(88981) <= 6820299;
srom_1(88982) <= 7387958;
srom_1(88983) <= 7960310;
srom_1(88984) <= 8534670;
srom_1(88985) <= 9108346;
srom_1(88986) <= 9678646;
srom_1(88987) <= 10242897;
srom_1(88988) <= 10798452;
srom_1(88989) <= 11342707;
srom_1(88990) <= 11873109;
srom_1(88991) <= 12387170;
srom_1(88992) <= 12882482;
srom_1(88993) <= 13356720;
srom_1(88994) <= 13807660;
srom_1(88995) <= 14233189;
srom_1(88996) <= 14631311;
srom_1(88997) <= 15000159;
srom_1(88998) <= 15338002;
srom_1(88999) <= 15643258;
srom_1(89000) <= 15914494;
srom_1(89001) <= 16150438;
srom_1(89002) <= 16349985;
srom_1(89003) <= 16512198;
srom_1(89004) <= 16636317;
srom_1(89005) <= 16721759;
srom_1(89006) <= 16768124;
srom_1(89007) <= 16775195;
srom_1(89008) <= 16742939;
srom_1(89009) <= 16671505;
srom_1(89010) <= 16561231;
srom_1(89011) <= 16412632;
srom_1(89012) <= 16226406;
srom_1(89013) <= 16003426;
srom_1(89014) <= 15744738;
srom_1(89015) <= 15451553;
srom_1(89016) <= 15125249;
srom_1(89017) <= 14767354;
srom_1(89018) <= 14379546;
srom_1(89019) <= 13963645;
srom_1(89020) <= 13521601;
srom_1(89021) <= 13055487;
srom_1(89022) <= 12567488;
srom_1(89023) <= 12059892;
srom_1(89024) <= 11535081;
srom_1(89025) <= 10995515;
srom_1(89026) <= 10443724;
srom_1(89027) <= 9882296;
srom_1(89028) <= 9313864;
srom_1(89029) <= 8741093;
srom_1(89030) <= 8166668;
srom_1(89031) <= 7593285;
srom_1(89032) <= 7023631;
srom_1(89033) <= 6460378;
srom_1(89034) <= 5906167;
srom_1(89035) <= 5363597;
srom_1(89036) <= 4835213;
srom_1(89037) <= 4323491;
srom_1(89038) <= 3830832;
srom_1(89039) <= 3359546;
srom_1(89040) <= 2911844;
srom_1(89041) <= 2489823;
srom_1(89042) <= 2095464;
srom_1(89043) <= 1730616;
srom_1(89044) <= 1396989;
srom_1(89045) <= 1096149;
srom_1(89046) <= 829505;
srom_1(89047) <= 598308;
srom_1(89048) <= 403643;
srom_1(89049) <= 246422;
srom_1(89050) <= 127383;
srom_1(89051) <= 47083;
srom_1(89052) <= 5900;
srom_1(89053) <= 4026;
srom_1(89054) <= 41470;
srom_1(89055) <= 118057;
srom_1(89056) <= 233427;
srom_1(89057) <= 387039;
srom_1(89058) <= 578174;
srom_1(89059) <= 805935;
srom_1(89060) <= 1069253;
srom_1(89061) <= 1366894;
srom_1(89062) <= 1697463;
srom_1(89063) <= 2059408;
srom_1(89064) <= 2451034;
srom_1(89065) <= 2870502;
srom_1(89066) <= 3315847;
srom_1(89067) <= 3784980;
srom_1(89068) <= 4275701;
srom_1(89069) <= 4785708;
srom_1(89070) <= 5312611;
srom_1(89071) <= 5853939;
srom_1(89072) <= 6407152;
srom_1(89073) <= 6969657;
srom_1(89074) <= 7538816;
srom_1(89075) <= 8111960;
srom_1(89076) <= 8686401;
srom_1(89077) <= 9259445;
srom_1(89078) <= 9828406;
srom_1(89079) <= 10390616;
srom_1(89080) <= 10943437;
srom_1(89081) <= 11484278;
srom_1(89082) <= 12010602;
srom_1(89083) <= 12519941;
srom_1(89084) <= 13009907;
srom_1(89085) <= 13478202;
srom_1(89086) <= 13922630;
srom_1(89087) <= 14341108;
srom_1(89088) <= 14731672;
srom_1(89089) <= 15092491;
srom_1(89090) <= 15421873;
srom_1(89091) <= 15718274;
srom_1(89092) <= 15980304;
srom_1(89093) <= 16206734;
srom_1(89094) <= 16396501;
srom_1(89095) <= 16548717;
srom_1(89096) <= 16662668;
srom_1(89097) <= 16737818;
srom_1(89098) <= 16773816;
srom_1(89099) <= 16770493;
srom_1(89100) <= 16727865;
srom_1(89101) <= 16646130;
srom_1(89102) <= 16525674;
srom_1(89103) <= 16367060;
srom_1(89104) <= 16171032;
srom_1(89105) <= 15938510;
srom_1(89106) <= 15670584;
srom_1(89107) <= 15368509;
srom_1(89108) <= 15033704;
srom_1(89109) <= 14667738;
srom_1(89110) <= 14272327;
srom_1(89111) <= 13849325;
srom_1(89112) <= 13400715;
srom_1(89113) <= 12928602;
srom_1(89114) <= 12435200;
srom_1(89115) <= 11922822;
srom_1(89116) <= 11393870;
srom_1(89117) <= 10850826;
srom_1(89118) <= 10296236;
srom_1(89119) <= 9732700;
srom_1(89120) <= 9162861;
srom_1(89121) <= 8589392;
srom_1(89122) <= 8014981;
srom_1(89123) <= 7442322;
srom_1(89124) <= 6874100;
srom_1(89125) <= 6312981;
srom_1(89126) <= 5761594;
srom_1(89127) <= 5222527;
srom_1(89128) <= 4698307;
srom_1(89129) <= 4191392;
srom_1(89130) <= 3704158;
srom_1(89131) <= 3238892;
srom_1(89132) <= 2797775;
srom_1(89133) <= 2382875;
srom_1(89134) <= 1996138;
srom_1(89135) <= 1639377;
srom_1(89136) <= 1314266;
srom_1(89137) <= 1022329;
srom_1(89138) <= 764935;
srom_1(89139) <= 543291;
srom_1(89140) <= 358436;
srom_1(89141) <= 211237;
srom_1(89142) <= 102385;
srom_1(89143) <= 32390;
srom_1(89144) <= 1580;
srom_1(89145) <= 10100;
srom_1(89146) <= 57910;
srom_1(89147) <= 144784;
srom_1(89148) <= 270317;
srom_1(89149) <= 433920;
srom_1(89150) <= 634825;
srom_1(89151) <= 872090;
srom_1(89152) <= 1144602;
srom_1(89153) <= 1451084;
srom_1(89154) <= 1790099;
srom_1(89155) <= 2160056;
srom_1(89156) <= 2559221;
srom_1(89157) <= 2985722;
srom_1(89158) <= 3437559;
srom_1(89159) <= 3912613;
srom_1(89160) <= 4408656;
srom_1(89161) <= 4923363;
srom_1(89162) <= 5454320;
srom_1(89163) <= 5999036;
srom_1(89164) <= 6554958;
srom_1(89165) <= 7119479;
srom_1(89166) <= 7689951;
srom_1(89167) <= 8263699;
srom_1(89168) <= 8838033;
srom_1(89169) <= 9410260;
srom_1(89170) <= 9977695;
srom_1(89171) <= 10537679;
srom_1(89172) <= 11087585;
srom_1(89173) <= 11624835;
srom_1(89174) <= 12146909;
srom_1(89175) <= 12651359;
srom_1(89176) <= 13135819;
srom_1(89177) <= 13598018;
srom_1(89178) <= 14035788;
srom_1(89179) <= 14447077;
srom_1(89180) <= 14829956;
srom_1(89181) <= 15182628;
srom_1(89182) <= 15503442;
srom_1(89183) <= 15790891;
srom_1(89184) <= 16043629;
srom_1(89185) <= 16260469;
srom_1(89186) <= 16440396;
srom_1(89187) <= 16582565;
srom_1(89188) <= 16686310;
srom_1(89189) <= 16751144;
srom_1(89190) <= 16776763;
srom_1(89191) <= 16763047;
srom_1(89192) <= 16710061;
srom_1(89193) <= 16618052;
srom_1(89194) <= 16487453;
srom_1(89195) <= 16318875;
srom_1(89196) <= 16113110;
srom_1(89197) <= 15871122;
srom_1(89198) <= 15594045;
srom_1(89199) <= 15283180;
srom_1(89200) <= 14939984;
srom_1(89201) <= 14566067;
srom_1(89202) <= 14163181;
srom_1(89203) <= 13733216;
srom_1(89204) <= 13278188;
srom_1(89205) <= 12800232;
srom_1(89206) <= 12301588;
srom_1(89207) <= 11784594;
srom_1(89208) <= 11251676;
srom_1(89209) <= 10705331;
srom_1(89210) <= 10148123;
srom_1(89211) <= 9582664;
srom_1(89212) <= 9011605;
srom_1(89213) <= 8437625;
srom_1(89214) <= 7863415;
srom_1(89215) <= 7291668;
srom_1(89216) <= 6725065;
srom_1(89217) <= 6166263;
srom_1(89218) <= 5617882;
srom_1(89219) <= 5082494;
srom_1(89220) <= 4562609;
srom_1(89221) <= 4060666;
srom_1(89222) <= 3579018;
srom_1(89223) <= 3119924;
srom_1(89224) <= 2685537;
srom_1(89225) <= 2277893;
srom_1(89226) <= 1898904;
srom_1(89227) <= 1550348;
srom_1(89228) <= 1233859;
srom_1(89229) <= 950921;
srom_1(89230) <= 702861;
srom_1(89231) <= 490841;
srom_1(89232) <= 315858;
srom_1(89233) <= 178730;
srom_1(89234) <= 80101;
srom_1(89235) <= 20433;
srom_1(89236) <= 7;
srom_1(89237) <= 18918;
srom_1(89238) <= 77077;
srom_1(89239) <= 174211;
srom_1(89240) <= 309866;
srom_1(89241) <= 483405;
srom_1(89242) <= 694014;
srom_1(89243) <= 940705;
srom_1(89244) <= 1222323;
srom_1(89245) <= 1537545;
srom_1(89246) <= 1884895;
srom_1(89247) <= 2262742;
srom_1(89248) <= 2669316;
srom_1(89249) <= 3102710;
srom_1(89250) <= 3560891;
srom_1(89251) <= 4041711;
srom_1(89252) <= 4542915;
srom_1(89253) <= 5062152;
srom_1(89254) <= 5596989;
srom_1(89255) <= 6144917;
srom_1(89256) <= 6703365;
srom_1(89257) <= 7269717;
srom_1(89258) <= 7841315;
srom_1(89259) <= 8415480;
srom_1(89260) <= 8989519;
srom_1(89261) <= 9560740;
srom_1(89262) <= 10126464;
srom_1(89263) <= 10684039;
srom_1(89264) <= 11230850;
srom_1(89265) <= 11764333;
srom_1(89266) <= 12281986;
srom_1(89267) <= 12781381;
srom_1(89268) <= 13260177;
srom_1(89269) <= 13716129;
srom_1(89270) <= 14147098;
srom_1(89271) <= 14551063;
srom_1(89272) <= 14926131;
srom_1(89273) <= 15270542;
srom_1(89274) <= 15582681;
srom_1(89275) <= 15861085;
srom_1(89276) <= 16104447;
srom_1(89277) <= 16311628;
srom_1(89278) <= 16481654;
srom_1(89279) <= 16613730;
srom_1(89280) <= 16707235;
srom_1(89281) <= 16761731;
srom_1(89282) <= 16776963;
srom_1(89283) <= 16752859;
srom_1(89284) <= 16689532;
srom_1(89285) <= 16587279;
srom_1(89286) <= 16446580;
srom_1(89287) <= 16268094;
srom_1(89288) <= 16052659;
srom_1(89289) <= 15801284;
srom_1(89290) <= 15515148;
srom_1(89291) <= 15195594;
srom_1(89292) <= 14844120;
srom_1(89293) <= 14462373;
srom_1(89294) <= 14052144;
srom_1(89295) <= 13615357;
srom_1(89296) <= 13154060;
srom_1(89297) <= 12670417;
srom_1(89298) <= 12166694;
srom_1(89299) <= 11645255;
srom_1(89300) <= 11108544;
srom_1(89301) <= 10559078;
srom_1(89302) <= 9999434;
srom_1(89303) <= 9432237;
srom_1(89304) <= 8860145;
srom_1(89305) <= 8285843;
srom_1(89306) <= 7712022;
srom_1(89307) <= 7141374;
srom_1(89308) <= 6576575;
srom_1(89309) <= 6020273;
srom_1(89310) <= 5475076;
srom_1(89311) <= 4943543;
srom_1(89312) <= 4428164;
srom_1(89313) <= 3931358;
srom_1(89314) <= 3455453;
srom_1(89315) <= 3002681;
srom_1(89316) <= 2575165;
srom_1(89317) <= 2174911;
srom_1(89318) <= 1803795;
srom_1(89319) <= 1463558;
srom_1(89320) <= 1155794;
srom_1(89321) <= 881948;
srom_1(89322) <= 643303;
srom_1(89323) <= 440978;
srom_1(89324) <= 275922;
srom_1(89325) <= 148910;
srom_1(89326) <= 60536;
srom_1(89327) <= 11216;
srom_1(89328) <= 1180;
srom_1(89329) <= 30475;
srom_1(89330) <= 98965;
srom_1(89331) <= 206327;
srom_1(89332) <= 352060;
srom_1(89333) <= 535478;
srom_1(89334) <= 755722;
srom_1(89335) <= 1011760;
srom_1(89336) <= 1302390;
srom_1(89337) <= 1626250;
srom_1(89338) <= 1981820;
srom_1(89339) <= 2367435;
srom_1(89340) <= 2781284;
srom_1(89341) <= 3221429;
srom_1(89342) <= 3685804;
srom_1(89343) <= 4172232;
srom_1(89344) <= 4678432;
srom_1(89345) <= 5202031;
srom_1(89346) <= 5740572;
srom_1(89347) <= 6291531;
srom_1(89348) <= 6852324;
srom_1(89349) <= 7420321;
srom_1(89350) <= 7992859;
srom_1(89351) <= 8567252;
srom_1(89352) <= 9140808;
srom_1(89353) <= 9710836;
srom_1(89354) <= 10274664;
srom_1(89355) <= 10829648;
srom_1(89356) <= 11373185;
srom_1(89357) <= 11902726;
srom_1(89358) <= 12415788;
srom_1(89359) <= 12909965;
srom_1(89360) <= 13382940;
srom_1(89361) <= 13832495;
srom_1(89362) <= 14256522;
srom_1(89363) <= 14653032;
srom_1(89364) <= 15020166;
srom_1(89365) <= 15356202;
srom_1(89366) <= 15659565;
srom_1(89367) <= 15928831;
srom_1(89368) <= 16162740;
srom_1(89369) <= 16360192;
srom_1(89370) <= 16520263;
srom_1(89371) <= 16642202;
srom_1(89372) <= 16725437;
srom_1(89373) <= 16769578;
srom_1(89374) <= 16774417;
srom_1(89375) <= 16739933;
srom_1(89376) <= 16666286;
srom_1(89377) <= 16553822;
srom_1(89378) <= 16403069;
srom_1(89379) <= 16214733;
srom_1(89380) <= 15989698;
srom_1(89381) <= 15729019;
srom_1(89382) <= 15433918;
srom_1(89383) <= 15105779;
srom_1(89384) <= 14746141;
srom_1(89385) <= 14356691;
srom_1(89386) <= 13939254;
srom_1(89387) <= 13495788;
srom_1(89388) <= 13028373;
srom_1(89389) <= 12539200;
srom_1(89390) <= 12030564;
srom_1(89391) <= 11504849;
srom_1(89392) <= 10964521;
srom_1(89393) <= 10412114;
srom_1(89394) <= 9850218;
srom_1(89395) <= 9281468;
srom_1(89396) <= 8708531;
srom_1(89397) <= 8134094;
srom_1(89398) <= 7560850;
srom_1(89399) <= 6991488;
srom_1(89400) <= 6428677;
srom_1(89401) <= 5875058;
srom_1(89402) <= 5333225;
srom_1(89403) <= 4805720;
srom_1(89404) <= 4295016;
srom_1(89405) <= 3803509;
srom_1(89406) <= 3333502;
srom_1(89407) <= 2887201;
srom_1(89408) <= 2466698;
srom_1(89409) <= 2073964;
srom_1(89410) <= 1710842;
srom_1(89411) <= 1379035;
srom_1(89412) <= 1080098;
srom_1(89413) <= 815432;
srom_1(89414) <= 586281;
srom_1(89415) <= 393716;
srom_1(89416) <= 238643;
srom_1(89417) <= 121788;
srom_1(89418) <= 43698;
srom_1(89419) <= 4741;
srom_1(89420) <= 5098;
srom_1(89421) <= 44769;
srom_1(89422) <= 123567;
srom_1(89423) <= 241122;
srom_1(89424) <= 396884;
srom_1(89425) <= 590122;
srom_1(89426) <= 819929;
srom_1(89427) <= 1085229;
srom_1(89428) <= 1384777;
srom_1(89429) <= 1717168;
srom_1(89430) <= 2080843;
srom_1(89431) <= 2474098;
srom_1(89432) <= 2895088;
srom_1(89433) <= 3341840;
srom_1(89434) <= 3812257;
srom_1(89435) <= 4304134;
srom_1(89436) <= 4815165;
srom_1(89437) <= 5342952;
srom_1(89438) <= 5885022;
srom_1(89439) <= 6438832;
srom_1(89440) <= 7001786;
srom_1(89441) <= 7571242;
srom_1(89442) <= 8144532;
srom_1(89443) <= 8718966;
srom_1(89444) <= 9291850;
srom_1(89445) <= 9860500;
srom_1(89446) <= 10422247;
srom_1(89447) <= 10974457;
srom_1(89448) <= 11514542;
srom_1(89449) <= 12039968;
srom_1(89450) <= 12548271;
srom_1(89451) <= 13037069;
srom_1(89452) <= 13504068;
srom_1(89453) <= 13947079;
srom_1(89454) <= 14364024;
srom_1(89455) <= 14752949;
srom_1(89456) <= 15112029;
srom_1(89457) <= 15439581;
srom_1(89458) <= 15734068;
srom_1(89459) <= 15994110;
srom_1(89460) <= 16218487;
srom_1(89461) <= 16406147;
srom_1(89462) <= 16556210;
srom_1(89463) <= 16667972;
srom_1(89464) <= 16740910;
srom_1(89465) <= 16774680;
srom_1(89466) <= 16769126;
srom_1(89467) <= 16724272;
srom_1(89468) <= 16640330;
srom_1(89469) <= 16517692;
srom_1(89470) <= 16356934;
srom_1(89471) <= 16158811;
srom_1(89472) <= 15924249;
srom_1(89473) <= 15654351;
srom_1(89474) <= 15350381;
srom_1(89475) <= 15013765;
srom_1(89476) <= 14646082;
srom_1(89477) <= 14249055;
srom_1(89478) <= 13824546;
srom_1(89479) <= 13374546;
srom_1(89480) <= 12901166;
srom_1(89481) <= 12406624;
srom_1(89482) <= 11893241;
srom_1(89483) <= 11363423;
srom_1(89484) <= 10819655;
srom_1(89485) <= 10264488;
srom_1(89486) <= 9700523;
srom_1(89487) <= 9130407;
srom_1(89488) <= 8556812;
srom_1(89489) <= 7982428;
srom_1(89490) <= 7409949;
srom_1(89491) <= 6842059;
srom_1(89492) <= 6281422;
srom_1(89493) <= 5730666;
srom_1(89494) <= 5192374;
srom_1(89495) <= 4669070;
srom_1(89496) <= 4163208;
srom_1(89497) <= 3677161;
srom_1(89498) <= 3213207;
srom_1(89499) <= 2773522;
srom_1(89500) <= 2360169;
srom_1(89501) <= 1975085;
srom_1(89502) <= 1620076;
srom_1(89503) <= 1296807;
srom_1(89504) <= 1006794;
srom_1(89505) <= 751396;
srom_1(89506) <= 531813;
srom_1(89507) <= 349072;
srom_1(89508) <= 204032;
srom_1(89509) <= 97372;
srom_1(89510) <= 29592;
srom_1(89511) <= 1011;
srom_1(89512) <= 11762;
srom_1(89513) <= 61795;
srom_1(89514) <= 150875;
srom_1(89515) <= 278585;
srom_1(89516) <= 444325;
srom_1(89517) <= 647319;
srom_1(89518) <= 886615;
srom_1(89519) <= 1161089;
srom_1(89520) <= 1469457;
srom_1(89521) <= 1810270;
srom_1(89522) <= 2181931;
srom_1(89523) <= 2582698;
srom_1(89524) <= 3010691;
srom_1(89525) <= 3463902;
srom_1(89526) <= 3940208;
srom_1(89527) <= 4437373;
srom_1(89528) <= 4953067;
srom_1(89529) <= 5484871;
srom_1(89530) <= 6030292;
srom_1(89531) <= 6586772;
srom_1(89532) <= 7151701;
srom_1(89533) <= 7722431;
srom_1(89534) <= 8296284;
srom_1(89535) <= 8870571;
srom_1(89536) <= 9442597;
srom_1(89537) <= 10009681;
srom_1(89538) <= 10569163;
srom_1(89539) <= 11118420;
srom_1(89540) <= 11654876;
srom_1(89541) <= 12176015;
srom_1(89542) <= 12679393;
srom_1(89543) <= 13162651;
srom_1(89544) <= 13623521;
srom_1(89545) <= 14059843;
srom_1(89546) <= 14469571;
srom_1(89547) <= 14850783;
srom_1(89548) <= 15201692;
srom_1(89549) <= 15520651;
srom_1(89550) <= 15806167;
srom_1(89551) <= 16056898;
srom_1(89552) <= 16271671;
srom_1(89553) <= 16449477;
srom_1(89554) <= 16589482;
srom_1(89555) <= 16691031;
srom_1(89556) <= 16753648;
srom_1(89557) <= 16777037;
srom_1(89558) <= 16761091;
srom_1(89559) <= 16705883;
srom_1(89560) <= 16611672;
srom_1(89561) <= 16478901;
srom_1(89562) <= 16308191;
srom_1(89563) <= 16100344;
srom_1(89564) <= 15856333;
srom_1(89565) <= 15577305;
srom_1(89566) <= 15264565;
srom_1(89567) <= 14919582;
srom_1(89568) <= 14543973;
srom_1(89569) <= 14139500;
srom_1(89570) <= 13708058;
srom_1(89571) <= 13251672;
srom_1(89572) <= 12772481;
srom_1(89573) <= 12272733;
srom_1(89574) <= 11754771;
srom_1(89575) <= 11221023;
srom_1(89576) <= 10673994;
srom_1(89577) <= 10116247;
srom_1(89578) <= 9550399;
srom_1(89579) <= 8979103;
srom_1(89580) <= 8405038;
srom_1(89581) <= 7830895;
srom_1(89582) <= 7259369;
srom_1(89583) <= 6693137;
srom_1(89584) <= 6134856;
srom_1(89585) <= 5587144;
srom_1(89586) <= 5052569;
srom_1(89587) <= 4533637;
srom_1(89588) <= 4032783;
srom_1(89589) <= 3552355;
srom_1(89590) <= 3094606;
srom_1(89591) <= 2661682;
srom_1(89592) <= 2255613;
srom_1(89593) <= 1878304;
srom_1(89594) <= 1531525;
srom_1(89595) <= 1216900;
srom_1(89596) <= 935906;
srom_1(89597) <= 689861;
srom_1(89598) <= 479917;
srom_1(89599) <= 307060;
srom_1(89600) <= 172101;
srom_1(89601) <= 75671;
srom_1(89602) <= 18223;
srom_1(89603) <= 27;
srom_1(89604) <= 21168;
srom_1(89605) <= 81547;
srom_1(89606) <= 180880;
srom_1(89607) <= 318702;
srom_1(89608) <= 494367;
srom_1(89609) <= 707051;
srom_1(89610) <= 955756;
srom_1(89611) <= 1239316;
srom_1(89612) <= 1556402;
srom_1(89613) <= 1905526;
srom_1(89614) <= 2285052;
srom_1(89615) <= 2693199;
srom_1(89616) <= 3128054;
srom_1(89617) <= 3587578;
srom_1(89618) <= 4069615;
srom_1(89619) <= 4571905;
srom_1(89620) <= 5092094;
srom_1(89621) <= 5627740;
srom_1(89622) <= 6176334;
srom_1(89623) <= 6735301;
srom_1(89624) <= 7302022;
srom_1(89625) <= 7873838;
srom_1(89626) <= 8448068;
srom_1(89627) <= 9022018;
srom_1(89628) <= 9592999;
srom_1(89629) <= 10158332;
srom_1(89630) <= 10715366;
srom_1(89631) <= 11261489;
srom_1(89632) <= 11794140;
srom_1(89633) <= 12310821;
srom_1(89634) <= 12809110;
srom_1(89635) <= 13286670;
srom_1(89636) <= 13741260;
srom_1(89637) <= 14170751;
srom_1(89638) <= 14573127;
srom_1(89639) <= 14946501;
srom_1(89640) <= 15289124;
srom_1(89641) <= 15599387;
srom_1(89642) <= 15875837;
srom_1(89643) <= 16117176;
srom_1(89644) <= 16322273;
srom_1(89645) <= 16490167;
srom_1(89646) <= 16620070;
srom_1(89647) <= 16711373;
srom_1(89648) <= 16763647;
srom_1(89649) <= 16776648;
srom_1(89650) <= 16750314;
srom_1(89651) <= 16684770;
srom_1(89652) <= 16580322;
srom_1(89653) <= 16437460;
srom_1(89654) <= 16256855;
srom_1(89655) <= 16039352;
srom_1(89656) <= 15785973;
srom_1(89657) <= 15497904;
srom_1(89658) <= 15176498;
srom_1(89659) <= 14823261;
srom_1(89660) <= 14439850;
srom_1(89661) <= 14028062;
srom_1(89662) <= 13589829;
srom_1(89663) <= 13127206;
srom_1(89664) <= 12642362;
srom_1(89665) <= 12137570;
srom_1(89666) <= 11615198;
srom_1(89667) <= 11077696;
srom_1(89668) <= 10527584;
srom_1(89669) <= 9967441;
srom_1(89670) <= 9399894;
srom_1(89671) <= 8827606;
srom_1(89672) <= 8253258;
srom_1(89673) <= 7679545;
srom_1(89674) <= 7109158;
srom_1(89675) <= 6544770;
srom_1(89676) <= 5989028;
srom_1(89677) <= 5444539;
srom_1(89678) <= 4913856;
srom_1(89679) <= 4399467;
srom_1(89680) <= 3903784;
srom_1(89681) <= 3429133;
srom_1(89682) <= 2977738;
srom_1(89683) <= 2551716;
srom_1(89684) <= 2153066;
srom_1(89685) <= 1783656;
srom_1(89686) <= 1445219;
srom_1(89687) <= 1139342;
srom_1(89688) <= 867459;
srom_1(89689) <= 630846;
srom_1(89690) <= 430611;
srom_1(89691) <= 267694;
srom_1(89692) <= 142859;
srom_1(89693) <= 56691;
srom_1(89694) <= 9594;
srom_1(89695) <= 1790;
srom_1(89696) <= 33313;
srom_1(89697) <= 104018;
srom_1(89698) <= 213572;
srom_1(89699) <= 361462;
srom_1(89700) <= 546994;
srom_1(89701) <= 769297;
srom_1(89702) <= 1027330;
srom_1(89703) <= 1319883;
srom_1(89704) <= 1645584;
srom_1(89705) <= 2002905;
srom_1(89706) <= 2390170;
srom_1(89707) <= 2805564;
srom_1(89708) <= 3247139;
srom_1(89709) <= 3712825;
srom_1(89710) <= 4200436;
srom_1(89711) <= 4707687;
srom_1(89712) <= 5232200;
srom_1(89713) <= 5771514;
srom_1(89714) <= 6323100;
srom_1(89715) <= 6884372;
srom_1(89716) <= 7452698;
srom_1(89717) <= 8025413;
srom_1(89718) <= 8599831;
srom_1(89719) <= 9173259;
srom_1(89720) <= 9743007;
srom_1(89721) <= 10306403;
srom_1(89722) <= 10860807;
srom_1(89723) <= 11403617;
srom_1(89724) <= 11932290;
srom_1(89725) <= 12444344;
srom_1(89726) <= 12937380;
srom_1(89727) <= 13409085;
srom_1(89728) <= 13857247;
srom_1(89729) <= 14279765;
srom_1(89730) <= 14674658;
srom_1(89731) <= 15040072;
srom_1(89732) <= 15374296;
srom_1(89733) <= 15675762;
srom_1(89734) <= 15943055;
srom_1(89735) <= 16174924;
srom_1(89736) <= 16370279;
srom_1(89737) <= 16528206;
srom_1(89738) <= 16647963;
srom_1(89739) <= 16728989;
srom_1(89740) <= 16770905;
srom_1(89741) <= 16773512;
srom_1(89742) <= 16736801;
srom_1(89743) <= 16660941;
srom_1(89744) <= 16546290;
srom_1(89745) <= 16393385;
srom_1(89746) <= 16202942;
srom_1(89747) <= 15975856;
srom_1(89748) <= 15713190;
srom_1(89749) <= 15416177;
srom_1(89750) <= 15086209;
srom_1(89751) <= 14724833;
srom_1(89752) <= 14333745;
srom_1(89753) <= 13914778;
srom_1(89754) <= 13469897;
srom_1(89755) <= 13001188;
srom_1(89756) <= 12510849;
srom_1(89757) <= 12001180;
srom_1(89758) <= 11474570;
srom_1(89759) <= 10933488;
srom_1(89760) <= 10380473;
srom_1(89761) <= 9818118;
srom_1(89762) <= 9249059;
srom_1(89763) <= 8675964;
srom_1(89764) <= 8101523;
srom_1(89765) <= 7528428;
srom_1(89766) <= 6959366;
srom_1(89767) <= 6397006;
srom_1(89768) <= 5843986;
srom_1(89769) <= 5302899;
srom_1(89770) <= 4776281;
srom_1(89771) <= 4266603;
srom_1(89772) <= 3776254;
srom_1(89773) <= 3307534;
srom_1(89774) <= 2862641;
srom_1(89775) <= 2443662;
srom_1(89776) <= 2052560;
srom_1(89777) <= 1691170;
srom_1(89778) <= 1361186;
srom_1(89779) <= 1064157;
srom_1(89780) <= 801474;
srom_1(89781) <= 574371;
srom_1(89782) <= 383910;
srom_1(89783) <= 230987;
srom_1(89784) <= 116317;
srom_1(89785) <= 40439;
srom_1(89786) <= 3709;
srom_1(89787) <= 6298;
srom_1(89788) <= 48194;
srom_1(89789) <= 129202;
srom_1(89790) <= 248941;
srom_1(89791) <= 406850;
srom_1(89792) <= 602187;
srom_1(89793) <= 834038;
srom_1(89794) <= 1101315;
srom_1(89795) <= 1402765;
srom_1(89796) <= 1736973;
srom_1(89797) <= 2102374;
srom_1(89798) <= 2497252;
srom_1(89799) <= 2919758;
srom_1(89800) <= 3367908;
srom_1(89801) <= 3839602;
srom_1(89802) <= 4332629;
srom_1(89803) <= 4844675;
srom_1(89804) <= 5373339;
srom_1(89805) <= 5916144;
srom_1(89806) <= 6470542;
srom_1(89807) <= 7033935;
srom_1(89808) <= 7603681;
srom_1(89809) <= 8177107;
srom_1(89810) <= 8751526;
srom_1(89811) <= 9324242;
srom_1(89812) <= 9892571;
srom_1(89813) <= 10453847;
srom_1(89814) <= 11005438;
srom_1(89815) <= 11544759;
srom_1(89816) <= 12069279;
srom_1(89817) <= 12576539;
srom_1(89818) <= 13064160;
srom_1(89819) <= 13529857;
srom_1(89820) <= 13971444;
srom_1(89821) <= 14386851;
srom_1(89822) <= 14774130;
srom_1(89823) <= 15131466;
srom_1(89824) <= 15457182;
srom_1(89825) <= 15749751;
srom_1(89826) <= 16007801;
srom_1(89827) <= 16230122;
srom_1(89828) <= 16415671;
srom_1(89829) <= 16563579;
srom_1(89830) <= 16673152;
srom_1(89831) <= 16743875;
srom_1(89832) <= 16775418;
srom_1(89833) <= 16767632;
srom_1(89834) <= 16720554;
srom_1(89835) <= 16634404;
srom_1(89836) <= 16509588;
srom_1(89837) <= 16346689;
srom_1(89838) <= 16146472;
srom_1(89839) <= 15909875;
srom_1(89840) <= 15638009;
srom_1(89841) <= 15332148;
srom_1(89842) <= 14993726;
srom_1(89843) <= 14624331;
srom_1(89844) <= 14225694;
srom_1(89845) <= 13799685;
srom_1(89846) <= 13348302;
srom_1(89847) <= 12873661;
srom_1(89848) <= 12377988;
srom_1(89849) <= 11863607;
srom_1(89850) <= 11332931;
srom_1(89851) <= 10788448;
srom_1(89852) <= 10232711;
srom_1(89853) <= 9668327;
srom_1(89854) <= 9097941;
srom_1(89855) <= 8524229;
srom_1(89856) <= 7949882;
srom_1(89857) <= 7377591;
srom_1(89858) <= 6810042;
srom_1(89859) <= 6249895;
srom_1(89860) <= 5699777;
srom_1(89861) <= 5162268;
srom_1(89862) <= 4639889;
srom_1(89863) <= 4135088;
srom_1(89864) <= 3650234;
srom_1(89865) <= 3187599;
srom_1(89866) <= 2749354;
srom_1(89867) <= 2337553;
srom_1(89868) <= 1954128;
srom_1(89869) <= 1600876;
srom_1(89870) <= 1279454;
srom_1(89871) <= 991370;
srom_1(89872) <= 737973;
srom_1(89873) <= 520454;
srom_1(89874) <= 339830;
srom_1(89875) <= 196950;
srom_1(89876) <= 92484;
srom_1(89877) <= 26921;
srom_1(89878) <= 568;
srom_1(89879) <= 13550;
srom_1(89880) <= 65806;
srom_1(89881) <= 157090;
srom_1(89882) <= 286975;
srom_1(89883) <= 454850;
srom_1(89884) <= 659930;
srom_1(89885) <= 901253;
srom_1(89886) <= 1177686;
srom_1(89887) <= 1487933;
srom_1(89888) <= 1830541;
srom_1(89889) <= 2203901;
srom_1(89890) <= 2606263;
srom_1(89891) <= 3035741;
srom_1(89892) <= 3490321;
srom_1(89893) <= 3967870;
srom_1(89894) <= 4466149;
srom_1(89895) <= 4982822;
srom_1(89896) <= 5515466;
srom_1(89897) <= 6061583;
srom_1(89898) <= 6618613;
srom_1(89899) <= 7183942;
srom_1(89900) <= 7754921;
srom_1(89901) <= 8328871;
srom_1(89902) <= 8903101;
srom_1(89903) <= 9474919;
srom_1(89904) <= 10041642;
srom_1(89905) <= 10600614;
srom_1(89906) <= 11149213;
srom_1(89907) <= 11684867;
srom_1(89908) <= 12205063;
srom_1(89909) <= 12707363;
srom_1(89910) <= 13189410;
srom_1(89911) <= 13648945;
srom_1(89912) <= 14083812;
srom_1(89913) <= 14491973;
srom_1(89914) <= 14871513;
srom_1(89915) <= 15220652;
srom_1(89916) <= 15537753;
srom_1(89917) <= 15821330;
srom_1(89918) <= 16070052;
srom_1(89919) <= 16282753;
srom_1(89920) <= 16458436;
srom_1(89921) <= 16596276;
srom_1(89922) <= 16695628;
srom_1(89923) <= 16756025;
srom_1(89924) <= 16777185;
srom_1(89925) <= 16759008;
srom_1(89926) <= 16701579;
srom_1(89927) <= 16605168;
srom_1(89928) <= 16470226;
srom_1(89929) <= 16297387;
srom_1(89930) <= 16087461;
srom_1(89931) <= 15841433;
srom_1(89932) <= 15560455;
srom_1(89933) <= 15245846;
srom_1(89934) <= 14899082;
srom_1(89935) <= 14521787;
srom_1(89936) <= 14115732;
srom_1(89937) <= 13682820;
srom_1(89938) <= 13225082;
srom_1(89939) <= 12744665;
srom_1(89940) <= 12243820;
srom_1(89941) <= 11724896;
srom_1(89942) <= 11190328;
srom_1(89943) <= 10642621;
srom_1(89944) <= 10084345;
srom_1(89945) <= 9518116;
srom_1(89946) <= 8946591;
srom_1(89947) <= 8372450;
srom_1(89948) <= 7798384;
srom_1(89949) <= 7227086;
srom_1(89950) <= 6661235;
srom_1(89951) <= 6103484;
srom_1(89952) <= 5556448;
srom_1(89953) <= 5022694;
srom_1(89954) <= 4504723;
srom_1(89955) <= 4004966;
srom_1(89956) <= 3525765;
srom_1(89957) <= 3069367;
srom_1(89958) <= 2637913;
srom_1(89959) <= 2233426;
srom_1(89960) <= 1857803;
srom_1(89961) <= 1512805;
srom_1(89962) <= 1200050;
srom_1(89963) <= 921005;
srom_1(89964) <= 676977;
srom_1(89965) <= 469113;
srom_1(89966) <= 298385;
srom_1(89967) <= 165595;
srom_1(89968) <= 71366;
srom_1(89969) <= 16139;
srom_1(89970) <= 174;
srom_1(89971) <= 23545;
srom_1(89972) <= 86142;
srom_1(89973) <= 187673;
srom_1(89974) <= 327660;
srom_1(89975) <= 505449;
srom_1(89976) <= 720204;
srom_1(89977) <= 970918;
srom_1(89978) <= 1256417;
srom_1(89979) <= 1575361;
srom_1(89980) <= 1926255;
srom_1(89981) <= 2307453;
srom_1(89982) <= 2717167;
srom_1(89983) <= 3153477;
srom_1(89984) <= 3614337;
srom_1(89985) <= 4097584;
srom_1(89986) <= 4600953;
srom_1(89987) <= 5122085;
srom_1(89988) <= 5658533;
srom_1(89989) <= 6207785;
srom_1(89990) <= 6767262;
srom_1(89991) <= 7334343;
srom_1(89992) <= 7906368;
srom_1(89993) <= 8480654;
srom_1(89994) <= 9054508;
srom_1(89995) <= 9625240;
srom_1(89996) <= 10190173;
srom_1(89997) <= 10746657;
srom_1(89998) <= 11292084;
srom_1(89999) <= 11823896;
srom_1(90000) <= 12339598;
srom_1(90001) <= 12836773;
srom_1(90002) <= 13313088;
srom_1(90003) <= 13766311;
srom_1(90004) <= 14194317;
srom_1(90005) <= 14595097;
srom_1(90006) <= 14966773;
srom_1(90007) <= 15307601;
srom_1(90008) <= 15615984;
srom_1(90009) <= 15890476;
srom_1(90010) <= 16129788;
srom_1(90011) <= 16332800;
srom_1(90012) <= 16498558;
srom_1(90013) <= 16626286;
srom_1(90014) <= 16715385;
srom_1(90015) <= 16765436;
srom_1(90016) <= 16776206;
srom_1(90017) <= 16747644;
srom_1(90018) <= 16679883;
srom_1(90019) <= 16573241;
srom_1(90020) <= 16428219;
srom_1(90021) <= 16245496;
srom_1(90022) <= 16025930;
srom_1(90023) <= 15770550;
srom_1(90024) <= 15480553;
srom_1(90025) <= 15157300;
srom_1(90026) <= 14802305;
srom_1(90027) <= 14417235;
srom_1(90028) <= 14003895;
srom_1(90029) <= 13564222;
srom_1(90030) <= 13100280;
srom_1(90031) <= 12614242;
srom_1(90032) <= 12108389;
srom_1(90033) <= 11585093;
srom_1(90034) <= 11046808;
srom_1(90035) <= 10496057;
srom_1(90036) <= 9935424;
srom_1(90037) <= 9367537;
srom_1(90038) <= 8795059;
srom_1(90039) <= 8220676;
srom_1(90040) <= 7647080;
srom_1(90041) <= 7076961;
srom_1(90042) <= 6512993;
srom_1(90043) <= 5957820;
srom_1(90044) <= 5414047;
srom_1(90045) <= 4884222;
srom_1(90046) <= 4370830;
srom_1(90047) <= 3876279;
srom_1(90048) <= 3402888;
srom_1(90049) <= 2952876;
srom_1(90050) <= 2528355;
srom_1(90051) <= 2131314;
srom_1(90052) <= 1763616;
srom_1(90053) <= 1426985;
srom_1(90054) <= 1122999;
srom_1(90055) <= 853084;
srom_1(90056) <= 618506;
srom_1(90057) <= 420364;
srom_1(90058) <= 259589;
srom_1(90059) <= 136933;
srom_1(90060) <= 52972;
srom_1(90061) <= 8099;
srom_1(90062) <= 2526;
srom_1(90063) <= 36278;
srom_1(90064) <= 109197;
srom_1(90065) <= 220941;
srom_1(90066) <= 370985;
srom_1(90067) <= 558628;
srom_1(90068) <= 782987;
srom_1(90069) <= 1043012;
srom_1(90070) <= 1337483;
srom_1(90071) <= 1665020;
srom_1(90072) <= 2024085;
srom_1(90073) <= 2412996;
srom_1(90074) <= 2829928;
srom_1(90075) <= 3272927;
srom_1(90076) <= 3739916;
srom_1(90077) <= 4228703;
srom_1(90078) <= 4736998;
srom_1(90079) <= 5262416;
srom_1(90080) <= 5802495;
srom_1(90081) <= 6354700;
srom_1(90082) <= 6916443;
srom_1(90083) <= 7485090;
srom_1(90084) <= 8057973;
srom_1(90085) <= 8632407;
srom_1(90086) <= 9205698;
srom_1(90087) <= 9775157;
srom_1(90088) <= 10338114;
srom_1(90089) <= 10891929;
srom_1(90090) <= 11434005;
srom_1(90091) <= 11961800;
srom_1(90092) <= 12472839;
srom_1(90093) <= 12964726;
srom_1(90094) <= 13435154;
srom_1(90095) <= 13881917;
srom_1(90096) <= 14302920;
srom_1(90097) <= 14696189;
srom_1(90098) <= 15059879;
srom_1(90099) <= 15392285;
srom_1(90100) <= 15691849;
srom_1(90101) <= 15957165;
srom_1(90102) <= 16186990;
srom_1(90103) <= 16380245;
srom_1(90104) <= 16536025;
srom_1(90105) <= 16653599;
srom_1(90106) <= 16732416;
srom_1(90107) <= 16772105;
srom_1(90108) <= 16772481;
srom_1(90109) <= 16733543;
srom_1(90110) <= 16655472;
srom_1(90111) <= 16538635;
srom_1(90112) <= 16383580;
srom_1(90113) <= 16191033;
srom_1(90114) <= 15961899;
srom_1(90115) <= 15697250;
srom_1(90116) <= 15398329;
srom_1(90117) <= 15066537;
srom_1(90118) <= 14703429;
srom_1(90119) <= 14310710;
srom_1(90120) <= 13890219;
srom_1(90121) <= 13443930;
srom_1(90122) <= 12973934;
srom_1(90123) <= 12482437;
srom_1(90124) <= 11971742;
srom_1(90125) <= 11444244;
srom_1(90126) <= 10902417;
srom_1(90127) <= 10348803;
srom_1(90128) <= 9785996;
srom_1(90129) <= 9216636;
srom_1(90130) <= 8643394;
srom_1(90131) <= 8068956;
srom_1(90132) <= 7496018;
srom_1(90133) <= 6927265;
srom_1(90134) <= 6365365;
srom_1(90135) <= 5812953;
srom_1(90136) <= 5272619;
srom_1(90137) <= 4746897;
srom_1(90138) <= 4238252;
srom_1(90139) <= 3749069;
srom_1(90140) <= 3281643;
srom_1(90141) <= 2838165;
srom_1(90142) <= 2420715;
srom_1(90143) <= 2031251;
srom_1(90144) <= 1671598;
srom_1(90145) <= 1343444;
srom_1(90146) <= 1048327;
srom_1(90147) <= 787631;
srom_1(90148) <= 562578;
srom_1(90149) <= 374225;
srom_1(90150) <= 223454;
srom_1(90151) <= 110972;
srom_1(90152) <= 37306;
srom_1(90153) <= 2803;
srom_1(90154) <= 7624;
srom_1(90155) <= 51746;
srom_1(90156) <= 134962;
srom_1(90157) <= 256882;
srom_1(90158) <= 416935;
srom_1(90159) <= 614370;
srom_1(90160) <= 848261;
srom_1(90161) <= 1117511;
srom_1(90162) <= 1420858;
srom_1(90163) <= 1756879;
srom_1(90164) <= 2123999;
srom_1(90165) <= 2520495;
srom_1(90166) <= 2944509;
srom_1(90167) <= 3394052;
srom_1(90168) <= 3867017;
srom_1(90169) <= 4361185;
srom_1(90170) <= 4874238;
srom_1(90171) <= 5403772;
srom_1(90172) <= 5947303;
srom_1(90173) <= 6502281;
srom_1(90174) <= 7066106;
srom_1(90175) <= 7636132;
srom_1(90176) <= 8209686;
srom_1(90177) <= 8784080;
srom_1(90178) <= 9356619;
srom_1(90179) <= 9924619;
srom_1(90180) <= 10485416;
srom_1(90181) <= 11036380;
srom_1(90182) <= 11574928;
srom_1(90183) <= 12098534;
srom_1(90184) <= 12604743;
srom_1(90185) <= 13091182;
srom_1(90186) <= 13555568;
srom_1(90187) <= 13995724;
srom_1(90188) <= 14409587;
srom_1(90189) <= 14795215;
srom_1(90190) <= 15150801;
srom_1(90191) <= 15474676;
srom_1(90192) <= 15765323;
srom_1(90193) <= 16021377;
srom_1(90194) <= 16241639;
srom_1(90195) <= 16425075;
srom_1(90196) <= 16570825;
srom_1(90197) <= 16678206;
srom_1(90198) <= 16746714;
srom_1(90199) <= 16776029;
srom_1(90200) <= 16766012;
srom_1(90201) <= 16716710;
srom_1(90202) <= 16628355;
srom_1(90203) <= 16501361;
srom_1(90204) <= 16336323;
srom_1(90205) <= 16134016;
srom_1(90206) <= 15895388;
srom_1(90207) <= 15621558;
srom_1(90208) <= 15313810;
srom_1(90209) <= 14973588;
srom_1(90210) <= 14602486;
srom_1(90211) <= 14202245;
srom_1(90212) <= 13774743;
srom_1(90213) <= 13321982;
srom_1(90214) <= 12846088;
srom_1(90215) <= 12349291;
srom_1(90216) <= 11833921;
srom_1(90217) <= 11302394;
srom_1(90218) <= 10757204;
srom_1(90219) <= 10200906;
srom_1(90220) <= 9636111;
srom_1(90221) <= 9065465;
srom_1(90222) <= 8491645;
srom_1(90223) <= 7917342;
srom_1(90224) <= 7345249;
srom_1(90225) <= 6778048;
srom_1(90226) <= 6218400;
srom_1(90227) <= 5668929;
srom_1(90228) <= 5132211;
srom_1(90229) <= 4610764;
srom_1(90230) <= 4107032;
srom_1(90231) <= 3623378;
srom_1(90232) <= 3162070;
srom_1(90233) <= 2725271;
srom_1(90234) <= 2315029;
srom_1(90235) <= 1933269;
srom_1(90236) <= 1581779;
srom_1(90237) <= 1262209;
srom_1(90238) <= 976058;
srom_1(90239) <= 724666;
srom_1(90240) <= 509213;
srom_1(90241) <= 330709;
srom_1(90242) <= 189992;
srom_1(90243) <= 87721;
srom_1(90244) <= 24375;
srom_1(90245) <= 252;
srom_1(90246) <= 15465;
srom_1(90247) <= 69943;
srom_1(90248) <= 163429;
srom_1(90249) <= 295486;
srom_1(90250) <= 465495;
srom_1(90251) <= 672658;
srom_1(90252) <= 916004;
srom_1(90253) <= 1194391;
srom_1(90254) <= 1506514;
srom_1(90255) <= 1850910;
srom_1(90256) <= 2225964;
srom_1(90257) <= 2629916;
srom_1(90258) <= 3060872;
srom_1(90259) <= 3516813;
srom_1(90260) <= 3995598;
srom_1(90261) <= 4494984;
srom_1(90262) <= 5012629;
srom_1(90263) <= 5546105;
srom_1(90264) <= 6092910;
srom_1(90265) <= 6650480;
srom_1(90266) <= 7216201;
srom_1(90267) <= 7787420;
srom_1(90268) <= 8361458;
srom_1(90269) <= 8935624;
srom_1(90270) <= 9507224;
srom_1(90271) <= 10073579;
srom_1(90272) <= 10632032;
srom_1(90273) <= 11179965;
srom_1(90274) <= 11714808;
srom_1(90275) <= 12234054;
srom_1(90276) <= 12735267;
srom_1(90277) <= 13216097;
srom_1(90278) <= 13674290;
srom_1(90279) <= 14107696;
srom_1(90280) <= 14514283;
srom_1(90281) <= 14892145;
srom_1(90282) <= 15239509;
srom_1(90283) <= 15554747;
srom_1(90284) <= 15836381;
srom_1(90285) <= 16083090;
srom_1(90286) <= 16293716;
srom_1(90287) <= 16467273;
srom_1(90288) <= 16602946;
srom_1(90289) <= 16700099;
srom_1(90290) <= 16758277;
srom_1(90291) <= 16777207;
srom_1(90292) <= 16756799;
srom_1(90293) <= 16697150;
srom_1(90294) <= 16598540;
srom_1(90295) <= 16461430;
srom_1(90296) <= 16286464;
srom_1(90297) <= 16074462;
srom_1(90298) <= 15826419;
srom_1(90299) <= 15543497;
srom_1(90300) <= 15227024;
srom_1(90301) <= 14878483;
srom_1(90302) <= 14499508;
srom_1(90303) <= 14091878;
srom_1(90304) <= 13657503;
srom_1(90305) <= 13198420;
srom_1(90306) <= 12716782;
srom_1(90307) <= 12214848;
srom_1(90308) <= 11694972;
srom_1(90309) <= 11159590;
srom_1(90310) <= 10611215;
srom_1(90311) <= 10052417;
srom_1(90312) <= 9485817;
srom_1(90313) <= 8914072;
srom_1(90314) <= 8339862;
srom_1(90315) <= 7765882;
srom_1(90316) <= 7194821;
srom_1(90317) <= 6629358;
srom_1(90318) <= 6072146;
srom_1(90319) <= 5525795;
srom_1(90320) <= 4992870;
srom_1(90321) <= 4475868;
srom_1(90322) <= 3977215;
srom_1(90323) <= 3499248;
srom_1(90324) <= 3044209;
srom_1(90325) <= 2614231;
srom_1(90326) <= 2211332;
srom_1(90327) <= 1837400;
srom_1(90328) <= 1494189;
srom_1(90329) <= 1183308;
srom_1(90330) <= 906215;
srom_1(90331) <= 664210;
srom_1(90332) <= 458427;
srom_1(90333) <= 289832;
srom_1(90334) <= 159214;
srom_1(90335) <= 67187;
srom_1(90336) <= 14182;
srom_1(90337) <= 447;
srom_1(90338) <= 26048;
srom_1(90339) <= 90863;
srom_1(90340) <= 194589;
srom_1(90341) <= 336740;
srom_1(90342) <= 516649;
srom_1(90343) <= 733472;
srom_1(90344) <= 986193;
srom_1(90345) <= 1273626;
srom_1(90346) <= 1594424;
srom_1(90347) <= 1947081;
srom_1(90348) <= 2329946;
srom_1(90349) <= 2741222;
srom_1(90350) <= 3178980;
srom_1(90351) <= 3641168;
srom_1(90352) <= 4125618;
srom_1(90353) <= 4630059;
srom_1(90354) <= 5152125;
srom_1(90355) <= 5689368;
srom_1(90356) <= 6239268;
srom_1(90357) <= 6799248;
srom_1(90358) <= 7366681;
srom_1(90359) <= 7938905;
srom_1(90360) <= 8513239;
srom_1(90361) <= 9086988;
srom_1(90362) <= 9657463;
srom_1(90363) <= 10221987;
srom_1(90364) <= 10777913;
srom_1(90365) <= 11322636;
srom_1(90366) <= 11853600;
srom_1(90367) <= 12368315;
srom_1(90368) <= 12864368;
srom_1(90369) <= 13339433;
srom_1(90370) <= 13791281;
srom_1(90371) <= 14217795;
srom_1(90372) <= 14616973;
srom_1(90373) <= 14986945;
srom_1(90374) <= 15325975;
srom_1(90375) <= 15632472;
srom_1(90376) <= 15905001;
srom_1(90377) <= 16142283;
srom_1(90378) <= 16343206;
srom_1(90379) <= 16506826;
srom_1(90380) <= 16632378;
srom_1(90381) <= 16719271;
srom_1(90382) <= 16767099;
srom_1(90383) <= 16775638;
srom_1(90384) <= 16744847;
srom_1(90385) <= 16674870;
srom_1(90386) <= 16566037;
srom_1(90387) <= 16418857;
srom_1(90388) <= 16234020;
srom_1(90389) <= 16012393;
srom_1(90390) <= 15755016;
srom_1(90391) <= 15463095;
srom_1(90392) <= 15137999;
srom_1(90393) <= 14781253;
srom_1(90394) <= 14394530;
srom_1(90395) <= 13979643;
srom_1(90396) <= 13538538;
srom_1(90397) <= 13073282;
srom_1(90398) <= 12586059;
srom_1(90399) <= 12079153;
srom_1(90400) <= 11554940;
srom_1(90401) <= 11015879;
srom_1(90402) <= 10464498;
srom_1(90403) <= 9903383;
srom_1(90404) <= 9335164;
srom_1(90405) <= 8762507;
srom_1(90406) <= 8188096;
srom_1(90407) <= 7614625;
srom_1(90408) <= 7044784;
srom_1(90409) <= 6481244;
srom_1(90410) <= 5926649;
srom_1(90411) <= 5383599;
srom_1(90412) <= 4854640;
srom_1(90413) <= 4342253;
srom_1(90414) <= 3848841;
srom_1(90415) <= 3376718;
srom_1(90416) <= 2928097;
srom_1(90417) <= 2505082;
srom_1(90418) <= 2109657;
srom_1(90419) <= 1743676;
srom_1(90420) <= 1408856;
srom_1(90421) <= 1106766;
srom_1(90422) <= 838823;
srom_1(90423) <= 606283;
srom_1(90424) <= 410238;
srom_1(90425) <= 251606;
srom_1(90426) <= 131131;
srom_1(90427) <= 49378;
srom_1(90428) <= 6731;
srom_1(90429) <= 3389;
srom_1(90430) <= 39368;
srom_1(90431) <= 114500;
srom_1(90432) <= 228432;
srom_1(90433) <= 380630;
srom_1(90434) <= 570380;
srom_1(90435) <= 796792;
srom_1(90436) <= 1058805;
srom_1(90437) <= 1355190;
srom_1(90438) <= 1684557;
srom_1(90439) <= 2045362;
srom_1(90440) <= 2435912;
srom_1(90441) <= 2854376;
srom_1(90442) <= 3298793;
srom_1(90443) <= 3767077;
srom_1(90444) <= 4257033;
srom_1(90445) <= 4766364;
srom_1(90446) <= 5292680;
srom_1(90447) <= 5833515;
srom_1(90448) <= 6386331;
srom_1(90449) <= 6948536;
srom_1(90450) <= 7517495;
srom_1(90451) <= 8090538;
srom_1(90452) <= 8664979;
srom_1(90453) <= 9238124;
srom_1(90454) <= 9807286;
srom_1(90455) <= 10369794;
srom_1(90456) <= 10923013;
srom_1(90457) <= 11464346;
srom_1(90458) <= 11991257;
srom_1(90459) <= 12501273;
srom_1(90460) <= 12992004;
srom_1(90461) <= 13461147;
srom_1(90462) <= 13906504;
srom_1(90463) <= 14325986;
srom_1(90464) <= 14717625;
srom_1(90465) <= 15079585;
srom_1(90466) <= 15410169;
srom_1(90467) <= 15707826;
srom_1(90468) <= 15971161;
srom_1(90469) <= 16198939;
srom_1(90470) <= 16390091;
srom_1(90471) <= 16543722;
srom_1(90472) <= 16659111;
srom_1(90473) <= 16735716;
srom_1(90474) <= 16773179;
srom_1(90475) <= 16771324;
srom_1(90476) <= 16730159;
srom_1(90477) <= 16649878;
srom_1(90478) <= 16530857;
srom_1(90479) <= 16373654;
srom_1(90480) <= 16179007;
srom_1(90481) <= 15947827;
srom_1(90482) <= 15681200;
srom_1(90483) <= 15380376;
srom_1(90484) <= 15046764;
srom_1(90485) <= 14681930;
srom_1(90486) <= 14287585;
srom_1(90487) <= 13865577;
srom_1(90488) <= 13417886;
srom_1(90489) <= 12946611;
srom_1(90490) <= 12453962;
srom_1(90491) <= 11942249;
srom_1(90492) <= 11413872;
srom_1(90493) <= 10871308;
srom_1(90494) <= 10317102;
srom_1(90495) <= 9753853;
srom_1(90496) <= 9184201;
srom_1(90497) <= 8610819;
srom_1(90498) <= 8036395;
srom_1(90499) <= 7463622;
srom_1(90500) <= 6895187;
srom_1(90501) <= 6333755;
srom_1(90502) <= 5781959;
srom_1(90503) <= 5242386;
srom_1(90504) <= 4717567;
srom_1(90505) <= 4209963;
srom_1(90506) <= 3721954;
srom_1(90507) <= 3255829;
srom_1(90508) <= 2813773;
srom_1(90509) <= 2397859;
srom_1(90510) <= 2010038;
srom_1(90511) <= 1652128;
srom_1(90512) <= 1325808;
srom_1(90513) <= 1032607;
srom_1(90514) <= 773902;
srom_1(90515) <= 550904;
srom_1(90516) <= 364661;
srom_1(90517) <= 216044;
srom_1(90518) <= 105751;
srom_1(90519) <= 34299;
srom_1(90520) <= 2024;
srom_1(90521) <= 9076;
srom_1(90522) <= 55422;
srom_1(90523) <= 140846;
srom_1(90524) <= 264947;
srom_1(90525) <= 427142;
srom_1(90526) <= 626671;
srom_1(90527) <= 862598;
srom_1(90528) <= 1133817;
srom_1(90529) <= 1439057;
srom_1(90530) <= 1776885;
srom_1(90531) <= 2145719;
srom_1(90532) <= 2543827;
srom_1(90533) <= 2969343;
srom_1(90534) <= 3420272;
srom_1(90535) <= 3894499;
srom_1(90536) <= 4389801;
srom_1(90537) <= 4903855;
srom_1(90538) <= 5434249;
srom_1(90539) <= 5978498;
srom_1(90540) <= 6534049;
srom_1(90541) <= 7098296;
srom_1(90542) <= 7668594;
srom_1(90543) <= 8242268;
srom_1(90544) <= 8816629;
srom_1(90545) <= 9388982;
srom_1(90546) <= 9956644;
srom_1(90547) <= 10516953;
srom_1(90548) <= 11067282;
srom_1(90549) <= 11605050;
srom_1(90550) <= 12127734;
srom_1(90551) <= 12632884;
srom_1(90552) <= 13118132;
srom_1(90553) <= 13581201;
srom_1(90554) <= 14019920;
srom_1(90555) <= 14432232;
srom_1(90556) <= 14816204;
srom_1(90557) <= 15170034;
srom_1(90558) <= 15492064;
srom_1(90559) <= 15780783;
srom_1(90560) <= 16034838;
srom_1(90561) <= 16253037;
srom_1(90562) <= 16434357;
srom_1(90563) <= 16577948;
srom_1(90564) <= 16683136;
srom_1(90565) <= 16749428;
srom_1(90566) <= 16776513;
srom_1(90567) <= 16764265;
srom_1(90568) <= 16712740;
srom_1(90569) <= 16622181;
srom_1(90570) <= 16493011;
srom_1(90571) <= 16325837;
srom_1(90572) <= 16121443;
srom_1(90573) <= 15880787;
srom_1(90574) <= 15604997;
srom_1(90575) <= 15295368;
srom_1(90576) <= 14953350;
srom_1(90577) <= 14580547;
srom_1(90578) <= 14178709;
srom_1(90579) <= 13749719;
srom_1(90580) <= 13295589;
srom_1(90581) <= 12818448;
srom_1(90582) <= 12320534;
srom_1(90583) <= 11804182;
srom_1(90584) <= 11271813;
srom_1(90585) <= 10725924;
srom_1(90586) <= 10169075;
srom_1(90587) <= 9603876;
srom_1(90588) <= 9032978;
srom_1(90589) <= 8459059;
srom_1(90590) <= 7884809;
srom_1(90591) <= 7312922;
srom_1(90592) <= 6746079;
srom_1(90593) <= 6186938;
srom_1(90594) <= 5638122;
srom_1(90595) <= 5102204;
srom_1(90596) <= 4581697;
srom_1(90597) <= 4079041;
srom_1(90598) <= 3596595;
srom_1(90599) <= 3136620;
srom_1(90600) <= 2701274;
srom_1(90601) <= 2292597;
srom_1(90602) <= 1912507;
srom_1(90603) <= 1562785;
srom_1(90604) <= 1245072;
srom_1(90605) <= 960857;
srom_1(90606) <= 711474;
srom_1(90607) <= 498092;
srom_1(90608) <= 321710;
srom_1(90609) <= 183157;
srom_1(90610) <= 83083;
srom_1(90611) <= 21956;
srom_1(90612) <= 62;
srom_1(90613) <= 17506;
srom_1(90614) <= 74205;
srom_1(90615) <= 169893;
srom_1(90616) <= 304121;
srom_1(90617) <= 476260;
srom_1(90618) <= 685502;
srom_1(90619) <= 930868;
srom_1(90620) <= 1211205;
srom_1(90621) <= 1525199;
srom_1(90622) <= 1871379;
srom_1(90623) <= 2248119;
srom_1(90624) <= 2653655;
srom_1(90625) <= 3086084;
srom_1(90626) <= 3543378;
srom_1(90627) <= 4023393;
srom_1(90628) <= 4523878;
srom_1(90629) <= 5042487;
srom_1(90630) <= 5576786;
srom_1(90631) <= 6124271;
srom_1(90632) <= 6682374;
srom_1(90633) <= 7248478;
srom_1(90634) <= 7819929;
srom_1(90635) <= 8394046;
srom_1(90636) <= 8968138;
srom_1(90637) <= 9539512;
srom_1(90638) <= 10105490;
srom_1(90639) <= 10663416;
srom_1(90640) <= 11210675;
srom_1(90641) <= 11744700;
srom_1(90642) <= 12262987;
srom_1(90643) <= 12763106;
srom_1(90644) <= 13242712;
srom_1(90645) <= 13699555;
srom_1(90646) <= 14131493;
srom_1(90647) <= 14536500;
srom_1(90648) <= 14912679;
srom_1(90649) <= 15258263;
srom_1(90650) <= 15571633;
srom_1(90651) <= 15851320;
srom_1(90652) <= 16096012;
srom_1(90653) <= 16304560;
srom_1(90654) <= 16475988;
srom_1(90655) <= 16609492;
srom_1(90656) <= 16704445;
srom_1(90657) <= 16760402;
srom_1(90658) <= 16777101;
srom_1(90659) <= 16754464;
srom_1(90660) <= 16692596;
srom_1(90661) <= 16591788;
srom_1(90662) <= 16452512;
srom_1(90663) <= 16275422;
srom_1(90664) <= 16061348;
srom_1(90665) <= 15811294;
srom_1(90666) <= 15526432;
srom_1(90667) <= 15208098;
srom_1(90668) <= 14857786;
srom_1(90669) <= 14477137;
srom_1(90670) <= 14067937;
srom_1(90671) <= 13632105;
srom_1(90672) <= 13171685;
srom_1(90673) <= 12688834;
srom_1(90674) <= 12185819;
srom_1(90675) <= 11664997;
srom_1(90676) <= 11128811;
srom_1(90677) <= 10579775;
srom_1(90678) <= 10020464;
srom_1(90679) <= 9453501;
srom_1(90680) <= 8881544;
srom_1(90681) <= 8307275;
srom_1(90682) <= 7733388;
srom_1(90683) <= 7162574;
srom_1(90684) <= 6597509;
srom_1(90685) <= 6040842;
srom_1(90686) <= 5495186;
srom_1(90687) <= 4963097;
srom_1(90688) <= 4447072;
srom_1(90689) <= 3949530;
srom_1(90690) <= 3472805;
srom_1(90691) <= 3019131;
srom_1(90692) <= 2590637;
srom_1(90693) <= 2189331;
srom_1(90694) <= 1817096;
srom_1(90695) <= 1475677;
srom_1(90696) <= 1166675;
srom_1(90697) <= 891539;
srom_1(90698) <= 651560;
srom_1(90699) <= 447862;
srom_1(90700) <= 281401;
srom_1(90701) <= 152957;
srom_1(90702) <= 63134;
srom_1(90703) <= 12351;
srom_1(90704) <= 848;
srom_1(90705) <= 28677;
srom_1(90706) <= 95709;
srom_1(90707) <= 201630;
srom_1(90708) <= 345941;
srom_1(90709) <= 527968;
srom_1(90710) <= 746856;
srom_1(90711) <= 1001579;
srom_1(90712) <= 1290942;
srom_1(90713) <= 1613588;
srom_1(90714) <= 1968005;
srom_1(90715) <= 2352530;
srom_1(90716) <= 2765361;
srom_1(90717) <= 3204561;
srom_1(90718) <= 3668070;
srom_1(90719) <= 4153716;
srom_1(90720) <= 4659221;
srom_1(90721) <= 5182214;
srom_1(90722) <= 5720243;
srom_1(90723) <= 6270784;
srom_1(90724) <= 6831257;
srom_1(90725) <= 7399033;
srom_1(90726) <= 7971450;
srom_1(90727) <= 8545822;
srom_1(90728) <= 9119458;
srom_1(90729) <= 9689666;
srom_1(90730) <= 10253773;
srom_1(90731) <= 10809133;
srom_1(90732) <= 11353143;
srom_1(90733) <= 11883251;
srom_1(90734) <= 12396972;
srom_1(90735) <= 12891896;
srom_1(90736) <= 13365702;
srom_1(90737) <= 13816170;
srom_1(90738) <= 14241185;
srom_1(90739) <= 14638756;
srom_1(90740) <= 15007017;
srom_1(90741) <= 15344243;
srom_1(90742) <= 15648851;
srom_1(90743) <= 15919414;
srom_1(90744) <= 16154662;
srom_1(90745) <= 16353492;
srom_1(90746) <= 16514972;
srom_1(90747) <= 16638345;
srom_1(90748) <= 16723032;
srom_1(90749) <= 16768636;
srom_1(90750) <= 16774943;
srom_1(90751) <= 16741924;
srom_1(90752) <= 16669733;
srom_1(90753) <= 16558709;
srom_1(90754) <= 16409373;
srom_1(90755) <= 16222424;
srom_1(90756) <= 15998741;
srom_1(90757) <= 15739370;
srom_1(90758) <= 15445529;
srom_1(90759) <= 15118596;
srom_1(90760) <= 14760104;
srom_1(90761) <= 14371734;
srom_1(90762) <= 13955306;
srom_1(90763) <= 13512775;
srom_1(90764) <= 13046214;
srom_1(90765) <= 12557813;
srom_1(90766) <= 12049860;
srom_1(90767) <= 11524739;
srom_1(90768) <= 10984911;
srom_1(90769) <= 10432909;
srom_1(90770) <= 9871319;
srom_1(90771) <= 9302777;
srom_1(90772) <= 8729948;
srom_1(90773) <= 8155519;
srom_1(90774) <= 7582182;
srom_1(90775) <= 7012627;
srom_1(90776) <= 6449525;
srom_1(90777) <= 5895515;
srom_1(90778) <= 5353197;
srom_1(90779) <= 4825112;
srom_1(90780) <= 4313738;
srom_1(90781) <= 3821472;
srom_1(90782) <= 3350624;
srom_1(90783) <= 2903400;
srom_1(90784) <= 2481898;
srom_1(90785) <= 2088095;
srom_1(90786) <= 1723837;
srom_1(90787) <= 1390832;
srom_1(90788) <= 1090642;
srom_1(90789) <= 824675;
srom_1(90790) <= 594178;
srom_1(90791) <= 400232;
srom_1(90792) <= 243746;
srom_1(90793) <= 125454;
srom_1(90794) <= 45910;
srom_1(90795) <= 5489;
srom_1(90796) <= 4379;
srom_1(90797) <= 42585;
srom_1(90798) <= 119929;
srom_1(90799) <= 236047;
srom_1(90800) <= 390395;
srom_1(90801) <= 582250;
srom_1(90802) <= 810712;
srom_1(90803) <= 1074709;
srom_1(90804) <= 1373003;
srom_1(90805) <= 1704196;
srom_1(90806) <= 2066734;
srom_1(90807) <= 2458918;
srom_1(90808) <= 2878908;
srom_1(90809) <= 3324735;
srom_1(90810) <= 3794308;
srom_1(90811) <= 4285426;
srom_1(90812) <= 4795784;
srom_1(90813) <= 5322991;
srom_1(90814) <= 5864573;
srom_1(90815) <= 6417992;
srom_1(90816) <= 6980651;
srom_1(90817) <= 7549913;
srom_1(90818) <= 8123107;
srom_1(90819) <= 8697547;
srom_1(90820) <= 9270538;
srom_1(90821) <= 9839393;
srom_1(90822) <= 10401445;
srom_1(90823) <= 10954058;
srom_1(90824) <= 11494641;
srom_1(90825) <= 12020659;
srom_1(90826) <= 12529644;
srom_1(90827) <= 13019211;
srom_1(90828) <= 13487064;
srom_1(90829) <= 13931008;
srom_1(90830) <= 14348961;
srom_1(90831) <= 14738965;
srom_1(90832) <= 15099190;
srom_1(90833) <= 15427946;
srom_1(90834) <= 15723692;
srom_1(90835) <= 15985042;
srom_1(90836) <= 16210770;
srom_1(90837) <= 16399816;
srom_1(90838) <= 16551296;
srom_1(90839) <= 16664497;
srom_1(90840) <= 16738890;
srom_1(90841) <= 16774126;
srom_1(90842) <= 16770039;
srom_1(90843) <= 16726649;
srom_1(90844) <= 16644159;
srom_1(90845) <= 16522956;
srom_1(90846) <= 16363608;
srom_1(90847) <= 16166862;
srom_1(90848) <= 15933642;
srom_1(90849) <= 15665040;
srom_1(90850) <= 15362317;
srom_1(90851) <= 15026891;
srom_1(90852) <= 14660336;
srom_1(90853) <= 14264371;
srom_1(90854) <= 13840853;
srom_1(90855) <= 13391767;
srom_1(90856) <= 12919219;
srom_1(90857) <= 12425426;
srom_1(90858) <= 11912703;
srom_1(90859) <= 11383454;
srom_1(90860) <= 10840162;
srom_1(90861) <= 10285373;
srom_1(90862) <= 9721689;
srom_1(90863) <= 9151755;
srom_1(90864) <= 8578241;
srom_1(90865) <= 8003838;
srom_1(90866) <= 7431240;
srom_1(90867) <= 6863131;
srom_1(90868) <= 6302176;
srom_1(90869) <= 5751004;
srom_1(90870) <= 5212201;
srom_1(90871) <= 4688294;
srom_1(90872) <= 4181738;
srom_1(90873) <= 3694910;
srom_1(90874) <= 3230092;
srom_1(90875) <= 2789464;
srom_1(90876) <= 2375093;
srom_1(90877) <= 1988921;
srom_1(90878) <= 1632759;
srom_1(90879) <= 1308278;
srom_1(90880) <= 1016999;
srom_1(90881) <= 760288;
srom_1(90882) <= 539349;
srom_1(90883) <= 355217;
srom_1(90884) <= 208757;
srom_1(90885) <= 100655;
srom_1(90886) <= 31418;
srom_1(90887) <= 1371;
srom_1(90888) <= 10655;
srom_1(90889) <= 59225;
srom_1(90890) <= 146855;
srom_1(90891) <= 273133;
srom_1(90892) <= 437468;
srom_1(90893) <= 639088;
srom_1(90894) <= 877048;
srom_1(90895) <= 1150233;
srom_1(90896) <= 1457361;
srom_1(90897) <= 1796991;
srom_1(90898) <= 2167533;
srom_1(90899) <= 2567246;
srom_1(90900) <= 2994259;
srom_1(90901) <= 3446567;
srom_1(90902) <= 3922050;
srom_1(90903) <= 4418478;
srom_1(90904) <= 4933524;
srom_1(90905) <= 5464772;
srom_1(90906) <= 6009730;
srom_1(90907) <= 6565844;
srom_1(90908) <= 7130506;
srom_1(90909) <= 7701067;
srom_1(90910) <= 8274852;
srom_1(90911) <= 8849171;
srom_1(90912) <= 9421330;
srom_1(90913) <= 9988646;
srom_1(90914) <= 10548459;
srom_1(90915) <= 11098144;
srom_1(90916) <= 11635122;
srom_1(90917) <= 12156877;
srom_1(90918) <= 12660961;
srom_1(90919) <= 13145011;
srom_1(90920) <= 13606756;
srom_1(90921) <= 14044031;
srom_1(90922) <= 14454786;
srom_1(90923) <= 14837095;
srom_1(90924) <= 15189165;
srom_1(90925) <= 15509344;
srom_1(90926) <= 15796132;
srom_1(90927) <= 16048183;
srom_1(90928) <= 16264316;
srom_1(90929) <= 16443518;
srom_1(90930) <= 16584946;
srom_1(90931) <= 16687940;
srom_1(90932) <= 16752015;
srom_1(90933) <= 16776871;
srom_1(90934) <= 16762392;
srom_1(90935) <= 16708645;
srom_1(90936) <= 16615882;
srom_1(90937) <= 16484539;
srom_1(90938) <= 16315232;
srom_1(90939) <= 16108754;
srom_1(90940) <= 15866073;
srom_1(90941) <= 15588328;
srom_1(90942) <= 15276821;
srom_1(90943) <= 14933013;
srom_1(90944) <= 14558515;
srom_1(90945) <= 14155085;
srom_1(90946) <= 13724614;
srom_1(90947) <= 13269121;
srom_1(90948) <= 12790741;
srom_1(90949) <= 12291718;
srom_1(90950) <= 11774392;
srom_1(90951) <= 11241189;
srom_1(90952) <= 10694609;
srom_1(90953) <= 10137216;
srom_1(90954) <= 9571623;
srom_1(90955) <= 9000482;
srom_1(90956) <= 8426472;
srom_1(90957) <= 7852284;
srom_1(90958) <= 7280611;
srom_1(90959) <= 6714134;
srom_1(90960) <= 6155510;
srom_1(90961) <= 5607357;
srom_1(90962) <= 5072246;
srom_1(90963) <= 4552687;
srom_1(90964) <= 4051115;
srom_1(90965) <= 3569884;
srom_1(90966) <= 3111249;
srom_1(90967) <= 2677362;
srom_1(90968) <= 2270257;
srom_1(90969) <= 1891843;
srom_1(90970) <= 1543894;
srom_1(90971) <= 1228042;
srom_1(90972) <= 945769;
srom_1(90973) <= 698398;
srom_1(90974) <= 487089;
srom_1(90975) <= 312833;
srom_1(90976) <= 176447;
srom_1(90977) <= 78570;
srom_1(90978) <= 19662;
srom_1(90979) <= 0;
srom_1(90980) <= 19674;
srom_1(90981) <= 78592;
srom_1(90982) <= 176480;
srom_1(90983) <= 312877;
srom_1(90984) <= 487143;
srom_1(90985) <= 698463;
srom_1(90986) <= 945844;
srom_1(90987) <= 1228127;
srom_1(90988) <= 1543988;
srom_1(90989) <= 1891945;
srom_1(90990) <= 2270368;
srom_1(90991) <= 2677481;
srom_1(90992) <= 3111375;
srom_1(90993) <= 3570017;
srom_1(90994) <= 4051254;
srom_1(90995) <= 4552831;
srom_1(90996) <= 5072395;
srom_1(90997) <= 5607510;
srom_1(90998) <= 6155666;
srom_1(90999) <= 6714293;
srom_1(91000) <= 7280772;
srom_1(91001) <= 7852446;
srom_1(91002) <= 8426634;
srom_1(91003) <= 9000643;
srom_1(91004) <= 9571783;
srom_1(91005) <= 10137374;
srom_1(91006) <= 10694765;
srom_1(91007) <= 11241342;
srom_1(91008) <= 11774541;
srom_1(91009) <= 12291862;
srom_1(91010) <= 12790879;
srom_1(91011) <= 13269253;
srom_1(91012) <= 13724739;
srom_1(91013) <= 14155203;
srom_1(91014) <= 14558625;
srom_1(91015) <= 14933114;
srom_1(91016) <= 15276913;
srom_1(91017) <= 15588411;
srom_1(91018) <= 15866146;
srom_1(91019) <= 16108817;
srom_1(91020) <= 16315285;
srom_1(91021) <= 16484582;
srom_1(91022) <= 16615914;
srom_1(91023) <= 16708665;
srom_1(91024) <= 16762401;
srom_1(91025) <= 16776869;
srom_1(91026) <= 16752002;
srom_1(91027) <= 16687916;
srom_1(91028) <= 16584912;
srom_1(91029) <= 16443472;
srom_1(91030) <= 16264261;
srom_1(91031) <= 16048117;
srom_1(91032) <= 15796056;
srom_1(91033) <= 15509258;
srom_1(91034) <= 15189070;
srom_1(91035) <= 14836991;
srom_1(91036) <= 14454674;
srom_1(91037) <= 14043911;
srom_1(91038) <= 13606629;
srom_1(91039) <= 13144877;
srom_1(91040) <= 12660822;
srom_1(91041) <= 12156732;
srom_1(91042) <= 11634973;
srom_1(91043) <= 11097990;
srom_1(91044) <= 10548302;
srom_1(91045) <= 9988487;
srom_1(91046) <= 9421169;
srom_1(91047) <= 8849009;
srom_1(91048) <= 8274690;
srom_1(91049) <= 7700905;
srom_1(91050) <= 7130345;
srom_1(91051) <= 6565686;
srom_1(91052) <= 6009575;
srom_1(91053) <= 5464620;
srom_1(91054) <= 4933376;
srom_1(91055) <= 4418335;
srom_1(91056) <= 3921913;
srom_1(91057) <= 3446436;
srom_1(91058) <= 2994134;
srom_1(91059) <= 2567130;
srom_1(91060) <= 2167424;
srom_1(91061) <= 1796891;
srom_1(91062) <= 1457269;
srom_1(91063) <= 1150151;
srom_1(91064) <= 876976;
srom_1(91065) <= 639026;
srom_1(91066) <= 437416;
srom_1(91067) <= 273092;
srom_1(91068) <= 146825;
srom_1(91069) <= 59206;
srom_1(91070) <= 10646;
srom_1(91071) <= 1374;
srom_1(91072) <= 31432;
srom_1(91073) <= 100680;
srom_1(91074) <= 208793;
srom_1(91075) <= 355264;
srom_1(91076) <= 539406;
srom_1(91077) <= 760355;
srom_1(91078) <= 1017077;
srom_1(91079) <= 1308365;
srom_1(91080) <= 1632855;
srom_1(91081) <= 1989026;
srom_1(91082) <= 2375206;
srom_1(91083) <= 2789585;
srom_1(91084) <= 3230220;
srom_1(91085) <= 3695044;
srom_1(91086) <= 4181878;
srom_1(91087) <= 4688439;
srom_1(91088) <= 5212351;
srom_1(91089) <= 5751158;
srom_1(91090) <= 6302333;
srom_1(91091) <= 6863290;
srom_1(91092) <= 7431401;
srom_1(91093) <= 8004000;
srom_1(91094) <= 8578403;
srom_1(91095) <= 9151916;
srom_1(91096) <= 9721849;
srom_1(91097) <= 10285531;
srom_1(91098) <= 10840317;
srom_1(91099) <= 11383606;
srom_1(91100) <= 11912850;
srom_1(91101) <= 12425568;
srom_1(91102) <= 12919356;
srom_1(91103) <= 13391897;
srom_1(91104) <= 13840976;
srom_1(91105) <= 14264487;
srom_1(91106) <= 14660444;
srom_1(91107) <= 15026990;
srom_1(91108) <= 15362407;
srom_1(91109) <= 15665121;
srom_1(91110) <= 15933713;
srom_1(91111) <= 16166923;
srom_1(91112) <= 16363658;
srom_1(91113) <= 16522995;
srom_1(91114) <= 16644188;
srom_1(91115) <= 16726667;
srom_1(91116) <= 16770046;
srom_1(91117) <= 16774122;
srom_1(91118) <= 16738875;
srom_1(91119) <= 16664471;
srom_1(91120) <= 16551258;
srom_1(91121) <= 16399768;
srom_1(91122) <= 16210711;
srom_1(91123) <= 15984973;
srom_1(91124) <= 15723614;
srom_1(91125) <= 15427858;
srom_1(91126) <= 15099092;
srom_1(91127) <= 14738859;
srom_1(91128) <= 14348847;
srom_1(91129) <= 13930886;
srom_1(91130) <= 13486935;
srom_1(91131) <= 13019076;
srom_1(91132) <= 12529503;
srom_1(91133) <= 12020513;
srom_1(91134) <= 11494491;
srom_1(91135) <= 10953904;
srom_1(91136) <= 10401288;
srom_1(91137) <= 9839234;
srom_1(91138) <= 9270377;
srom_1(91139) <= 8697385;
srom_1(91140) <= 8122945;
srom_1(91141) <= 7549751;
srom_1(91142) <= 6980491;
srom_1(91143) <= 6417834;
srom_1(91144) <= 5864419;
srom_1(91145) <= 5322840;
srom_1(91146) <= 4795638;
srom_1(91147) <= 4285284;
srom_1(91148) <= 3794172;
srom_1(91149) <= 3324606;
srom_1(91150) <= 2878786;
srom_1(91151) <= 2458803;
srom_1(91152) <= 2066627;
srom_1(91153) <= 1704098;
srom_1(91154) <= 1372914;
srom_1(91155) <= 1074629;
srom_1(91156) <= 810642;
srom_1(91157) <= 582191;
srom_1(91158) <= 390346;
srom_1(91159) <= 236009;
srom_1(91160) <= 119901;
srom_1(91161) <= 42569;
srom_1(91162) <= 4373;
srom_1(91163) <= 5495;
srom_1(91164) <= 45927;
srom_1(91165) <= 125482;
srom_1(91166) <= 243785;
srom_1(91167) <= 400281;
srom_1(91168) <= 594238;
srom_1(91169) <= 824746;
srom_1(91170) <= 1090722;
srom_1(91171) <= 1390921;
srom_1(91172) <= 1723935;
srom_1(91173) <= 2088202;
srom_1(91174) <= 2482013;
srom_1(91175) <= 2903523;
srom_1(91176) <= 3350753;
srom_1(91177) <= 3821608;
srom_1(91178) <= 4313880;
srom_1(91179) <= 4825259;
srom_1(91180) <= 5353348;
srom_1(91181) <= 5895670;
srom_1(91182) <= 6449682;
srom_1(91183) <= 7012787;
srom_1(91184) <= 7582344;
srom_1(91185) <= 8155681;
srom_1(91186) <= 8730110;
srom_1(91187) <= 9302938;
srom_1(91188) <= 9871479;
srom_1(91189) <= 10433066;
srom_1(91190) <= 10985065;
srom_1(91191) <= 11524889;
srom_1(91192) <= 12050006;
srom_1(91193) <= 12557953;
srom_1(91194) <= 13046349;
srom_1(91195) <= 13512903;
srom_1(91196) <= 13955428;
srom_1(91197) <= 14371847;
srom_1(91198) <= 14760210;
srom_1(91199) <= 15118693;
srom_1(91200) <= 15445617;
srom_1(91201) <= 15739448;
srom_1(91202) <= 15998809;
srom_1(91203) <= 16222482;
srom_1(91204) <= 16409420;
srom_1(91205) <= 16558746;
srom_1(91206) <= 16669759;
srom_1(91207) <= 16741939;
srom_1(91208) <= 16774947;
srom_1(91209) <= 16768629;
srom_1(91210) <= 16723014;
srom_1(91211) <= 16638316;
srom_1(91212) <= 16514932;
srom_1(91213) <= 16353441;
srom_1(91214) <= 16154601;
srom_1(91215) <= 15919342;
srom_1(91216) <= 15648770;
srom_1(91217) <= 15344153;
srom_1(91218) <= 15006918;
srom_1(91219) <= 14638648;
srom_1(91220) <= 14241069;
srom_1(91221) <= 13816046;
srom_1(91222) <= 13365572;
srom_1(91223) <= 12891759;
srom_1(91224) <= 12396830;
srom_1(91225) <= 11883104;
srom_1(91226) <= 11352992;
srom_1(91227) <= 10808978;
srom_1(91228) <= 10253615;
srom_1(91229) <= 9689506;
srom_1(91230) <= 9119296;
srom_1(91231) <= 8545660;
srom_1(91232) <= 7971288;
srom_1(91233) <= 7398872;
srom_1(91234) <= 6831098;
srom_1(91235) <= 6270628;
srom_1(91236) <= 5720089;
srom_1(91237) <= 5182064;
srom_1(91238) <= 4659076;
srom_1(91239) <= 4153576;
srom_1(91240) <= 3667936;
srom_1(91241) <= 3204433;
srom_1(91242) <= 2765241;
srom_1(91243) <= 2352418;
srom_1(91244) <= 1967901;
srom_1(91245) <= 1613493;
srom_1(91246) <= 1290856;
srom_1(91247) <= 1001502;
srom_1(91248) <= 746789;
srom_1(91249) <= 527912;
srom_1(91250) <= 345895;
srom_1(91251) <= 201594;
srom_1(91252) <= 95685;
srom_1(91253) <= 28664;
srom_1(91254) <= 845;
srom_1(91255) <= 12360;
srom_1(91256) <= 63154;
srom_1(91257) <= 152988;
srom_1(91258) <= 281443;
srom_1(91259) <= 447914;
srom_1(91260) <= 651622;
srom_1(91261) <= 891612;
srom_1(91262) <= 1166757;
srom_1(91263) <= 1475769;
srom_1(91264) <= 1817197;
srom_1(91265) <= 2189440;
srom_1(91266) <= 2590754;
srom_1(91267) <= 3019256;
srom_1(91268) <= 3472936;
srom_1(91269) <= 3949668;
srom_1(91270) <= 4447215;
srom_1(91271) <= 4963245;
srom_1(91272) <= 5495338;
srom_1(91273) <= 6040998;
srom_1(91274) <= 6597667;
srom_1(91275) <= 7162734;
srom_1(91276) <= 7733550;
srom_1(91277) <= 8307438;
srom_1(91278) <= 8881706;
srom_1(91279) <= 9453662;
srom_1(91280) <= 10020623;
srom_1(91281) <= 10579932;
srom_1(91282) <= 11128964;
srom_1(91283) <= 11665146;
srom_1(91284) <= 12185963;
srom_1(91285) <= 12688973;
srom_1(91286) <= 13171818;
srom_1(91287) <= 13632232;
srom_1(91288) <= 14068057;
srom_1(91289) <= 14477249;
srom_1(91290) <= 14857889;
srom_1(91291) <= 15208193;
srom_1(91292) <= 15526517;
srom_1(91293) <= 15811369;
srom_1(91294) <= 16061413;
srom_1(91295) <= 16275477;
srom_1(91296) <= 16452557;
srom_1(91297) <= 16591822;
srom_1(91298) <= 16692619;
srom_1(91299) <= 16754476;
srom_1(91300) <= 16777102;
srom_1(91301) <= 16760392;
srom_1(91302) <= 16704424;
srom_1(91303) <= 16609460;
srom_1(91304) <= 16475945;
srom_1(91305) <= 16304507;
srom_1(91306) <= 16095948;
srom_1(91307) <= 15851246;
srom_1(91308) <= 15571550;
srom_1(91309) <= 15258170;
srom_1(91310) <= 14912577;
srom_1(91311) <= 14536390;
srom_1(91312) <= 14131375;
srom_1(91313) <= 13699429;
srom_1(91314) <= 13242580;
srom_1(91315) <= 12762968;
srom_1(91316) <= 12262843;
srom_1(91317) <= 11744551;
srom_1(91318) <= 11210522;
srom_1(91319) <= 10663260;
srom_1(91320) <= 10105331;
srom_1(91321) <= 9539352;
srom_1(91322) <= 8967976;
srom_1(91323) <= 8393884;
srom_1(91324) <= 7819767;
srom_1(91325) <= 7248317;
srom_1(91326) <= 6682215;
srom_1(91327) <= 6124115;
srom_1(91328) <= 5576633;
srom_1(91329) <= 5042338;
srom_1(91330) <= 4523734;
srom_1(91331) <= 4023255;
srom_1(91332) <= 3543246;
srom_1(91333) <= 3085958;
srom_1(91334) <= 2653537;
srom_1(91335) <= 2248009;
srom_1(91336) <= 1871276;
srom_1(91337) <= 1525106;
srom_1(91338) <= 1211121;
srom_1(91339) <= 930793;
srom_1(91340) <= 685438;
srom_1(91341) <= 476206;
srom_1(91342) <= 304077;
srom_1(91343) <= 169860;
srom_1(91344) <= 74183;
srom_1(91345) <= 17496;
srom_1(91346) <= 63;
srom_1(91347) <= 21967;
srom_1(91348) <= 83106;
srom_1(91349) <= 183191;
srom_1(91350) <= 321755;
srom_1(91351) <= 498147;
srom_1(91352) <= 711539;
srom_1(91353) <= 960933;
srom_1(91354) <= 1245157;
srom_1(91355) <= 1562879;
srom_1(91356) <= 1912610;
srom_1(91357) <= 2292708;
srom_1(91358) <= 2701393;
srom_1(91359) <= 3136747;
srom_1(91360) <= 3596728;
srom_1(91361) <= 4079180;
srom_1(91362) <= 4581841;
srom_1(91363) <= 5102353;
srom_1(91364) <= 5638275;
srom_1(91365) <= 6187095;
srom_1(91366) <= 6746238;
srom_1(91367) <= 7313083;
srom_1(91368) <= 7884971;
srom_1(91369) <= 8459221;
srom_1(91370) <= 9033140;
srom_1(91371) <= 9604036;
srom_1(91372) <= 10169233;
srom_1(91373) <= 10726080;
srom_1(91374) <= 11271966;
srom_1(91375) <= 11804330;
srom_1(91376) <= 12320677;
srom_1(91377) <= 12818586;
srom_1(91378) <= 13295720;
srom_1(91379) <= 13749844;
srom_1(91380) <= 14178826;
srom_1(91381) <= 14580657;
srom_1(91382) <= 14953451;
srom_1(91383) <= 15295460;
srom_1(91384) <= 15605080;
srom_1(91385) <= 15880860;
srom_1(91386) <= 16121506;
srom_1(91387) <= 16325890;
srom_1(91388) <= 16493053;
srom_1(91389) <= 16622212;
srom_1(91390) <= 16712760;
srom_1(91391) <= 16764274;
srom_1(91392) <= 16776511;
srom_1(91393) <= 16749415;
srom_1(91394) <= 16683111;
srom_1(91395) <= 16577912;
srom_1(91396) <= 16434311;
srom_1(91397) <= 16252980;
srom_1(91398) <= 16034771;
srom_1(91399) <= 15780706;
srom_1(91400) <= 15491978;
srom_1(91401) <= 15169939;
srom_1(91402) <= 14816100;
srom_1(91403) <= 14432120;
srom_1(91404) <= 14019800;
srom_1(91405) <= 13581074;
srom_1(91406) <= 13117998;
srom_1(91407) <= 12632745;
srom_1(91408) <= 12127589;
srom_1(91409) <= 11604900;
srom_1(91410) <= 11067129;
srom_1(91411) <= 10516797;
srom_1(91412) <= 9956485;
srom_1(91413) <= 9388821;
srom_1(91414) <= 8816467;
srom_1(91415) <= 8242106;
srom_1(91416) <= 7668432;
srom_1(91417) <= 7098136;
srom_1(91418) <= 6533891;
srom_1(91419) <= 5978343;
srom_1(91420) <= 5434098;
srom_1(91421) <= 4903707;
srom_1(91422) <= 4389659;
srom_1(91423) <= 3894363;
srom_1(91424) <= 3420142;
srom_1(91425) <= 2969219;
srom_1(91426) <= 2543710;
srom_1(91427) <= 2145610;
srom_1(91428) <= 1776786;
srom_1(91429) <= 1438966;
srom_1(91430) <= 1133736;
srom_1(91431) <= 862526;
srom_1(91432) <= 626609;
srom_1(91433) <= 427090;
srom_1(91434) <= 264906;
srom_1(91435) <= 140817;
srom_1(91436) <= 55404;
srom_1(91437) <= 9068;
srom_1(91438) <= 2027;
srom_1(91439) <= 34314;
srom_1(91440) <= 105777;
srom_1(91441) <= 216080;
srom_1(91442) <= 364708;
srom_1(91443) <= 550962;
srom_1(91444) <= 773970;
srom_1(91445) <= 1032685;
srom_1(91446) <= 1325895;
srom_1(91447) <= 1652225;
srom_1(91448) <= 2010143;
srom_1(91449) <= 2397972;
srom_1(91450) <= 2813894;
srom_1(91451) <= 3255957;
srom_1(91452) <= 3722089;
srom_1(91453) <= 4210104;
srom_1(91454) <= 4717713;
srom_1(91455) <= 5242537;
srom_1(91456) <= 5782113;
srom_1(91457) <= 6333912;
srom_1(91458) <= 6895346;
srom_1(91459) <= 7463783;
srom_1(91460) <= 8036557;
srom_1(91461) <= 8610981;
srom_1(91462) <= 9184363;
srom_1(91463) <= 9754013;
srom_1(91464) <= 10317260;
srom_1(91465) <= 10871463;
srom_1(91466) <= 11414023;
srom_1(91467) <= 11942396;
srom_1(91468) <= 12454104;
srom_1(91469) <= 12946747;
srom_1(91470) <= 13418016;
srom_1(91471) <= 13865700;
srom_1(91472) <= 14287700;
srom_1(91473) <= 14682038;
srom_1(91474) <= 15046863;
srom_1(91475) <= 15380465;
srom_1(91476) <= 15681280;
srom_1(91477) <= 15947898;
srom_1(91478) <= 16179067;
srom_1(91479) <= 16373704;
srom_1(91480) <= 16530896;
srom_1(91481) <= 16649906;
srom_1(91482) <= 16730176;
srom_1(91483) <= 16771330;
srom_1(91484) <= 16773174;
srom_1(91485) <= 16735700;
srom_1(91486) <= 16659083;
srom_1(91487) <= 16543684;
srom_1(91488) <= 16390042;
srom_1(91489) <= 16198880;
srom_1(91490) <= 15971092;
srom_1(91491) <= 15707747;
srom_1(91492) <= 15410080;
srom_1(91493) <= 15079487;
srom_1(91494) <= 14717518;
srom_1(91495) <= 14325871;
srom_1(91496) <= 13906382;
srom_1(91497) <= 13461018;
srom_1(91498) <= 12991868;
srom_1(91499) <= 12501132;
srom_1(91500) <= 11991110;
srom_1(91501) <= 11464195;
srom_1(91502) <= 10922858;
srom_1(91503) <= 10369637;
srom_1(91504) <= 9807126;
srom_1(91505) <= 9237963;
srom_1(91506) <= 8664817;
srom_1(91507) <= 8090376;
srom_1(91508) <= 7517333;
srom_1(91509) <= 6948377;
srom_1(91510) <= 6386173;
srom_1(91511) <= 5833360;
srom_1(91512) <= 5292530;
srom_1(91513) <= 4766218;
srom_1(91514) <= 4256892;
srom_1(91515) <= 3766942;
srom_1(91516) <= 3298664;
srom_1(91517) <= 2854255;
srom_1(91518) <= 2435798;
srom_1(91519) <= 2045256;
srom_1(91520) <= 1684460;
srom_1(91521) <= 1355102;
srom_1(91522) <= 1058726;
srom_1(91523) <= 796723;
srom_1(91524) <= 570321;
srom_1(91525) <= 380582;
srom_1(91526) <= 228395;
srom_1(91527) <= 114474;
srom_1(91528) <= 39353;
srom_1(91529) <= 3384;
srom_1(91530) <= 6737;
srom_1(91531) <= 49396;
srom_1(91532) <= 131159;
srom_1(91533) <= 251645;
srom_1(91534) <= 410288;
srom_1(91535) <= 606344;
srom_1(91536) <= 838894;
srom_1(91537) <= 1106846;
srom_1(91538) <= 1408946;
srom_1(91539) <= 1743775;
srom_1(91540) <= 2109765;
srom_1(91541) <= 2505198;
srom_1(91542) <= 2928220;
srom_1(91543) <= 3376848;
srom_1(91544) <= 3848978;
srom_1(91545) <= 4342395;
srom_1(91546) <= 4854787;
srom_1(91547) <= 5383750;
srom_1(91548) <= 5926804;
srom_1(91549) <= 6481402;
srom_1(91550) <= 7044944;
srom_1(91551) <= 7614787;
srom_1(91552) <= 8188258;
srom_1(91553) <= 8762669;
srom_1(91554) <= 9335325;
srom_1(91555) <= 9903542;
srom_1(91556) <= 10464655;
srom_1(91557) <= 11016033;
srom_1(91558) <= 11555090;
srom_1(91559) <= 12079298;
srom_1(91560) <= 12586200;
srom_1(91561) <= 13073417;
srom_1(91562) <= 13538665;
srom_1(91563) <= 13979764;
srom_1(91564) <= 14394643;
srom_1(91565) <= 14781358;
srom_1(91566) <= 15138095;
srom_1(91567) <= 15463182;
srom_1(91568) <= 15755093;
srom_1(91569) <= 16012460;
srom_1(91570) <= 16234077;
srom_1(91571) <= 16418903;
srom_1(91572) <= 16566073;
srom_1(91573) <= 16674896;
srom_1(91574) <= 16744861;
srom_1(91575) <= 16775641;
srom_1(91576) <= 16767091;
srom_1(91577) <= 16719252;
srom_1(91578) <= 16632348;
srom_1(91579) <= 16506786;
srom_1(91580) <= 16343154;
srom_1(91581) <= 16142222;
srom_1(91582) <= 15904929;
srom_1(91583) <= 15632391;
srom_1(91584) <= 15325883;
srom_1(91585) <= 14986845;
srom_1(91586) <= 14616865;
srom_1(91587) <= 14217678;
srom_1(91588) <= 13791157;
srom_1(91589) <= 13339302;
srom_1(91590) <= 12864231;
srom_1(91591) <= 12368172;
srom_1(91592) <= 11853452;
srom_1(91593) <= 11322484;
srom_1(91594) <= 10777758;
srom_1(91595) <= 10221828;
srom_1(91596) <= 9657302;
srom_1(91597) <= 9086827;
srom_1(91598) <= 8513077;
srom_1(91599) <= 7938744;
srom_1(91600) <= 7366520;
srom_1(91601) <= 6799089;
srom_1(91602) <= 6239112;
srom_1(91603) <= 5689214;
srom_1(91604) <= 5151975;
srom_1(91605) <= 4629914;
srom_1(91606) <= 4125478;
srom_1(91607) <= 3641034;
srom_1(91608) <= 3178853;
srom_1(91609) <= 2741102;
srom_1(91610) <= 2329834;
srom_1(91611) <= 1946978;
srom_1(91612) <= 1594328;
srom_1(91613) <= 1273540;
srom_1(91614) <= 986116;
srom_1(91615) <= 733406;
srom_1(91616) <= 516593;
srom_1(91617) <= 336695;
srom_1(91618) <= 194555;
srom_1(91619) <= 90839;
srom_1(91620) <= 26035;
srom_1(91621) <= 446;
srom_1(91622) <= 14191;
srom_1(91623) <= 67208;
srom_1(91624) <= 159246;
srom_1(91625) <= 289874;
srom_1(91626) <= 458480;
srom_1(91627) <= 664273;
srom_1(91628) <= 906289;
srom_1(91629) <= 1183391;
srom_1(91630) <= 1494281;
srom_1(91631) <= 1837501;
srom_1(91632) <= 2211442;
srom_1(91633) <= 2614349;
srom_1(91634) <= 3044334;
srom_1(91635) <= 3499380;
srom_1(91636) <= 3977353;
srom_1(91637) <= 4476012;
srom_1(91638) <= 4993018;
srom_1(91639) <= 5525948;
srom_1(91640) <= 6072301;
srom_1(91641) <= 6629517;
srom_1(91642) <= 7194981;
srom_1(91643) <= 7766043;
srom_1(91644) <= 8340024;
srom_1(91645) <= 8914233;
srom_1(91646) <= 9485978;
srom_1(91647) <= 10052576;
srom_1(91648) <= 10611371;
srom_1(91649) <= 11159743;
srom_1(91650) <= 11695120;
srom_1(91651) <= 12214992;
srom_1(91652) <= 12716921;
srom_1(91653) <= 13198553;
srom_1(91654) <= 13657629;
srom_1(91655) <= 14091997;
srom_1(91656) <= 14499619;
srom_1(91657) <= 14878585;
srom_1(91658) <= 15227118;
srom_1(91659) <= 15543582;
srom_1(91660) <= 15826494;
srom_1(91661) <= 16074527;
srom_1(91662) <= 16286519;
srom_1(91663) <= 16461474;
srom_1(91664) <= 16598573;
srom_1(91665) <= 16697173;
srom_1(91666) <= 16756810;
srom_1(91667) <= 16777207;
srom_1(91668) <= 16758266;
srom_1(91669) <= 16700077;
srom_1(91670) <= 16602913;
srom_1(91671) <= 16467229;
srom_1(91672) <= 16293662;
srom_1(91673) <= 16083025;
srom_1(91674) <= 15836307;
srom_1(91675) <= 15554663;
srom_1(91676) <= 15239416;
srom_1(91677) <= 14892042;
srom_1(91678) <= 14514172;
srom_1(91679) <= 14107577;
srom_1(91680) <= 13674164;
srom_1(91681) <= 13215965;
srom_1(91682) <= 12735129;
srom_1(91683) <= 12233910;
srom_1(91684) <= 11714660;
srom_1(91685) <= 11179812;
srom_1(91686) <= 10631876;
srom_1(91687) <= 10073420;
srom_1(91688) <= 9507063;
srom_1(91689) <= 8935462;
srom_1(91690) <= 8361296;
srom_1(91691) <= 7787259;
srom_1(91692) <= 7216041;
srom_1(91693) <= 6650322;
srom_1(91694) <= 6092754;
srom_1(91695) <= 5545952;
srom_1(91696) <= 5012480;
srom_1(91697) <= 4494841;
srom_1(91698) <= 3995460;
srom_1(91699) <= 3516681;
srom_1(91700) <= 3060747;
srom_1(91701) <= 2629798;
srom_1(91702) <= 2225854;
srom_1(91703) <= 1850809;
srom_1(91704) <= 1506422;
srom_1(91705) <= 1194308;
srom_1(91706) <= 915930;
srom_1(91707) <= 672594;
srom_1(91708) <= 465442;
srom_1(91709) <= 295444;
srom_1(91710) <= 163397;
srom_1(91711) <= 69922;
srom_1(91712) <= 15455;
srom_1(91713) <= 253;
srom_1(91714) <= 24387;
srom_1(91715) <= 87744;
srom_1(91716) <= 190026;
srom_1(91717) <= 330754;
srom_1(91718) <= 509269;
srom_1(91719) <= 724732;
srom_1(91720) <= 976134;
srom_1(91721) <= 1262295;
srom_1(91722) <= 1581874;
srom_1(91723) <= 1933372;
srom_1(91724) <= 2315141;
srom_1(91725) <= 2725391;
srom_1(91726) <= 3162197;
srom_1(91727) <= 3623512;
srom_1(91728) <= 4107172;
srom_1(91729) <= 4610909;
srom_1(91730) <= 5132361;
srom_1(91731) <= 5669082;
srom_1(91732) <= 6218557;
srom_1(91733) <= 6778207;
srom_1(91734) <= 7345410;
srom_1(91735) <= 7917504;
srom_1(91736) <= 8491807;
srom_1(91737) <= 9065626;
srom_1(91738) <= 9636271;
srom_1(91739) <= 10201065;
srom_1(91740) <= 10757359;
srom_1(91741) <= 11302546;
srom_1(91742) <= 11834068;
srom_1(91743) <= 12349434;
srom_1(91744) <= 12846225;
srom_1(91745) <= 13322114;
srom_1(91746) <= 13774867;
srom_1(91747) <= 14202362;
srom_1(91748) <= 14602595;
srom_1(91749) <= 14973688;
srom_1(91750) <= 15313902;
srom_1(91751) <= 15621640;
srom_1(91752) <= 15895460;
srom_1(91753) <= 16134078;
srom_1(91754) <= 16336375;
srom_1(91755) <= 16501402;
srom_1(91756) <= 16628385;
srom_1(91757) <= 16716729;
srom_1(91758) <= 16766020;
srom_1(91759) <= 16776026;
srom_1(91760) <= 16746701;
srom_1(91761) <= 16678181;
srom_1(91762) <= 16570789;
srom_1(91763) <= 16425028;
srom_1(91764) <= 16241582;
srom_1(91765) <= 16021310;
srom_1(91766) <= 15765245;
srom_1(91767) <= 15474590;
srom_1(91768) <= 15150705;
srom_1(91769) <= 14795111;
srom_1(91770) <= 14409474;
srom_1(91771) <= 13995604;
srom_1(91772) <= 13555440;
srom_1(91773) <= 13091047;
srom_1(91774) <= 12604603;
srom_1(91775) <= 12098389;
srom_1(91776) <= 11574778;
srom_1(91777) <= 11036226;
srom_1(91778) <= 10485259;
srom_1(91779) <= 9924460;
srom_1(91780) <= 9356458;
srom_1(91781) <= 8783918;
srom_1(91782) <= 8209524;
srom_1(91783) <= 7635970;
srom_1(91784) <= 7065946;
srom_1(91785) <= 6502123;
srom_1(91786) <= 5947147;
srom_1(91787) <= 5403620;
srom_1(91788) <= 4874091;
srom_1(91789) <= 4361042;
srom_1(91790) <= 3866880;
srom_1(91791) <= 3393922;
srom_1(91792) <= 2944386;
srom_1(91793) <= 2520379;
srom_1(91794) <= 2123891;
srom_1(91795) <= 1756780;
srom_1(91796) <= 1420768;
srom_1(91797) <= 1117431;
srom_1(91798) <= 848190;
srom_1(91799) <= 614309;
srom_1(91800) <= 416885;
srom_1(91801) <= 256843;
srom_1(91802) <= 134933;
srom_1(91803) <= 51728;
srom_1(91804) <= 7617;
srom_1(91805) <= 2807;
srom_1(91806) <= 37322;
srom_1(91807) <= 110998;
srom_1(91808) <= 223491;
srom_1(91809) <= 374273;
srom_1(91810) <= 562637;
srom_1(91811) <= 787699;
srom_1(91812) <= 1048405;
srom_1(91813) <= 1343532;
srom_1(91814) <= 1671695;
srom_1(91815) <= 2031357;
srom_1(91816) <= 2420829;
srom_1(91817) <= 2838287;
srom_1(91818) <= 3281772;
srom_1(91819) <= 3749204;
srom_1(91820) <= 4238393;
srom_1(91821) <= 4747043;
srom_1(91822) <= 5272769;
srom_1(91823) <= 5813107;
srom_1(91824) <= 6365523;
srom_1(91825) <= 6927425;
srom_1(91826) <= 7496179;
srom_1(91827) <= 8069118;
srom_1(91828) <= 8643556;
srom_1(91829) <= 9216798;
srom_1(91830) <= 9786156;
srom_1(91831) <= 10348960;
srom_1(91832) <= 10902572;
srom_1(91833) <= 11444395;
srom_1(91834) <= 11971888;
srom_1(91835) <= 12482578;
srom_1(91836) <= 12974070;
srom_1(91837) <= 13444059;
srom_1(91838) <= 13890342;
srom_1(91839) <= 14310825;
srom_1(91840) <= 14703536;
srom_1(91841) <= 15066635;
srom_1(91842) <= 15398418;
srom_1(91843) <= 15697330;
srom_1(91844) <= 15961968;
srom_1(91845) <= 16191093;
srom_1(91846) <= 16383629;
srom_1(91847) <= 16538673;
srom_1(91848) <= 16655499;
srom_1(91849) <= 16733559;
srom_1(91850) <= 16772487;
srom_1(91851) <= 16772099;
srom_1(91852) <= 16732399;
srom_1(91853) <= 16653571;
srom_1(91854) <= 16535987;
srom_1(91855) <= 16380196;
srom_1(91856) <= 16186930;
srom_1(91857) <= 15957095;
srom_1(91858) <= 15691769;
srom_1(91859) <= 15392196;
srom_1(91860) <= 15059781;
srom_1(91861) <= 14696082;
srom_1(91862) <= 14302805;
srom_1(91863) <= 13881795;
srom_1(91864) <= 13435025;
srom_1(91865) <= 12964590;
srom_1(91866) <= 12472698;
srom_1(91867) <= 11961653;
srom_1(91868) <= 11433854;
srom_1(91869) <= 10891774;
srom_1(91870) <= 10337956;
srom_1(91871) <= 9774997;
srom_1(91872) <= 9205536;
srom_1(91873) <= 8632245;
srom_1(91874) <= 8057811;
srom_1(91875) <= 7484928;
srom_1(91876) <= 6916284;
srom_1(91877) <= 6354543;
srom_1(91878) <= 5802340;
srom_1(91879) <= 5262266;
srom_1(91880) <= 4736852;
srom_1(91881) <= 4228563;
srom_1(91882) <= 3739781;
srom_1(91883) <= 3272799;
srom_1(91884) <= 2829807;
srom_1(91885) <= 2412882;
srom_1(91886) <= 2023979;
srom_1(91887) <= 1664923;
srom_1(91888) <= 1337396;
srom_1(91889) <= 1042934;
srom_1(91890) <= 782919;
srom_1(91891) <= 558570;
srom_1(91892) <= 370938;
srom_1(91893) <= 220904;
srom_1(91894) <= 109171;
srom_1(91895) <= 36263;
srom_1(91896) <= 2522;
srom_1(91897) <= 8106;
srom_1(91898) <= 52990;
srom_1(91899) <= 136962;
srom_1(91900) <= 259629;
srom_1(91901) <= 420415;
srom_1(91902) <= 618567;
srom_1(91903) <= 853155;
srom_1(91904) <= 1123080;
srom_1(91905) <= 1427075;
srom_1(91906) <= 1763716;
srom_1(91907) <= 2131422;
srom_1(91908) <= 2528471;
srom_1(91909) <= 2953000;
srom_1(91910) <= 3403018;
srom_1(91911) <= 3876416;
srom_1(91912) <= 4370972;
srom_1(91913) <= 4884369;
srom_1(91914) <= 5414198;
srom_1(91915) <= 5957976;
srom_1(91916) <= 6513151;
srom_1(91917) <= 7077121;
srom_1(91918) <= 7647241;
srom_1(91919) <= 8220838;
srom_1(91920) <= 8795221;
srom_1(91921) <= 9367698;
srom_1(91922) <= 9935583;
srom_1(91923) <= 10496214;
srom_1(91924) <= 11046961;
srom_1(91925) <= 11585243;
srom_1(91926) <= 12108535;
srom_1(91927) <= 12614382;
srom_1(91928) <= 13100414;
srom_1(91929) <= 13564350;
srom_1(91930) <= 14004015;
srom_1(91931) <= 14417348;
srom_1(91932) <= 14802410;
srom_1(91933) <= 15157395;
srom_1(91934) <= 15480640;
srom_1(91935) <= 15770627;
srom_1(91936) <= 16025997;
srom_1(91937) <= 16245553;
srom_1(91938) <= 16428265;
srom_1(91939) <= 16573277;
srom_1(91940) <= 16679907;
srom_1(91941) <= 16747657;
srom_1(91942) <= 16776209;
srom_1(91943) <= 16765428;
srom_1(91944) <= 16715365;
srom_1(91945) <= 16626255;
srom_1(91946) <= 16498517;
srom_1(91947) <= 16332748;
srom_1(91948) <= 16129726;
srom_1(91949) <= 15890403;
srom_1(91950) <= 15615902;
srom_1(91951) <= 15307510;
srom_1(91952) <= 14966672;
srom_1(91953) <= 14594988;
srom_1(91954) <= 14194200;
srom_1(91955) <= 13766187;
srom_1(91956) <= 13312957;
srom_1(91957) <= 12836635;
srom_1(91958) <= 12339455;
srom_1(91959) <= 11823748;
srom_1(91960) <= 11291932;
srom_1(91961) <= 10746502;
srom_1(91962) <= 10190015;
srom_1(91963) <= 9625080;
srom_1(91964) <= 9054347;
srom_1(91965) <= 8480492;
srom_1(91966) <= 7906206;
srom_1(91967) <= 7334183;
srom_1(91968) <= 6767103;
srom_1(91969) <= 6207628;
srom_1(91970) <= 5658380;
srom_1(91971) <= 5121935;
srom_1(91972) <= 4600809;
srom_1(91973) <= 4097445;
srom_1(91974) <= 3614203;
srom_1(91975) <= 3153351;
srom_1(91976) <= 2717048;
srom_1(91977) <= 2307341;
srom_1(91978) <= 1926152;
srom_1(91979) <= 1575267;
srom_1(91980) <= 1256332;
srom_1(91981) <= 970843;
srom_1(91982) <= 720138;
srom_1(91983) <= 505393;
srom_1(91984) <= 327616;
srom_1(91985) <= 187639;
srom_1(91986) <= 86119;
srom_1(91987) <= 23533;
srom_1(91988) <= 173;
srom_1(91989) <= 16149;
srom_1(91990) <= 71387;
srom_1(91991) <= 165627;
srom_1(91992) <= 298428;
srom_1(91993) <= 469166;
srom_1(91994) <= 677041;
srom_1(91995) <= 921078;
srom_1(91996) <= 1200134;
srom_1(91997) <= 1512898;
srom_1(91998) <= 1857905;
srom_1(91999) <= 2233536;
srom_1(92000) <= 2638031;
srom_1(92001) <= 3069492;
srom_1(92002) <= 3525897;
srom_1(92003) <= 4005104;
srom_1(92004) <= 4504867;
srom_1(92005) <= 5022842;
srom_1(92006) <= 5556601;
srom_1(92007) <= 6103640;
srom_1(92008) <= 6661393;
srom_1(92009) <= 7227247;
srom_1(92010) <= 7798546;
srom_1(92011) <= 8372612;
srom_1(92012) <= 8946753;
srom_1(92013) <= 9518277;
srom_1(92014) <= 10084504;
srom_1(92015) <= 10642777;
srom_1(92016) <= 11190481;
srom_1(92017) <= 11725045;
srom_1(92018) <= 12243964;
srom_1(92019) <= 12744803;
srom_1(92020) <= 13225215;
srom_1(92021) <= 13682946;
srom_1(92022) <= 14115850;
srom_1(92023) <= 14521898;
srom_1(92024) <= 14899184;
srom_1(92025) <= 15245940;
srom_1(92026) <= 15560539;
srom_1(92027) <= 15841507;
srom_1(92028) <= 16087526;
srom_1(92029) <= 16297441;
srom_1(92030) <= 16470270;
srom_1(92031) <= 16605200;
srom_1(92032) <= 16701601;
srom_1(92033) <= 16759019;
srom_1(92034) <= 16777185;
srom_1(92035) <= 16756014;
srom_1(92036) <= 16695606;
srom_1(92037) <= 16596243;
srom_1(92038) <= 16458391;
srom_1(92039) <= 16282698;
srom_1(92040) <= 16069987;
srom_1(92041) <= 15821255;
srom_1(92042) <= 15537669;
srom_1(92043) <= 15220558;
srom_1(92044) <= 14871410;
srom_1(92045) <= 14491862;
srom_1(92046) <= 14083693;
srom_1(92047) <= 13648819;
srom_1(92048) <= 13189277;
srom_1(92049) <= 12707224;
srom_1(92050) <= 12204919;
srom_1(92051) <= 11684718;
srom_1(92052) <= 11149060;
srom_1(92053) <= 10600458;
srom_1(92054) <= 10041483;
srom_1(92055) <= 9474758;
srom_1(92056) <= 8902939;
srom_1(92057) <= 8328709;
srom_1(92058) <= 7754759;
srom_1(92059) <= 7183782;
srom_1(92060) <= 6618454;
srom_1(92061) <= 6061428;
srom_1(92062) <= 5515314;
srom_1(92063) <= 4982674;
srom_1(92064) <= 4466006;
srom_1(92065) <= 3967732;
srom_1(92066) <= 3490189;
srom_1(92067) <= 3035616;
srom_1(92068) <= 2606146;
srom_1(92069) <= 2203791;
srom_1(92070) <= 1830440;
srom_1(92071) <= 1487841;
srom_1(92072) <= 1177603;
srom_1(92073) <= 901180;
srom_1(92074) <= 659867;
srom_1(92075) <= 454798;
srom_1(92076) <= 286932;
srom_1(92077) <= 157059;
srom_1(92078) <= 65786;
srom_1(92079) <= 13541;
srom_1(92080) <= 570;
srom_1(92081) <= 26934;
srom_1(92082) <= 92508;
srom_1(92083) <= 196985;
srom_1(92084) <= 339876;
srom_1(92085) <= 520510;
srom_1(92086) <= 738040;
srom_1(92087) <= 991446;
srom_1(92088) <= 1279540;
srom_1(92089) <= 1600971;
srom_1(92090) <= 1954232;
srom_1(92091) <= 2337666;
srom_1(92092) <= 2749474;
srom_1(92093) <= 3187726;
srom_1(92094) <= 3650367;
srom_1(92095) <= 4135228;
srom_1(92096) <= 4640034;
srom_1(92097) <= 5162418;
srom_1(92098) <= 5699931;
srom_1(92099) <= 6250052;
srom_1(92100) <= 6810201;
srom_1(92101) <= 7377752;
srom_1(92102) <= 7950044;
srom_1(92103) <= 8524391;
srom_1(92104) <= 9098103;
srom_1(92105) <= 9668487;
srom_1(92106) <= 10232869;
srom_1(92107) <= 10788603;
srom_1(92108) <= 11333083;
srom_1(92109) <= 11863754;
srom_1(92110) <= 12378130;
srom_1(92111) <= 12873798;
srom_1(92112) <= 13348432;
srom_1(92113) <= 13799809;
srom_1(92114) <= 14225810;
srom_1(92115) <= 14624439;
srom_1(92116) <= 14993826;
srom_1(92117) <= 15332239;
srom_1(92118) <= 15638091;
srom_1(92119) <= 15909947;
srom_1(92120) <= 16146533;
srom_1(92121) <= 16346740;
srom_1(92122) <= 16509628;
srom_1(92123) <= 16634434;
srom_1(92124) <= 16720573;
srom_1(92125) <= 16767640;
srom_1(92126) <= 16775414;
srom_1(92127) <= 16743861;
srom_1(92128) <= 16673126;
srom_1(92129) <= 16563543;
srom_1(92130) <= 16415624;
srom_1(92131) <= 16230064;
srom_1(92132) <= 16007733;
srom_1(92133) <= 15749673;
srom_1(92134) <= 15457095;
srom_1(92135) <= 15131370;
srom_1(92136) <= 14774025;
srom_1(92137) <= 14386738;
srom_1(92138) <= 13971323;
srom_1(92139) <= 13529729;
srom_1(92140) <= 13064026;
srom_1(92141) <= 12576399;
srom_1(92142) <= 12069133;
srom_1(92143) <= 11544609;
srom_1(92144) <= 11005284;
srom_1(92145) <= 10453690;
srom_1(92146) <= 9892411;
srom_1(92147) <= 9324081;
srom_1(92148) <= 8751364;
srom_1(92149) <= 8176945;
srom_1(92150) <= 7603520;
srom_1(92151) <= 7033775;
srom_1(92152) <= 6470385;
srom_1(92153) <= 5915989;
srom_1(92154) <= 5373188;
srom_1(92155) <= 4844528;
srom_1(92156) <= 4332487;
srom_1(92157) <= 3839466;
srom_1(92158) <= 3367778;
srom_1(92159) <= 2919635;
srom_1(92160) <= 2497137;
srom_1(92161) <= 2102266;
srom_1(92162) <= 1736875;
srom_1(92163) <= 1402675;
srom_1(92164) <= 1101235;
srom_1(92165) <= 833968;
srom_1(92166) <= 602127;
srom_1(92167) <= 406800;
srom_1(92168) <= 248902;
srom_1(92169) <= 129174;
srom_1(92170) <= 48177;
srom_1(92171) <= 6292;
srom_1(92172) <= 3713;
srom_1(92173) <= 40455;
srom_1(92174) <= 116344;
srom_1(92175) <= 231025;
srom_1(92176) <= 383959;
srom_1(92177) <= 574429;
srom_1(92178) <= 801544;
srom_1(92179) <= 1064236;
srom_1(92180) <= 1361275;
srom_1(92181) <= 1691267;
srom_1(92182) <= 2052666;
srom_1(92183) <= 2443776;
srom_1(92184) <= 2862763;
srom_1(92185) <= 3307663;
srom_1(92186) <= 3776389;
srom_1(92187) <= 4266744;
srom_1(92188) <= 4776427;
srom_1(92189) <= 5303049;
srom_1(92190) <= 5844141;
srom_1(92191) <= 6397164;
srom_1(92192) <= 6959526;
srom_1(92193) <= 7528589;
srom_1(92194) <= 8101685;
srom_1(92195) <= 8676127;
srom_1(92196) <= 9249220;
srom_1(92197) <= 9818277;
srom_1(92198) <= 10380631;
srom_1(92199) <= 10933643;
srom_1(92200) <= 11474720;
srom_1(92201) <= 12001326;
srom_1(92202) <= 12510991;
srom_1(92203) <= 13001324;
srom_1(92204) <= 13470026;
srom_1(92205) <= 13914900;
srom_1(92206) <= 14333859;
srom_1(92207) <= 14724939;
srom_1(92208) <= 15086306;
srom_1(92209) <= 15416265;
srom_1(92210) <= 15713269;
srom_1(92211) <= 15975925;
srom_1(92212) <= 16203001;
srom_1(92213) <= 16393433;
srom_1(92214) <= 16546328;
srom_1(92215) <= 16660968;
srom_1(92216) <= 16736817;
srom_1(92217) <= 16773517;
srom_1(92218) <= 16770898;
srom_1(92219) <= 16728972;
srom_1(92220) <= 16647935;
srom_1(92221) <= 16528166;
srom_1(92222) <= 16370229;
srom_1(92223) <= 16174863;
srom_1(92224) <= 15942985;
srom_1(92225) <= 15675681;
srom_1(92226) <= 15374206;
srom_1(92227) <= 15039974;
srom_1(92228) <= 14674550;
srom_1(92229) <= 14279650;
srom_1(92230) <= 13857124;
srom_1(92231) <= 13408955;
srom_1(92232) <= 12937244;
srom_1(92233) <= 12444202;
srom_1(92234) <= 11932143;
srom_1(92235) <= 11403466;
srom_1(92236) <= 10860652;
srom_1(92237) <= 10306246;
srom_1(92238) <= 9742847;
srom_1(92239) <= 9173097;
srom_1(92240) <= 8599669;
srom_1(92241) <= 8025251;
srom_1(92242) <= 7452537;
srom_1(92243) <= 6884213;
srom_1(92244) <= 6322943;
srom_1(92245) <= 5771360;
srom_1(92246) <= 5232050;
srom_1(92247) <= 4707542;
srom_1(92248) <= 4200296;
srom_1(92249) <= 3712690;
srom_1(92250) <= 3247011;
srom_1(92251) <= 2805443;
srom_1(92252) <= 2390057;
srom_1(92253) <= 2002799;
srom_1(92254) <= 1645487;
srom_1(92255) <= 1319796;
srom_1(92256) <= 1027253;
srom_1(92257) <= 769229;
srom_1(92258) <= 546936;
srom_1(92259) <= 361415;
srom_1(92260) <= 213536;
srom_1(92261) <= 103993;
srom_1(92262) <= 33299;
srom_1(92263) <= 1786;
srom_1(92264) <= 9602;
srom_1(92265) <= 56710;
srom_1(92266) <= 142889;
srom_1(92267) <= 267735;
srom_1(92268) <= 430662;
srom_1(92269) <= 630907;
srom_1(92270) <= 867531;
srom_1(92271) <= 1139424;
srom_1(92272) <= 1445310;
srom_1(92273) <= 1783756;
srom_1(92274) <= 2153174;
srom_1(92275) <= 2551833;
srom_1(92276) <= 2977862;
srom_1(92277) <= 3429263;
srom_1(92278) <= 3903921;
srom_1(92279) <= 4399610;
srom_1(92280) <= 4914004;
srom_1(92281) <= 5444691;
srom_1(92282) <= 5989184;
srom_1(92283) <= 6544928;
srom_1(92284) <= 7109318;
srom_1(92285) <= 7679707;
srom_1(92286) <= 8253420;
srom_1(92287) <= 8827767;
srom_1(92288) <= 9400055;
srom_1(92289) <= 9967600;
srom_1(92290) <= 10527740;
srom_1(92291) <= 11077850;
srom_1(92292) <= 11615348;
srom_1(92293) <= 12137715;
srom_1(92294) <= 12642501;
srom_1(92295) <= 13127340;
srom_1(92296) <= 13589956;
srom_1(92297) <= 14028182;
srom_1(92298) <= 14439962;
srom_1(92299) <= 14823365;
srom_1(92300) <= 15176593;
srom_1(92301) <= 15497990;
srom_1(92302) <= 15786049;
srom_1(92303) <= 16039419;
srom_1(92304) <= 16256911;
srom_1(92305) <= 16437506;
srom_1(92306) <= 16580357;
srom_1(92307) <= 16684794;
srom_1(92308) <= 16750327;
srom_1(92309) <= 16776650;
srom_1(92310) <= 16763638;
srom_1(92311) <= 16711352;
srom_1(92312) <= 16620039;
srom_1(92313) <= 16490125;
srom_1(92314) <= 16322221;
srom_1(92315) <= 16117113;
srom_1(92316) <= 15875763;
srom_1(92317) <= 15599304;
srom_1(92318) <= 15289031;
srom_1(92319) <= 14946400;
srom_1(92320) <= 14573017;
srom_1(92321) <= 14170633;
srom_1(92322) <= 13741136;
srom_1(92323) <= 13286538;
srom_1(92324) <= 12808972;
srom_1(92325) <= 12310678;
srom_1(92326) <= 11793992;
srom_1(92327) <= 11261337;
srom_1(92328) <= 10715210;
srom_1(92329) <= 10158173;
srom_1(92330) <= 9592839;
srom_1(92331) <= 9021857;
srom_1(92332) <= 8447905;
srom_1(92333) <= 7873676;
srom_1(92334) <= 7301861;
srom_1(92335) <= 6735143;
srom_1(92336) <= 6176178;
srom_1(92337) <= 5627587;
srom_1(92338) <= 5091945;
srom_1(92339) <= 4571761;
srom_1(92340) <= 4069476;
srom_1(92341) <= 3587445;
srom_1(92342) <= 3127928;
srom_1(92343) <= 2693080;
srom_1(92344) <= 2284940;
srom_1(92345) <= 1905423;
srom_1(92346) <= 1556308;
srom_1(92347) <= 1239231;
srom_1(92348) <= 955681;
srom_1(92349) <= 706986;
srom_1(92350) <= 494312;
srom_1(92351) <= 318658;
srom_1(92352) <= 180847;
srom_1(92353) <= 81524;
srom_1(92354) <= 21157;
srom_1(92355) <= 27;
srom_1(92356) <= 18234;
srom_1(92357) <= 75692;
srom_1(92358) <= 172133;
srom_1(92359) <= 307104;
srom_1(92360) <= 479971;
srom_1(92361) <= 689925;
srom_1(92362) <= 935981;
srom_1(92363) <= 1216984;
srom_1(92364) <= 1531618;
srom_1(92365) <= 1878407;
srom_1(92366) <= 2255724;
srom_1(92367) <= 2661800;
srom_1(92368) <= 3094731;
srom_1(92369) <= 3552487;
srom_1(92370) <= 4032922;
srom_1(92371) <= 4533781;
srom_1(92372) <= 5052717;
srom_1(92373) <= 5587297;
srom_1(92374) <= 6135012;
srom_1(92375) <= 6693296;
srom_1(92376) <= 7259529;
srom_1(92377) <= 7831057;
srom_1(92378) <= 8405200;
srom_1(92379) <= 8979265;
srom_1(92380) <= 9550559;
srom_1(92381) <= 10116406;
srom_1(92382) <= 10674150;
srom_1(92383) <= 11221176;
srom_1(92384) <= 11754919;
srom_1(92385) <= 12272877;
srom_1(92386) <= 12772619;
srom_1(92387) <= 13251804;
srom_1(92388) <= 13708184;
srom_1(92389) <= 14139618;
srom_1(92390) <= 14544083;
srom_1(92391) <= 14919684;
srom_1(92392) <= 15264658;
srom_1(92393) <= 15577388;
srom_1(92394) <= 15856407;
srom_1(92395) <= 16100407;
srom_1(92396) <= 16308244;
srom_1(92397) <= 16478943;
srom_1(92398) <= 16611704;
srom_1(92399) <= 16705904;
srom_1(92400) <= 16761101;
srom_1(92401) <= 16777036;
srom_1(92402) <= 16753635;
srom_1(92403) <= 16691008;
srom_1(92404) <= 16589448;
srom_1(92405) <= 16449432;
srom_1(92406) <= 16271615;
srom_1(92407) <= 16056832;
srom_1(92408) <= 15806091;
srom_1(92409) <= 15520566;
srom_1(92410) <= 15201597;
srom_1(92411) <= 14850680;
srom_1(92412) <= 14469459;
srom_1(92413) <= 14059724;
srom_1(92414) <= 13623394;
srom_1(92415) <= 13162517;
srom_1(92416) <= 12679254;
srom_1(92417) <= 12175870;
srom_1(92418) <= 11654726;
srom_1(92419) <= 11118267;
srom_1(92420) <= 10569007;
srom_1(92421) <= 10009522;
srom_1(92422) <= 9442436;
srom_1(92423) <= 8870409;
srom_1(92424) <= 8296122;
srom_1(92425) <= 7722269;
srom_1(92426) <= 7151541;
srom_1(92427) <= 6586614;
srom_1(92428) <= 6030136;
srom_1(92429) <= 5484719;
srom_1(92430) <= 4952919;
srom_1(92431) <= 4437230;
srom_1(92432) <= 3940070;
srom_1(92433) <= 3463771;
srom_1(92434) <= 3010566;
srom_1(92435) <= 2582581;
srom_1(92436) <= 2181822;
srom_1(92437) <= 1810169;
srom_1(92438) <= 1469365;
srom_1(92439) <= 1161007;
srom_1(92440) <= 886542;
srom_1(92441) <= 647257;
srom_1(92442) <= 444273;
srom_1(92443) <= 278543;
srom_1(92444) <= 150844;
srom_1(92445) <= 61775;
srom_1(92446) <= 11753;
srom_1(92447) <= 1014;
srom_1(92448) <= 29606;
srom_1(92449) <= 97397;
srom_1(92450) <= 204068;
srom_1(92451) <= 349119;
srom_1(92452) <= 531870;
srom_1(92453) <= 751464;
srom_1(92454) <= 1006871;
srom_1(92455) <= 1296893;
srom_1(92456) <= 1620171;
srom_1(92457) <= 1975189;
srom_1(92458) <= 2360281;
srom_1(92459) <= 2773643;
srom_1(92460) <= 3213334;
srom_1(92461) <= 3677295;
srom_1(92462) <= 4163348;
srom_1(92463) <= 4669215;
srom_1(92464) <= 5192523;
srom_1(92465) <= 5730819;
srom_1(92466) <= 6281579;
srom_1(92467) <= 6842219;
srom_1(92468) <= 7410110;
srom_1(92469) <= 7982590;
srom_1(92470) <= 8556974;
srom_1(92471) <= 9130568;
srom_1(92472) <= 9700683;
srom_1(92473) <= 10264646;
srom_1(92474) <= 10819810;
srom_1(92475) <= 11363575;
srom_1(92476) <= 11893388;
srom_1(92477) <= 12406766;
srom_1(92478) <= 12901302;
srom_1(92479) <= 13374676;
srom_1(92480) <= 13824669;
srom_1(92481) <= 14249171;
srom_1(92482) <= 14646190;
srom_1(92483) <= 15013865;
srom_1(92484) <= 15350472;
srom_1(92485) <= 15654432;
srom_1(92486) <= 15924321;
srom_1(92487) <= 16158872;
srom_1(92488) <= 16356985;
srom_1(92489) <= 16517732;
srom_1(92490) <= 16640359;
srom_1(92491) <= 16724290;
srom_1(92492) <= 16769133;
srom_1(92493) <= 16774676;
srom_1(92494) <= 16740894;
srom_1(92495) <= 16667946;
srom_1(92496) <= 16556173;
srom_1(92497) <= 16406099;
srom_1(92498) <= 16218429;
srom_1(92499) <= 15994041;
srom_1(92500) <= 15733990;
srom_1(92501) <= 15439493;
srom_1(92502) <= 15111932;
srom_1(92503) <= 14752843;
srom_1(92504) <= 14363911;
srom_1(92505) <= 13946958;
srom_1(92506) <= 13503939;
srom_1(92507) <= 13036934;
srom_1(92508) <= 12548131;
srom_1(92509) <= 12039822;
srom_1(92510) <= 11514391;
srom_1(92511) <= 10974303;
srom_1(92512) <= 10422089;
srom_1(92513) <= 9860340;
srom_1(92514) <= 9291689;
srom_1(92515) <= 8718804;
srom_1(92516) <= 8144370;
srom_1(92517) <= 7571081;
srom_1(92518) <= 7001626;
srom_1(92519) <= 6438675;
srom_1(92520) <= 5884868;
srom_1(92521) <= 5342801;
srom_1(92522) <= 4815018;
srom_1(92523) <= 4303992;
srom_1(92524) <= 3812121;
srom_1(92525) <= 3341710;
srom_1(92526) <= 2894966;
srom_1(92527) <= 2473983;
srom_1(92528) <= 2080736;
srom_1(92529) <= 1717069;
srom_1(92530) <= 1384687;
srom_1(92531) <= 1085149;
srom_1(92532) <= 819859;
srom_1(92533) <= 590062;
srom_1(92534) <= 396835;
srom_1(92535) <= 241084;
srom_1(92536) <= 123539;
srom_1(92537) <= 44752;
srom_1(92538) <= 5093;
srom_1(92539) <= 4746;
srom_1(92540) <= 43715;
srom_1(92541) <= 121815;
srom_1(92542) <= 238681;
srom_1(92543) <= 393765;
srom_1(92544) <= 586340;
srom_1(92545) <= 815502;
srom_1(92546) <= 1080177;
srom_1(92547) <= 1379124;
srom_1(92548) <= 1710940;
srom_1(92549) <= 2074071;
srom_1(92550) <= 2466812;
srom_1(92551) <= 2887323;
srom_1(92552) <= 3333632;
srom_1(92553) <= 3803644;
srom_1(92554) <= 4295157;
srom_1(92555) <= 4805866;
srom_1(92556) <= 5333376;
srom_1(92557) <= 5875212;
srom_1(92558) <= 6428835;
srom_1(92559) <= 6991648;
srom_1(92560) <= 7561011;
srom_1(92561) <= 8134256;
srom_1(92562) <= 8708693;
srom_1(92563) <= 9281629;
srom_1(92564) <= 9850378;
srom_1(92565) <= 10412271;
srom_1(92566) <= 10964675;
srom_1(92567) <= 11504999;
srom_1(92568) <= 12030710;
srom_1(92569) <= 12539341;
srom_1(92570) <= 13028508;
srom_1(92571) <= 13495916;
srom_1(92572) <= 13939375;
srom_1(92573) <= 14356805;
srom_1(92574) <= 14746247;
srom_1(92575) <= 15105876;
srom_1(92576) <= 15434006;
srom_1(92577) <= 15729098;
srom_1(92578) <= 15989767;
srom_1(92579) <= 16214792;
srom_1(92580) <= 16403117;
srom_1(92581) <= 16553859;
srom_1(92582) <= 16666312;
srom_1(92583) <= 16739948;
srom_1(92584) <= 16774421;
srom_1(92585) <= 16769571;
srom_1(92586) <= 16725419;
srom_1(92587) <= 16642173;
srom_1(92588) <= 16520223;
srom_1(92589) <= 16360142;
srom_1(92590) <= 16162679;
srom_1(92591) <= 15928760;
srom_1(92592) <= 15659484;
srom_1(92593) <= 15356112;
srom_1(92594) <= 15020066;
srom_1(92595) <= 14652924;
srom_1(92596) <= 14256406;
srom_1(92597) <= 13832372;
srom_1(92598) <= 13382810;
srom_1(92599) <= 12909828;
srom_1(92600) <= 12415645;
srom_1(92601) <= 11902578;
srom_1(92602) <= 11373033;
srom_1(92603) <= 10829493;
srom_1(92604) <= 10274506;
srom_1(92605) <= 9710676;
srom_1(92606) <= 9140646;
srom_1(92607) <= 8567090;
srom_1(92608) <= 7992697;
srom_1(92609) <= 7420160;
srom_1(92610) <= 6852165;
srom_1(92611) <= 6291374;
srom_1(92612) <= 5740418;
srom_1(92613) <= 5201881;
srom_1(92614) <= 4678287;
srom_1(92615) <= 4172092;
srom_1(92616) <= 3685670;
srom_1(92617) <= 3221301;
srom_1(92618) <= 2781164;
srom_1(92619) <= 2367322;
srom_1(92620) <= 1981716;
srom_1(92621) <= 1626154;
srom_1(92622) <= 1302303;
srom_1(92623) <= 1011682;
srom_1(92624) <= 755655;
srom_1(92625) <= 535421;
srom_1(92626) <= 352013;
srom_1(92627) <= 206292;
srom_1(92628) <= 98940;
srom_1(92629) <= 30461;
srom_1(92630) <= 1177;
srom_1(92631) <= 11224;
srom_1(92632) <= 60556;
srom_1(92633) <= 148940;
srom_1(92634) <= 275964;
srom_1(92635) <= 441030;
srom_1(92636) <= 643365;
srom_1(92637) <= 882020;
srom_1(92638) <= 1155876;
srom_1(92639) <= 1463649;
srom_1(92640) <= 1803896;
srom_1(92641) <= 2175020;
srom_1(92642) <= 2575282;
srom_1(92643) <= 3002805;
srom_1(92644) <= 3455584;
srom_1(92645) <= 3931495;
srom_1(92646) <= 4428307;
srom_1(92647) <= 4943691;
srom_1(92648) <= 5475228;
srom_1(92649) <= 6020428;
srom_1(92650) <= 6576733;
srom_1(92651) <= 7141534;
srom_1(92652) <= 7712183;
srom_1(92653) <= 8286005;
srom_1(92654) <= 8860307;
srom_1(92655) <= 9432398;
srom_1(92656) <= 9999593;
srom_1(92657) <= 10559235;
srom_1(92658) <= 11108697;
srom_1(92659) <= 11645404;
srom_1(92660) <= 12166839;
srom_1(92661) <= 12670556;
srom_1(92662) <= 13154194;
srom_1(92663) <= 13615484;
srom_1(92664) <= 14052264;
srom_1(92665) <= 14462485;
srom_1(92666) <= 14844223;
srom_1(92667) <= 15195689;
srom_1(92668) <= 15515234;
srom_1(92669) <= 15801360;
srom_1(92670) <= 16052725;
srom_1(92671) <= 16268150;
srom_1(92672) <= 16446625;
srom_1(92673) <= 16587313;
srom_1(92674) <= 16689555;
srom_1(92675) <= 16752871;
srom_1(92676) <= 16776964;
srom_1(92677) <= 16761721;
srom_1(92678) <= 16707214;
srom_1(92679) <= 16613698;
srom_1(92680) <= 16481612;
srom_1(92681) <= 16311574;
srom_1(92682) <= 16104384;
srom_1(92683) <= 15861011;
srom_1(92684) <= 15582597;
srom_1(92685) <= 15270449;
srom_1(92686) <= 14926029;
srom_1(92687) <= 14550953;
srom_1(92688) <= 14146980;
srom_1(92689) <= 13716003;
srom_1(92690) <= 13260045;
srom_1(92691) <= 12781243;
srom_1(92692) <= 12281842;
srom_1(92693) <= 11764184;
srom_1(92694) <= 11230698;
srom_1(92695) <= 10683883;
srom_1(92696) <= 10126306;
srom_1(92697) <= 9560579;
srom_1(92698) <= 8989357;
srom_1(92699) <= 8415318;
srom_1(92700) <= 7841154;
srom_1(92701) <= 7269556;
srom_1(92702) <= 6703207;
srom_1(92703) <= 6144760;
srom_1(92704) <= 5596836;
srom_1(92705) <= 5062004;
srom_1(92706) <= 4542771;
srom_1(92707) <= 4041572;
srom_1(92708) <= 3560758;
srom_1(92709) <= 3102584;
srom_1(92710) <= 2669198;
srom_1(92711) <= 2262632;
srom_1(92712) <= 1884792;
srom_1(92713) <= 1537452;
srom_1(92714) <= 1222239;
srom_1(92715) <= 940631;
srom_1(92716) <= 693949;
srom_1(92717) <= 483351;
srom_1(92718) <= 309822;
srom_1(92719) <= 174178;
srom_1(92720) <= 77055;
srom_1(92721) <= 18907;
srom_1(92722) <= 7;
srom_1(92723) <= 20444;
srom_1(92724) <= 80123;
srom_1(92725) <= 178763;
srom_1(92726) <= 315902;
srom_1(92727) <= 490896;
srom_1(92728) <= 702926;
srom_1(92729) <= 950996;
srom_1(92730) <= 1233944;
srom_1(92731) <= 1550442;
srom_1(92732) <= 1899007;
srom_1(92733) <= 2278004;
srom_1(92734) <= 2685655;
srom_1(92735) <= 3120050;
srom_1(92736) <= 3579151;
srom_1(92737) <= 4060805;
srom_1(92738) <= 4562754;
srom_1(92739) <= 5082643;
srom_1(92740) <= 5618035;
srom_1(92741) <= 6166419;
srom_1(92742) <= 6725224;
srom_1(92743) <= 7291829;
srom_1(92744) <= 7863577;
srom_1(92745) <= 8437787;
srom_1(92746) <= 9011767;
srom_1(92747) <= 9582824;
srom_1(92748) <= 10148282;
srom_1(92749) <= 10705487;
srom_1(92750) <= 11251828;
srom_1(92751) <= 11784742;
srom_1(92752) <= 12301731;
srom_1(92753) <= 12800370;
srom_1(92754) <= 13278320;
srom_1(92755) <= 13733341;
srom_1(92756) <= 14163298;
srom_1(92757) <= 14566176;
srom_1(92758) <= 14940086;
srom_1(92759) <= 15283273;
srom_1(92760) <= 15594128;
srom_1(92761) <= 15871195;
srom_1(92762) <= 16113173;
srom_1(92763) <= 16318928;
srom_1(92764) <= 16487495;
srom_1(92765) <= 16618083;
srom_1(92766) <= 16710081;
srom_1(92767) <= 16763056;
srom_1(92768) <= 16776761;
srom_1(92769) <= 16751131;
srom_1(92770) <= 16686286;
srom_1(92771) <= 16582530;
srom_1(92772) <= 16440350;
srom_1(92773) <= 16260413;
srom_1(92774) <= 16043562;
srom_1(92775) <= 15790815;
srom_1(92776) <= 15503356;
srom_1(92777) <= 15182533;
srom_1(92778) <= 14829852;
srom_1(92779) <= 14446965;
srom_1(92780) <= 14035668;
srom_1(92781) <= 13597891;
srom_1(92782) <= 13135685;
srom_1(92783) <= 12651219;
srom_1(92784) <= 12146764;
srom_1(92785) <= 11624685;
srom_1(92786) <= 11087432;
srom_1(92787) <= 10537523;
srom_1(92788) <= 9977536;
srom_1(92789) <= 9410099;
srom_1(92790) <= 8837871;
srom_1(92791) <= 8263537;
srom_1(92792) <= 7689790;
srom_1(92793) <= 7119319;
srom_1(92794) <= 6554800;
srom_1(92795) <= 5998881;
srom_1(92796) <= 5454168;
srom_1(92797) <= 4923216;
srom_1(92798) <= 4408514;
srom_1(92799) <= 3912476;
srom_1(92800) <= 3437428;
srom_1(92801) <= 2985598;
srom_1(92802) <= 2559104;
srom_1(92803) <= 2159947;
srom_1(92804) <= 1789999;
srom_1(92805) <= 1450993;
srom_1(92806) <= 1144520;
srom_1(92807) <= 872018;
srom_1(92808) <= 634763;
srom_1(92809) <= 433869;
srom_1(92810) <= 270277;
srom_1(92811) <= 144754;
srom_1(92812) <= 57890;
srom_1(92813) <= 10092;
srom_1(92814) <= 1583;
srom_1(92815) <= 32404;
srom_1(92816) <= 102411;
srom_1(92817) <= 211273;
srom_1(92818) <= 358483;
srom_1(92819) <= 543348;
srom_1(92820) <= 765002;
srom_1(92821) <= 1022406;
srom_1(92822) <= 1314353;
srom_1(92823) <= 1639473;
srom_1(92824) <= 1996243;
srom_1(92825) <= 2382988;
srom_1(92826) <= 2797896;
srom_1(92827) <= 3239020;
srom_1(92828) <= 3704293;
srom_1(92829) <= 4191532;
srom_1(92830) <= 4698452;
srom_1(92831) <= 5222677;
srom_1(92832) <= 5761748;
srom_1(92833) <= 6313138;
srom_1(92834) <= 6874260;
srom_1(92835) <= 7442483;
srom_1(92836) <= 8015143;
srom_1(92837) <= 8589554;
srom_1(92838) <= 9163023;
srom_1(92839) <= 9732860;
srom_1(92840) <= 10296394;
srom_1(92841) <= 10850981;
srom_1(92842) <= 11394022;
srom_1(92843) <= 11922969;
srom_1(92844) <= 12435342;
srom_1(92845) <= 12928739;
srom_1(92846) <= 13400845;
srom_1(92847) <= 13849448;
srom_1(92848) <= 14272442;
srom_1(92849) <= 14667845;
srom_1(92850) <= 15033803;
srom_1(92851) <= 15368599;
srom_1(92852) <= 15670664;
srom_1(92853) <= 15938580;
srom_1(92854) <= 16171093;
srom_1(92855) <= 16367110;
srom_1(92856) <= 16525713;
srom_1(92857) <= 16646159;
srom_1(92858) <= 16727882;
srom_1(92859) <= 16770500;
srom_1(92860) <= 16773812;
srom_1(92861) <= 16737802;
srom_1(92862) <= 16662641;
srom_1(92863) <= 16548680;
srom_1(92864) <= 16396453;
srom_1(92865) <= 16206675;
srom_1(92866) <= 15980235;
srom_1(92867) <= 15718195;
srom_1(92868) <= 15421785;
srom_1(92869) <= 15092393;
srom_1(92870) <= 14731566;
srom_1(92871) <= 14340993;
srom_1(92872) <= 13922508;
srom_1(92873) <= 13478073;
srom_1(92874) <= 13009772;
srom_1(92875) <= 12519800;
srom_1(92876) <= 12010455;
srom_1(92877) <= 11484127;
srom_1(92878) <= 10943282;
srom_1(92879) <= 10390458;
srom_1(92880) <= 9828247;
srom_1(92881) <= 9259284;
srom_1(92882) <= 8686239;
srom_1(92883) <= 8111797;
srom_1(92884) <= 7538654;
srom_1(92885) <= 6969497;
srom_1(92886) <= 6406994;
srom_1(92887) <= 5853784;
srom_1(92888) <= 5312461;
srom_1(92889) <= 4785562;
srom_1(92890) <= 4275560;
srom_1(92891) <= 3784844;
srom_1(92892) <= 3315718;
srom_1(92893) <= 2870380;
srom_1(92894) <= 2450919;
srom_1(92895) <= 2059302;
srom_1(92896) <= 1697365;
srom_1(92897) <= 1366806;
srom_1(92898) <= 1069174;
srom_1(92899) <= 805865;
srom_1(92900) <= 578115;
srom_1(92901) <= 386991;
srom_1(92902) <= 233389;
srom_1(92903) <= 118029;
srom_1(92904) <= 41454;
srom_1(92905) <= 4021;
srom_1(92906) <= 5906;
srom_1(92907) <= 47100;
srom_1(92908) <= 127411;
srom_1(92909) <= 246461;
srom_1(92910) <= 403693;
srom_1(92911) <= 598368;
srom_1(92912) <= 829575;
srom_1(92913) <= 1096229;
srom_1(92914) <= 1397079;
srom_1(92915) <= 1730714;
srom_1(92916) <= 2095571;
srom_1(92917) <= 2489938;
srom_1(92918) <= 2911966;
srom_1(92919) <= 3359676;
srom_1(92920) <= 3830968;
srom_1(92921) <= 4323633;
srom_1(92922) <= 4835359;
srom_1(92923) <= 5363748;
srom_1(92924) <= 5906322;
srom_1(92925) <= 6460536;
srom_1(92926) <= 7023791;
srom_1(92927) <= 7593446;
srom_1(92928) <= 8166830;
srom_1(92929) <= 8741255;
srom_1(92930) <= 9314025;
srom_1(92931) <= 9882456;
srom_1(92932) <= 10443881;
srom_1(92933) <= 10995669;
srom_1(92934) <= 11535231;
srom_1(92935) <= 12060038;
srom_1(92936) <= 12567628;
srom_1(92937) <= 13055621;
srom_1(92938) <= 13521730;
srom_1(92939) <= 13963767;
srom_1(92940) <= 14379660;
srom_1(92941) <= 14767459;
srom_1(92942) <= 15125345;
srom_1(92943) <= 15451641;
srom_1(92944) <= 15744815;
srom_1(92945) <= 16003494;
srom_1(92946) <= 16226464;
srom_1(92947) <= 16412680;
srom_1(92948) <= 16561268;
srom_1(92949) <= 16671531;
srom_1(92950) <= 16742953;
srom_1(92951) <= 16775199;
srom_1(92952) <= 16768117;
srom_1(92953) <= 16721740;
srom_1(92954) <= 16636287;
srom_1(92955) <= 16512158;
srom_1(92956) <= 16349934;
srom_1(92957) <= 16150377;
srom_1(92958) <= 15914422;
srom_1(92959) <= 15643176;
srom_1(92960) <= 15337911;
srom_1(92961) <= 15000059;
srom_1(92962) <= 14631203;
srom_1(92963) <= 14233073;
srom_1(92964) <= 13807537;
srom_1(92965) <= 13356589;
srom_1(92966) <= 12882345;
srom_1(92967) <= 12387028;
srom_1(92968) <= 11872961;
srom_1(92969) <= 11342555;
srom_1(92970) <= 10798297;
srom_1(92971) <= 10242738;
srom_1(92972) <= 9678486;
srom_1(92973) <= 9108184;
srom_1(92974) <= 8534508;
srom_1(92975) <= 7960148;
srom_1(92976) <= 7387797;
srom_1(92977) <= 6820140;
srom_1(92978) <= 6259837;
srom_1(92979) <= 5709517;
srom_1(92980) <= 5171760;
srom_1(92981) <= 4649088;
srom_1(92982) <= 4143952;
srom_1(92983) <= 3658721;
srom_1(92984) <= 3195669;
srom_1(92985) <= 2756969;
srom_1(92986) <= 2344678;
srom_1(92987) <= 1960729;
srom_1(92988) <= 1606922;
srom_1(92989) <= 1284917;
srom_1(92990) <= 996224;
srom_1(92991) <= 742196;
srom_1(92992) <= 524024;
srom_1(92993) <= 342733;
srom_1(92994) <= 199171;
srom_1(92995) <= 94012;
srom_1(92996) <= 27750;
srom_1(92997) <= 694;
srom_1(92998) <= 12973;
srom_1(92999) <= 64527;
srom_1(93000) <= 155116;
srom_1(93001) <= 284315;
srom_1(93002) <= 451517;
srom_1(93003) <= 655939;
srom_1(93004) <= 896623;
srom_1(93005) <= 1172438;
srom_1(93006) <= 1482093;
srom_1(93007) <= 1824135;
srom_1(93008) <= 2196960;
srom_1(93009) <= 2598820;
srom_1(93010) <= 3027830;
srom_1(93011) <= 3481978;
srom_1(93012) <= 3959136;
srom_1(93013) <= 4457065;
srom_1(93014) <= 4973430;
srom_1(93015) <= 5505810;
srom_1(93016) <= 6051708;
srom_1(93017) <= 6608565;
srom_1(93018) <= 7173769;
srom_1(93019) <= 7744670;
srom_1(93020) <= 8318591;
srom_1(93021) <= 8892840;
srom_1(93022) <= 9464724;
srom_1(93023) <= 10031562;
srom_1(93024) <= 10590696;
srom_1(93025) <= 11139503;
srom_1(93026) <= 11675411;
srom_1(93027) <= 12195905;
srom_1(93028) <= 12698546;
srom_1(93029) <= 13180976;
srom_1(93030) <= 13640933;
srom_1(93031) <= 14076260;
srom_1(93032) <= 14484916;
srom_1(93033) <= 14864984;
srom_1(93034) <= 15214682;
srom_1(93035) <= 15532370;
srom_1(93036) <= 15816558;
srom_1(93037) <= 16065915;
srom_1(93038) <= 16279270;
srom_1(93039) <= 16455623;
srom_1(93040) <= 16594146;
srom_1(93041) <= 16694192;
srom_1(93042) <= 16755289;
srom_1(93043) <= 16777152;
srom_1(93044) <= 16759679;
srom_1(93045) <= 16702950;
srom_1(93046) <= 16607233;
srom_1(93047) <= 16472976;
srom_1(93048) <= 16300808;
srom_1(93049) <= 16091538;
srom_1(93050) <= 15846145;
srom_1(93051) <= 15565782;
srom_1(93052) <= 15251763;
srom_1(93053) <= 14905560;
srom_1(93054) <= 14528796;
srom_1(93055) <= 14123239;
srom_1(93056) <= 13690791;
srom_1(93057) <= 13233478;
srom_1(93058) <= 12753447;
srom_1(93059) <= 12252947;
srom_1(93060) <= 11734326;
srom_1(93061) <= 11200016;
srom_1(93062) <= 10652522;
srom_1(93063) <= 10094412;
srom_1(93064) <= 9528302;
srom_1(93065) <= 8956849;
srom_1(93066) <= 8382730;
srom_1(93067) <= 7808639;
srom_1(93068) <= 7237268;
srom_1(93069) <= 6671296;
srom_1(93070) <= 6113377;
srom_1(93071) <= 5566127;
srom_1(93072) <= 5032113;
srom_1(93073) <= 4513839;
srom_1(93074) <= 4013734;
srom_1(93075) <= 3534145;
srom_1(93076) <= 3077320;
srom_1(93077) <= 2645402;
srom_1(93078) <= 2240415;
srom_1(93079) <= 1864260;
srom_1(93080) <= 1518699;
srom_1(93081) <= 1205354;
srom_1(93082) <= 925693;
srom_1(93083) <= 681029;
srom_1(93084) <= 472508;
srom_1(93085) <= 301109;
srom_1(93086) <= 167634;
srom_1(93087) <= 72711;
srom_1(93088) <= 16783;
srom_1(93089) <= 114;
srom_1(93090) <= 22781;
srom_1(93091) <= 84679;
srom_1(93092) <= 185517;
srom_1(93093) <= 324821;
srom_1(93094) <= 501940;
srom_1(93095) <= 716042;
srom_1(93096) <= 966123;
srom_1(93097) <= 1251011;
srom_1(93098) <= 1569369;
srom_1(93099) <= 1919705;
srom_1(93100) <= 2300376;
srom_1(93101) <= 2709597;
srom_1(93102) <= 3145449;
srom_1(93103) <= 3605887;
srom_1(93104) <= 4088754;
srom_1(93105) <= 4591784;
srom_1(93106) <= 5112618;
srom_1(93107) <= 5648815;
srom_1(93108) <= 6197859;
srom_1(93109) <= 6757177;
srom_1(93110) <= 7324145;
srom_1(93111) <= 7896105;
srom_1(93112) <= 8470374;
srom_1(93113) <= 9044260;
srom_1(93114) <= 9615071;
srom_1(93115) <= 10180131;
srom_1(93116) <= 10736790;
srom_1(93117) <= 11282437;
srom_1(93118) <= 11814514;
srom_1(93119) <= 12330526;
srom_1(93120) <= 12828053;
srom_1(93121) <= 13304762;
srom_1(93122) <= 13758417;
srom_1(93123) <= 14186892;
srom_1(93124) <= 14588176;
srom_1(93125) <= 14960388;
srom_1(93126) <= 15301783;
srom_1(93127) <= 15610760;
srom_1(93128) <= 15885870;
srom_1(93129) <= 16125822;
srom_1(93130) <= 16329492;
srom_1(93131) <= 16495924;
srom_1(93132) <= 16624339;
srom_1(93133) <= 16714133;
srom_1(93134) <= 16764886;
srom_1(93135) <= 16776359;
srom_1(93136) <= 16748500;
srom_1(93137) <= 16681438;
srom_1(93138) <= 16575488;
srom_1(93139) <= 16431147;
srom_1(93140) <= 16249092;
srom_1(93141) <= 16030177;
srom_1(93142) <= 15775427;
srom_1(93143) <= 15486038;
srom_1(93144) <= 15163367;
srom_1(93145) <= 14808927;
srom_1(93146) <= 14424379;
srom_1(93147) <= 14011528;
srom_1(93148) <= 13572309;
srom_1(93149) <= 13108782;
srom_1(93150) <= 12623120;
srom_1(93151) <= 12117601;
srom_1(93152) <= 11594596;
srom_1(93153) <= 11056556;
srom_1(93154) <= 10506006;
srom_1(93155) <= 9945526;
srom_1(93156) <= 9377746;
srom_1(93157) <= 8805327;
srom_1(93158) <= 8230954;
srom_1(93159) <= 7657320;
srom_1(93160) <= 7087116;
srom_1(93161) <= 6523015;
srom_1(93162) <= 5967662;
srom_1(93163) <= 5423661;
srom_1(93164) <= 4893565;
srom_1(93165) <= 4379857;
srom_1(93166) <= 3884949;
srom_1(93167) <= 3411159;
srom_1(93168) <= 2960710;
srom_1(93169) <= 2535715;
srom_1(93170) <= 2138166;
srom_1(93171) <= 1769927;
srom_1(93172) <= 1432726;
srom_1(93173) <= 1128143;
srom_1(93174) <= 857607;
srom_1(93175) <= 622386;
srom_1(93176) <= 423584;
srom_1(93177) <= 262132;
srom_1(93178) <= 138789;
srom_1(93179) <= 54131;
srom_1(93180) <= 8557;
srom_1(93181) <= 2280;
srom_1(93182) <= 35329;
srom_1(93183) <= 107550;
srom_1(93184) <= 218603;
srom_1(93185) <= 367968;
srom_1(93186) <= 554945;
srom_1(93187) <= 778656;
srom_1(93188) <= 1038053;
srom_1(93189) <= 1331920;
srom_1(93190) <= 1658877;
srom_1(93191) <= 2017393;
srom_1(93192) <= 2405785;
srom_1(93193) <= 2822233;
srom_1(93194) <= 3264784;
srom_1(93195) <= 3731362;
srom_1(93196) <= 4219779;
srom_1(93197) <= 4727746;
srom_1(93198) <= 5252879;
srom_1(93199) <= 5792717;
srom_1(93200) <= 6344728;
srom_1(93201) <= 6906323;
srom_1(93202) <= 7474870;
srom_1(93203) <= 8047701;
srom_1(93204) <= 8622131;
srom_1(93205) <= 9195465;
srom_1(93206) <= 9765017;
srom_1(93207) <= 10328113;
srom_1(93208) <= 10882115;
srom_1(93209) <= 11424424;
srom_1(93210) <= 11952496;
srom_1(93211) <= 12463857;
srom_1(93212) <= 12956107;
srom_1(93213) <= 13426938;
srom_1(93214) <= 13874144;
srom_1(93215) <= 14295625;
srom_1(93216) <= 14689407;
srom_1(93217) <= 15053641;
srom_1(93218) <= 15386622;
srom_1(93219) <= 15686786;
srom_1(93220) <= 15952726;
srom_1(93221) <= 16183196;
srom_1(93222) <= 16377114;
srom_1(93223) <= 16533572;
srom_1(93224) <= 16651834;
srom_1(93225) <= 16731348;
srom_1(93226) <= 16771740;
srom_1(93227) <= 16772820;
srom_1(93228) <= 16734584;
srom_1(93229) <= 16657211;
srom_1(93230) <= 16541063;
srom_1(93231) <= 16386686;
srom_1(93232) <= 16194803;
srom_1(93233) <= 15966314;
srom_1(93234) <= 15702291;
srom_1(93235) <= 15403971;
srom_1(93236) <= 15072753;
srom_1(93237) <= 14710192;
srom_1(93238) <= 14317986;
srom_1(93239) <= 13897976;
srom_1(93240) <= 13452130;
srom_1(93241) <= 12982540;
srom_1(93242) <= 12491407;
srom_1(93243) <= 11981034;
srom_1(93244) <= 11453816;
srom_1(93245) <= 10912223;
srom_1(93246) <= 10358797;
srom_1(93247) <= 9796131;
srom_1(93248) <= 9226866;
srom_1(93249) <= 8653669;
srom_1(93250) <= 8079230;
srom_1(93251) <= 7506241;
srom_1(93252) <= 6937390;
srom_1(93253) <= 6375344;
srom_1(93254) <= 5822739;
srom_1(93255) <= 5282166;
srom_1(93256) <= 4756161;
srom_1(93257) <= 4247189;
srom_1(93258) <= 3757638;
srom_1(93259) <= 3289803;
srom_1(93260) <= 2845878;
srom_1(93261) <= 2427944;
srom_1(93262) <= 2037963;
srom_1(93263) <= 1677761;
srom_1(93264) <= 1349030;
srom_1(93265) <= 1053309;
srom_1(93266) <= 791986;
srom_1(93267) <= 566286;
srom_1(93268) <= 377267;
srom_1(93269) <= 225817;
srom_1(93270) <= 112645;
srom_1(93271) <= 38281;
srom_1(93272) <= 3075;
srom_1(93273) <= 7192;
srom_1(93274) <= 50612;
srom_1(93275) <= 133131;
srom_1(93276) <= 254364;
srom_1(93277) <= 413741;
srom_1(93278) <= 610514;
srom_1(93279) <= 843762;
srom_1(93280) <= 1112390;
srom_1(93281) <= 1415139;
srom_1(93282) <= 1750589;
srom_1(93283) <= 2117167;
srom_1(93284) <= 2513153;
srom_1(93285) <= 2936692;
srom_1(93286) <= 3385797;
srom_1(93287) <= 3858361;
srom_1(93288) <= 4352169;
srom_1(93289) <= 4864906;
srom_1(93290) <= 5394167;
srom_1(93291) <= 5937469;
srom_1(93292) <= 6492266;
srom_1(93293) <= 7055955;
srom_1(93294) <= 7625893;
srom_1(93295) <= 8199408;
srom_1(93296) <= 8773811;
srom_1(93297) <= 9346407;
srom_1(93298) <= 9914511;
srom_1(93299) <= 10475460;
srom_1(93300) <= 11026623;
srom_1(93301) <= 11565416;
srom_1(93302) <= 12089311;
srom_1(93303) <= 12595853;
srom_1(93304) <= 13082665;
srom_1(93305) <= 13547465;
srom_1(93306) <= 13988074;
srom_1(93307) <= 14402424;
srom_1(93308) <= 14788574;
srom_1(93309) <= 15144712;
srom_1(93310) <= 15469169;
srom_1(93311) <= 15760422;
srom_1(93312) <= 16017107;
srom_1(93313) <= 16238018;
srom_1(93314) <= 16422121;
srom_1(93315) <= 16568553;
srom_1(93316) <= 16676625;
srom_1(93317) <= 16745832;
srom_1(93318) <= 16775850;
srom_1(93319) <= 16766536;
srom_1(93320) <= 16717936;
srom_1(93321) <= 16630277;
srom_1(93322) <= 16503969;
srom_1(93323) <= 16339606;
srom_1(93324) <= 16137958;
srom_1(93325) <= 15899970;
srom_1(93326) <= 15626759;
srom_1(93327) <= 15319606;
srom_1(93328) <= 14979952;
srom_1(93329) <= 14609388;
srom_1(93330) <= 14209652;
srom_1(93331) <= 13782620;
srom_1(93332) <= 13330293;
srom_1(93333) <= 12854793;
srom_1(93334) <= 12358350;
srom_1(93335) <= 11843291;
srom_1(93336) <= 11312032;
srom_1(93337) <= 10767064;
srom_1(93338) <= 10210943;
srom_1(93339) <= 9646276;
srom_1(93340) <= 9075711;
srom_1(93341) <= 8501924;
srom_1(93342) <= 7927606;
srom_1(93343) <= 7355450;
srom_1(93344) <= 6788139;
srom_1(93345) <= 6228332;
srom_1(93346) <= 5678656;
srom_1(93347) <= 5141688;
srom_1(93348) <= 4619946;
srom_1(93349) <= 4115876;
srom_1(93350) <= 3631843;
srom_1(93351) <= 3170115;
srom_1(93352) <= 2732859;
srom_1(93353) <= 2322125;
srom_1(93354) <= 1939839;
srom_1(93355) <= 1587793;
srom_1(93356) <= 1267638;
srom_1(93357) <= 980876;
srom_1(93358) <= 728852;
srom_1(93359) <= 512746;
srom_1(93360) <= 333574;
srom_1(93361) <= 192174;
srom_1(93362) <= 89210;
srom_1(93363) <= 25164;
srom_1(93364) <= 338;
srom_1(93365) <= 14847;
srom_1(93366) <= 68624;
srom_1(93367) <= 161416;
srom_1(93368) <= 292788;
srom_1(93369) <= 462124;
srom_1(93370) <= 668630;
srom_1(93371) <= 911338;
srom_1(93372) <= 1189109;
srom_1(93373) <= 1500641;
srom_1(93374) <= 1844474;
srom_1(93375) <= 2218993;
srom_1(93376) <= 2622445;
srom_1(93377) <= 3052936;
srom_1(93378) <= 3508447;
srom_1(93379) <= 3986844;
srom_1(93380) <= 4485881;
srom_1(93381) <= 5003220;
srom_1(93382) <= 5536434;
srom_1(93383) <= 6083023;
srom_1(93384) <= 6640424;
srom_1(93385) <= 7206023;
srom_1(93386) <= 7777167;
srom_1(93387) <= 8351178;
srom_1(93388) <= 8925365;
srom_1(93389) <= 9497035;
srom_1(93390) <= 10063507;
srom_1(93391) <= 10622124;
srom_1(93392) <= 11170268;
srom_1(93393) <= 11705368;
srom_1(93394) <= 12224915;
srom_1(93395) <= 12726471;
srom_1(93396) <= 13207686;
srom_1(93397) <= 13666303;
srom_1(93398) <= 14100171;
srom_1(93399) <= 14507255;
srom_1(93400) <= 14885647;
srom_1(93401) <= 15233572;
srom_1(93402) <= 15549398;
srom_1(93403) <= 15831645;
srom_1(93404) <= 16078989;
srom_1(93405) <= 16290271;
srom_1(93406) <= 16464498;
srom_1(93407) <= 16600855;
srom_1(93408) <= 16698702;
srom_1(93409) <= 16757580;
srom_1(93410) <= 16777213;
srom_1(93411) <= 16757510;
srom_1(93412) <= 16698561;
srom_1(93413) <= 16600644;
srom_1(93414) <= 16464218;
srom_1(93415) <= 16289923;
srom_1(93416) <= 16078576;
srom_1(93417) <= 15831168;
srom_1(93418) <= 15548859;
srom_1(93419) <= 15232973;
srom_1(93420) <= 14884992;
srom_1(93421) <= 14506546;
srom_1(93422) <= 14099412;
srom_1(93423) <= 13665498;
srom_1(93424) <= 13206839;
srom_1(93425) <= 12725585;
srom_1(93426) <= 12223994;
srom_1(93427) <= 11704417;
srom_1(93428) <= 11169292;
srom_1(93429) <= 10621126;
srom_1(93430) <= 10062492;
srom_1(93431) <= 9496008;
srom_1(93432) <= 8924331;
srom_1(93433) <= 8350143;
srom_1(93434) <= 7776134;
srom_1(93435) <= 7204998;
srom_1(93436) <= 6639411;
srom_1(93437) <= 6082028;
srom_1(93438) <= 5535461;
srom_1(93439) <= 5002273;
srom_1(93440) <= 4484965;
srom_1(93441) <= 3985962;
srom_1(93442) <= 3507605;
srom_1(93443) <= 3052137;
srom_1(93444) <= 2621693;
srom_1(93445) <= 2218292;
srom_1(93446) <= 1843826;
srom_1(93447) <= 1500050;
srom_1(93448) <= 1188578;
srom_1(93449) <= 910869;
srom_1(93450) <= 668225;
srom_1(93451) <= 461785;
srom_1(93452) <= 292517;
srom_1(93453) <= 161214;
srom_1(93454) <= 68492;
srom_1(93455) <= 14786;
srom_1(93456) <= 348;
srom_1(93457) <= 25245;
srom_1(93458) <= 89360;
srom_1(93459) <= 192394;
srom_1(93460) <= 333863;
srom_1(93461) <= 513103;
srom_1(93462) <= 729274;
srom_1(93463) <= 981362;
srom_1(93464) <= 1268185;
srom_1(93465) <= 1588399;
srom_1(93466) <= 1940501;
srom_1(93467) <= 2322840;
srom_1(93468) <= 2733624;
srom_1(93469) <= 3170926;
srom_1(93470) <= 3632696;
srom_1(93471) <= 4116767;
srom_1(93472) <= 4620871;
srom_1(93473) <= 5142643;
srom_1(93474) <= 5679636;
srom_1(93475) <= 6229333;
srom_1(93476) <= 6789155;
srom_1(93477) <= 7356478;
srom_1(93478) <= 7928640;
srom_1(93479) <= 8502960;
srom_1(93480) <= 9076743;
srom_1(93481) <= 9647299;
srom_1(93482) <= 10211953;
srom_1(93483) <= 10768057;
srom_1(93484) <= 11313003;
srom_1(93485) <= 11844235;
srom_1(93486) <= 12359262;
srom_1(93487) <= 12855670;
srom_1(93488) <= 13331130;
srom_1(93489) <= 13783413;
srom_1(93490) <= 14210398;
srom_1(93491) <= 14610082;
srom_1(93492) <= 14980592;
srom_1(93493) <= 15320190;
srom_1(93494) <= 15627283;
srom_1(93495) <= 15900431;
srom_1(93496) <= 16138354;
srom_1(93497) <= 16339936;
srom_1(93498) <= 16504231;
srom_1(93499) <= 16630469;
srom_1(93500) <= 16718059;
srom_1(93501) <= 16766588;
srom_1(93502) <= 16775831;
srom_1(93503) <= 16745743;
srom_1(93504) <= 16676465;
srom_1(93505) <= 16568323;
srom_1(93506) <= 16421823;
srom_1(93507) <= 16237653;
srom_1(93508) <= 16016676;
srom_1(93509) <= 15759928;
srom_1(93510) <= 15468614;
srom_1(93511) <= 15144099;
srom_1(93512) <= 14787905;
srom_1(93513) <= 14401702;
srom_1(93514) <= 13987303;
srom_1(93515) <= 13546649;
srom_1(93516) <= 13081807;
srom_1(93517) <= 12594957;
srom_1(93518) <= 12088382;
srom_1(93519) <= 11564458;
srom_1(93520) <= 11025641;
srom_1(93521) <= 10474457;
srom_1(93522) <= 9913493;
srom_1(93523) <= 9345378;
srom_1(93524) <= 8772776;
srom_1(93525) <= 8198373;
srom_1(93526) <= 7624862;
srom_1(93527) <= 7054933;
srom_1(93528) <= 6491257;
srom_1(93529) <= 5936479;
srom_1(93530) <= 5393199;
srom_1(93531) <= 4863966;
srom_1(93532) <= 4351262;
srom_1(93533) <= 3857490;
srom_1(93534) <= 3384965;
srom_1(93535) <= 2935905;
srom_1(93536) <= 2512414;
srom_1(93537) <= 2116479;
srom_1(93538) <= 1749956;
srom_1(93539) <= 1414564;
srom_1(93540) <= 1111875;
srom_1(93541) <= 843310;
srom_1(93542) <= 610127;
srom_1(93543) <= 413420;
srom_1(93544) <= 254111;
srom_1(93545) <= 132948;
srom_1(93546) <= 50498;
srom_1(93547) <= 7149;
srom_1(93548) <= 3103;
srom_1(93549) <= 38380;
srom_1(93550) <= 112814;
srom_1(93551) <= 226056;
srom_1(93552) <= 377574;
srom_1(93553) <= 566660;
srom_1(93554) <= 792425;
srom_1(93555) <= 1053811;
srom_1(93556) <= 1349593;
srom_1(93557) <= 1678383;
srom_1(93558) <= 2038639;
srom_1(93559) <= 2428673;
srom_1(93560) <= 2846655;
srom_1(93561) <= 3290625;
srom_1(93562) <= 3758501;
srom_1(93563) <= 4248089;
srom_1(93564) <= 4757094;
srom_1(93565) <= 5283128;
srom_1(93566) <= 5823725;
srom_1(93567) <= 6376349;
srom_1(93568) <= 6938410;
srom_1(93569) <= 7507270;
srom_1(93570) <= 8080264;
srom_1(93571) <= 8654704;
srom_1(93572) <= 9227896;
srom_1(93573) <= 9797152;
srom_1(93574) <= 10359803;
srom_1(93575) <= 10913211;
srom_1(93576) <= 11454779;
srom_1(93577) <= 11981970;
srom_1(93578) <= 12492310;
srom_1(93579) <= 12983406;
srom_1(93580) <= 13452955;
srom_1(93581) <= 13898757;
srom_1(93582) <= 14318719;
srom_1(93583) <= 14710873;
srom_1(93584) <= 15073379;
srom_1(93585) <= 15404538;
srom_1(93586) <= 15702798;
srom_1(93587) <= 15966758;
srom_1(93588) <= 16195182;
srom_1(93589) <= 16386998;
srom_1(93590) <= 16541307;
srom_1(93591) <= 16657385;
srom_1(93592) <= 16734688;
srom_1(93593) <= 16772854;
srom_1(93594) <= 16771702;
srom_1(93595) <= 16731240;
srom_1(93596) <= 16651656;
srom_1(93597) <= 16533324;
srom_1(93598) <= 16376798;
srom_1(93599) <= 16182813;
srom_1(93600) <= 15952279;
srom_1(93601) <= 15686275;
srom_1(93602) <= 15386051;
srom_1(93603) <= 15053013;
srom_1(93604) <= 14688723;
srom_1(93605) <= 14294890;
srom_1(93606) <= 13873360;
srom_1(93607) <= 13426110;
srom_1(93608) <= 12955238;
srom_1(93609) <= 12462952;
srom_1(93610) <= 11951559;
srom_1(93611) <= 11423458;
srom_1(93612) <= 10881126;
srom_1(93613) <= 10327106;
srom_1(93614) <= 9763995;
srom_1(93615) <= 9194435;
srom_1(93616) <= 8621096;
srom_1(93617) <= 8046666;
srom_1(93618) <= 7473840;
srom_1(93619) <= 6905304;
srom_1(93620) <= 6343724;
srom_1(93621) <= 5791732;
srom_1(93622) <= 5251919;
srom_1(93623) <= 4726814;
srom_1(93624) <= 4218881;
srom_1(93625) <= 3730501;
srom_1(93626) <= 3263964;
srom_1(93627) <= 2821459;
srom_1(93628) <= 2405060;
srom_1(93629) <= 2016719;
srom_1(93630) <= 1658259;
srom_1(93631) <= 1331360;
srom_1(93632) <= 1037554;
srom_1(93633) <= 778221;
srom_1(93634) <= 554574;
srom_1(93635) <= 367665;
srom_1(93636) <= 218368;
srom_1(93637) <= 107384;
srom_1(93638) <= 35234;
srom_1(93639) <= 2256;
srom_1(93640) <= 8604;
srom_1(93641) <= 54249;
srom_1(93642) <= 138976;
srom_1(93643) <= 262389;
srom_1(93644) <= 423909;
srom_1(93645) <= 622778;
srom_1(93646) <= 858063;
srom_1(93647) <= 1128662;
srom_1(93648) <= 1433305;
srom_1(93649) <= 1770563;
srom_1(93650) <= 2138857;
srom_1(93651) <= 2536457;
srom_1(93652) <= 2961500;
srom_1(93653) <= 3411993;
srom_1(93654) <= 3885822;
srom_1(93655) <= 4380767;
srom_1(93656) <= 4894506;
srom_1(93657) <= 5424630;
srom_1(93658) <= 5968653;
srom_1(93659) <= 6524024;
srom_1(93660) <= 7088139;
srom_1(93661) <= 7658352;
srom_1(93662) <= 8231989;
srom_1(93663) <= 8806361;
srom_1(93664) <= 9378774;
srom_1(93665) <= 9946544;
srom_1(93666) <= 10507008;
srom_1(93667) <= 11057538;
srom_1(93668) <= 11595552;
srom_1(93669) <= 12118529;
srom_1(93670) <= 12624014;
srom_1(93671) <= 13109638;
srom_1(93672) <= 13573123;
srom_1(93673) <= 14012296;
srom_1(93674) <= 14425098;
srom_1(93675) <= 14809593;
srom_1(93676) <= 15163978;
srom_1(93677) <= 15486590;
srom_1(93678) <= 15775918;
srom_1(93679) <= 16030604;
srom_1(93680) <= 16249454;
srom_1(93681) <= 16431442;
srom_1(93682) <= 16575714;
srom_1(93683) <= 16681594;
srom_1(93684) <= 16748585;
srom_1(93685) <= 16776374;
srom_1(93686) <= 16764829;
srom_1(93687) <= 16714006;
srom_1(93688) <= 16624142;
srom_1(93689) <= 16495658;
srom_1(93690) <= 16329158;
srom_1(93691) <= 16125422;
srom_1(93692) <= 15885405;
srom_1(93693) <= 15610233;
srom_1(93694) <= 15301197;
srom_1(93695) <= 14959745;
srom_1(93696) <= 14587478;
srom_1(93697) <= 14186143;
srom_1(93698) <= 13757622;
srom_1(93699) <= 13303923;
srom_1(93700) <= 12827175;
srom_1(93701) <= 12329612;
srom_1(93702) <= 11813569;
srom_1(93703) <= 11281465;
srom_1(93704) <= 10735796;
srom_1(93705) <= 10179119;
srom_1(93706) <= 9614047;
srom_1(93707) <= 9043228;
srom_1(93708) <= 8469339;
srom_1(93709) <= 7895071;
srom_1(93710) <= 7323118;
srom_1(93711) <= 6756162;
srom_1(93712) <= 6196860;
srom_1(93713) <= 5647836;
srom_1(93714) <= 5111665;
srom_1(93715) <= 4590860;
srom_1(93716) <= 4087865;
srom_1(93717) <= 3605037;
srom_1(93718) <= 3144640;
srom_1(93719) <= 2708835;
srom_1(93720) <= 2299664;
srom_1(93721) <= 1919046;
srom_1(93722) <= 1568766;
srom_1(93723) <= 1250467;
srom_1(93724) <= 965641;
srom_1(93725) <= 715623;
srom_1(93726) <= 501587;
srom_1(93727) <= 324536;
srom_1(93728) <= 185300;
srom_1(93729) <= 84532;
srom_1(93730) <= 22705;
srom_1(93731) <= 109;
srom_1(93732) <= 16849;
srom_1(93733) <= 72847;
srom_1(93734) <= 167840;
srom_1(93735) <= 301384;
srom_1(93736) <= 472851;
srom_1(93737) <= 681438;
srom_1(93738) <= 926166;
srom_1(93739) <= 1205889;
srom_1(93740) <= 1519294;
srom_1(93741) <= 1864911;
srom_1(93742) <= 2241120;
srom_1(93743) <= 2646157;
srom_1(93744) <= 3078122;
srom_1(93745) <= 3534990;
srom_1(93746) <= 4014618;
srom_1(93747) <= 4514757;
srom_1(93748) <= 5033062;
srom_1(93749) <= 5567102;
srom_1(93750) <= 6114374;
srom_1(93751) <= 6672310;
srom_1(93752) <= 7238294;
srom_1(93753) <= 7809672;
srom_1(93754) <= 8383766;
srom_1(93755) <= 8957882;
srom_1(93756) <= 9529328;
srom_1(93757) <= 10095425;
srom_1(93758) <= 10653519;
srom_1(93759) <= 11200991;
srom_1(93760) <= 11735276;
srom_1(93761) <= 12253866;
srom_1(93762) <= 12754331;
srom_1(93763) <= 13234324;
srom_1(93764) <= 13691593;
srom_1(93765) <= 14123995;
srom_1(93766) <= 14529502;
srom_1(93767) <= 14906211;
srom_1(93768) <= 15252358;
srom_1(93769) <= 15566318;
srom_1(93770) <= 15846620;
srom_1(93771) <= 16091948;
srom_1(93772) <= 16301152;
srom_1(93773) <= 16473252;
srom_1(93774) <= 16607440;
srom_1(93775) <= 16703088;
srom_1(93776) <= 16759745;
srom_1(93777) <= 16777148;
srom_1(93778) <= 16755214;
srom_1(93779) <= 16694046;
srom_1(93780) <= 16593931;
srom_1(93781) <= 16455338;
srom_1(93782) <= 16278918;
srom_1(93783) <= 16065498;
srom_1(93784) <= 15816077;
srom_1(93785) <= 15531827;
srom_1(93786) <= 15214080;
srom_1(93787) <= 14864326;
srom_1(93788) <= 14484205;
srom_1(93789) <= 14075499;
srom_1(93790) <= 13640126;
srom_1(93791) <= 13180126;
srom_1(93792) <= 12697658;
srom_1(93793) <= 12194983;
srom_1(93794) <= 11674458;
srom_1(93795) <= 11138525;
srom_1(93796) <= 10589697;
srom_1(93797) <= 10030547;
srom_1(93798) <= 9463697;
srom_1(93799) <= 8891806;
srom_1(93800) <= 8317555;
srom_1(93801) <= 7743638;
srom_1(93802) <= 7172745;
srom_1(93803) <= 6607553;
srom_1(93804) <= 6050714;
srom_1(93805) <= 5504837;
srom_1(93806) <= 4972484;
srom_1(93807) <= 4456150;
srom_1(93808) <= 3958257;
srom_1(93809) <= 3481139;
srom_1(93810) <= 3027034;
srom_1(93811) <= 2598071;
srom_1(93812) <= 2196262;
srom_1(93813) <= 1823491;
srom_1(93814) <= 1481506;
srom_1(93815) <= 1171910;
srom_1(93816) <= 896157;
srom_1(93817) <= 655538;
srom_1(93818) <= 451182;
srom_1(93819) <= 284047;
srom_1(93820) <= 154918;
srom_1(93821) <= 64399;
srom_1(93822) <= 12915;
srom_1(93823) <= 708;
srom_1(93824) <= 27834;
srom_1(93825) <= 94167;
srom_1(93826) <= 199395;
srom_1(93827) <= 343026;
srom_1(93828) <= 524385;
srom_1(93829) <= 742621;
srom_1(93830) <= 996713;
srom_1(93831) <= 1285468;
srom_1(93832) <= 1607531;
srom_1(93833) <= 1961394;
srom_1(93834) <= 2345396;
srom_1(93835) <= 2757737;
srom_1(93836) <= 3196482;
srom_1(93837) <= 3659576;
srom_1(93838) <= 4144845;
srom_1(93839) <= 4650015;
srom_1(93840) <= 5172716;
srom_1(93841) <= 5710498;
srom_1(93842) <= 6260839;
srom_1(93843) <= 6821157;
srom_1(93844) <= 7388826;
srom_1(93845) <= 7961182;
srom_1(93846) <= 8535544;
srom_1(93847) <= 9109216;
srom_1(93848) <= 9679509;
srom_1(93849) <= 10243748;
srom_1(93850) <= 10799288;
srom_1(93851) <= 11343524;
srom_1(93852) <= 11873903;
srom_1(93853) <= 12387938;
srom_1(93854) <= 12883219;
srom_1(93855) <= 13357423;
srom_1(93856) <= 13808327;
srom_1(93857) <= 14233816;
srom_1(93858) <= 14631894;
srom_1(93859) <= 15000696;
srom_1(93860) <= 15338491;
srom_1(93861) <= 15643696;
srom_1(93862) <= 15914879;
srom_1(93863) <= 16150770;
srom_1(93864) <= 16350260;
srom_1(93865) <= 16512416;
srom_1(93866) <= 16636476;
srom_1(93867) <= 16721859;
srom_1(93868) <= 16768165;
srom_1(93869) <= 16775176;
srom_1(93870) <= 16742860;
srom_1(93871) <= 16671367;
srom_1(93872) <= 16561034;
srom_1(93873) <= 16412378;
srom_1(93874) <= 16226095;
srom_1(93875) <= 16003060;
srom_1(93876) <= 15744318;
srom_1(93877) <= 15451082;
srom_1(93878) <= 15124728;
srom_1(93879) <= 14766786;
srom_1(93880) <= 14378935;
srom_1(93881) <= 13962993;
srom_1(93882) <= 13520911;
srom_1(93883) <= 13054761;
srom_1(93884) <= 12566730;
srom_1(93885) <= 12059107;
srom_1(93886) <= 11534272;
srom_1(93887) <= 10994685;
srom_1(93888) <= 10442877;
srom_1(93889) <= 9881437;
srom_1(93890) <= 9312996;
srom_1(93891) <= 8740220;
srom_1(93892) <= 8165795;
srom_1(93893) <= 7592416;
srom_1(93894) <= 7022769;
srom_1(93895) <= 6459528;
srom_1(93896) <= 5905333;
srom_1(93897) <= 5362783;
srom_1(93898) <= 4834421;
srom_1(93899) <= 4322727;
srom_1(93900) <= 3830099;
srom_1(93901) <= 3358847;
srom_1(93902) <= 2911182;
srom_1(93903) <= 2489202;
srom_1(93904) <= 2094887;
srom_1(93905) <= 1730085;
srom_1(93906) <= 1396507;
srom_1(93907) <= 1095717;
srom_1(93908) <= 829126;
srom_1(93909) <= 597984;
srom_1(93910) <= 403376;
srom_1(93911) <= 246212;
srom_1(93912) <= 127231;
srom_1(93913) <= 46991;
srom_1(93914) <= 5867;
srom_1(93915) <= 4053;
srom_1(93916) <= 41557;
srom_1(93917) <= 118203;
srom_1(93918) <= 233631;
srom_1(93919) <= 387302;
srom_1(93920) <= 578493;
srom_1(93921) <= 806308;
srom_1(93922) <= 1069680;
srom_1(93923) <= 1367372;
srom_1(93924) <= 1697989;
srom_1(93925) <= 2059981;
srom_1(93926) <= 2451650;
srom_1(93927) <= 2871160;
srom_1(93928) <= 3316543;
srom_1(93929) <= 3785710;
srom_1(93930) <= 4276462;
srom_1(93931) <= 4786497;
srom_1(93932) <= 5313424;
srom_1(93933) <= 5854771;
srom_1(93934) <= 6408000;
srom_1(93935) <= 6970518;
srom_1(93936) <= 7539685;
srom_1(93937) <= 8112832;
srom_1(93938) <= 8687273;
srom_1(93939) <= 9260314;
srom_1(93940) <= 9829267;
srom_1(93941) <= 10391464;
srom_1(93942) <= 10944269;
srom_1(93943) <= 11485089;
srom_1(93944) <= 12011389;
srom_1(93945) <= 12520701;
srom_1(93946) <= 13010636;
srom_1(93947) <= 13478896;
srom_1(93948) <= 13923287;
srom_1(93949) <= 14341723;
srom_1(93950) <= 14732243;
srom_1(93951) <= 15093016;
srom_1(93952) <= 15422349;
srom_1(93953) <= 15718699;
srom_1(93954) <= 15980675;
srom_1(93955) <= 16207050;
srom_1(93956) <= 16396761;
srom_1(93957) <= 16548920;
srom_1(93958) <= 16662811;
srom_1(93959) <= 16737903;
srom_1(93960) <= 16773841;
srom_1(93961) <= 16770458;
srom_1(93962) <= 16727770;
srom_1(93963) <= 16645977;
srom_1(93964) <= 16525462;
srom_1(93965) <= 16366790;
srom_1(93966) <= 16170706;
srom_1(93967) <= 15938129;
srom_1(93968) <= 15670150;
srom_1(93969) <= 15368025;
srom_1(93970) <= 15033171;
srom_1(93971) <= 14667159;
srom_1(93972) <= 14271704;
srom_1(93973) <= 13848662;
srom_1(93974) <= 13400015;
srom_1(93975) <= 12927868;
srom_1(93976) <= 12434435;
srom_1(93977) <= 11922030;
srom_1(93978) <= 11393055;
srom_1(93979) <= 10849991;
srom_1(93980) <= 10295385;
srom_1(93981) <= 9731838;
srom_1(93982) <= 9161992;
srom_1(93983) <= 8588519;
srom_1(93984) <= 8014108;
srom_1(93985) <= 7441454;
srom_1(93986) <= 6873241;
srom_1(93987) <= 6312134;
srom_1(93988) <= 5760765;
srom_1(93989) <= 5221718;
srom_1(93990) <= 4697523;
srom_1(93991) <= 4190635;
srom_1(93992) <= 3703434;
srom_1(93993) <= 3238203;
srom_1(93994) <= 2797124;
srom_1(93995) <= 2382265;
srom_1(93996) <= 1995572;
srom_1(93997) <= 1638859;
srom_1(93998) <= 1313797;
srom_1(93999) <= 1021911;
srom_1(94000) <= 764570;
srom_1(94001) <= 542981;
srom_1(94002) <= 358183;
srom_1(94003) <= 211043;
srom_1(94004) <= 102249;
srom_1(94005) <= 32314;
srom_1(94006) <= 1563;
srom_1(94007) <= 10143;
srom_1(94008) <= 58012;
srom_1(94009) <= 144946;
srom_1(94010) <= 270537;
srom_1(94011) <= 434197;
srom_1(94012) <= 635158;
srom_1(94013) <= 872477;
srom_1(94014) <= 1145042;
srom_1(94015) <= 1451575;
srom_1(94016) <= 1790638;
srom_1(94017) <= 2160641;
srom_1(94018) <= 2559849;
srom_1(94019) <= 2986390;
srom_1(94020) <= 3438264;
srom_1(94021) <= 3913351;
srom_1(94022) <= 4409425;
srom_1(94023) <= 4924159;
srom_1(94024) <= 5455138;
srom_1(94025) <= 5999874;
srom_1(94026) <= 6555811;
srom_1(94027) <= 7120342;
srom_1(94028) <= 7690821;
srom_1(94029) <= 8264573;
srom_1(94030) <= 8838905;
srom_1(94031) <= 9411127;
srom_1(94032) <= 9978553;
srom_1(94033) <= 10538523;
srom_1(94034) <= 11088412;
srom_1(94035) <= 11625641;
srom_1(94036) <= 12147690;
srom_1(94037) <= 12652111;
srom_1(94038) <= 13136539;
srom_1(94039) <= 13598703;
srom_1(94040) <= 14036434;
srom_1(94041) <= 14447681;
srom_1(94042) <= 14830515;
srom_1(94043) <= 15183141;
srom_1(94044) <= 15503904;
srom_1(94045) <= 15791302;
srom_1(94046) <= 16043986;
srom_1(94047) <= 16260771;
srom_1(94048) <= 16440641;
srom_1(94049) <= 16582752;
srom_1(94050) <= 16686438;
srom_1(94051) <= 16751212;
srom_1(94052) <= 16776772;
srom_1(94053) <= 16762996;
srom_1(94054) <= 16709950;
srom_1(94055) <= 16617883;
srom_1(94056) <= 16487225;
srom_1(94057) <= 16318590;
srom_1(94058) <= 16112769;
srom_1(94059) <= 15870727;
srom_1(94060) <= 15593598;
srom_1(94061) <= 15282683;
srom_1(94062) <= 14939439;
srom_1(94063) <= 14565476;
srom_1(94064) <= 14162547;
srom_1(94065) <= 13732543;
srom_1(94066) <= 13277479;
srom_1(94067) <= 12799489;
srom_1(94068) <= 12300815;
srom_1(94069) <= 11783796;
srom_1(94070) <= 11250855;
srom_1(94071) <= 10704492;
srom_1(94072) <= 10147269;
srom_1(94073) <= 9581799;
srom_1(94074) <= 9010734;
srom_1(94075) <= 8436752;
srom_1(94076) <= 7862544;
srom_1(94077) <= 7290802;
srom_1(94078) <= 6724209;
srom_1(94079) <= 6165421;
srom_1(94080) <= 5617058;
srom_1(94081) <= 5081691;
srom_1(94082) <= 4561832;
srom_1(94083) <= 4059918;
srom_1(94084) <= 3578303;
srom_1(94085) <= 3119245;
srom_1(94086) <= 2684896;
srom_1(94087) <= 2277295;
srom_1(94088) <= 1898351;
srom_1(94089) <= 1549842;
srom_1(94090) <= 1233403;
srom_1(94091) <= 950517;
srom_1(94092) <= 702511;
srom_1(94093) <= 490547;
srom_1(94094) <= 315620;
srom_1(94095) <= 178550;
srom_1(94096) <= 79980;
srom_1(94097) <= 20372;
srom_1(94098) <= 6;
srom_1(94099) <= 18976;
srom_1(94100) <= 77195;
srom_1(94101) <= 174388;
srom_1(94102) <= 310101;
srom_1(94103) <= 483697;
srom_1(94104) <= 694362;
srom_1(94105) <= 941107;
srom_1(94106) <= 1222777;
srom_1(94107) <= 1538049;
srom_1(94108) <= 1885446;
srom_1(94109) <= 2263339;
srom_1(94110) <= 2669955;
srom_1(94111) <= 3103388;
srom_1(94112) <= 3561605;
srom_1(94113) <= 4042458;
srom_1(94114) <= 4543691;
srom_1(94115) <= 5062954;
srom_1(94116) <= 5597813;
srom_1(94117) <= 6145758;
srom_1(94118) <= 6704221;
srom_1(94119) <= 7270582;
srom_1(94120) <= 7842187;
srom_1(94121) <= 8416353;
srom_1(94122) <= 8990390;
srom_1(94123) <= 9561605;
srom_1(94124) <= 10127319;
srom_1(94125) <= 10684879;
srom_1(94126) <= 11231672;
srom_1(94127) <= 11765132;
srom_1(94128) <= 12282759;
srom_1(94129) <= 12782125;
srom_1(94130) <= 13260888;
srom_1(94131) <= 13716803;
srom_1(94132) <= 14147733;
srom_1(94133) <= 14551656;
srom_1(94134) <= 14926678;
srom_1(94135) <= 15271041;
srom_1(94136) <= 15583130;
srom_1(94137) <= 15861481;
srom_1(94138) <= 16104790;
srom_1(94139) <= 16311914;
srom_1(94140) <= 16481884;
srom_1(94141) <= 16613901;
srom_1(94142) <= 16707348;
srom_1(94143) <= 16761784;
srom_1(94144) <= 16776956;
srom_1(94145) <= 16752792;
srom_1(94146) <= 16689406;
srom_1(94147) <= 16587094;
srom_1(94148) <= 16446337;
srom_1(94149) <= 16267794;
srom_1(94150) <= 16052304;
srom_1(94151) <= 15800875;
srom_1(94152) <= 15514688;
srom_1(94153) <= 15195084;
srom_1(94154) <= 14843562;
srom_1(94155) <= 14461771;
srom_1(94156) <= 14051500;
srom_1(94157) <= 13614674;
srom_1(94158) <= 13153342;
srom_1(94159) <= 12669666;
srom_1(94160) <= 12165914;
srom_1(94161) <= 11644450;
srom_1(94162) <= 11107718;
srom_1(94163) <= 10558234;
srom_1(94164) <= 9998577;
srom_1(94165) <= 9431370;
srom_1(94166) <= 8859273;
srom_1(94167) <= 8284969;
srom_1(94168) <= 7711151;
srom_1(94169) <= 7140510;
srom_1(94170) <= 6575722;
srom_1(94171) <= 6019435;
srom_1(94172) <= 5474257;
srom_1(94173) <= 4942747;
srom_1(94174) <= 4427394;
srom_1(94175) <= 3930618;
srom_1(94176) <= 3454746;
srom_1(94177) <= 3002011;
srom_1(94178) <= 2574536;
srom_1(94179) <= 2174325;
srom_1(94180) <= 1803254;
srom_1(94181) <= 1463065;
srom_1(94182) <= 1155352;
srom_1(94183) <= 881558;
srom_1(94184) <= 642967;
srom_1(94185) <= 440698;
srom_1(94186) <= 275700;
srom_1(94187) <= 148746;
srom_1(94188) <= 60431;
srom_1(94189) <= 11171;
srom_1(94190) <= 1194;
srom_1(94191) <= 30550;
srom_1(94192) <= 99099;
srom_1(94193) <= 206520;
srom_1(94194) <= 352310;
srom_1(94195) <= 535785;
srom_1(94196) <= 756084;
srom_1(94197) <= 1012175;
srom_1(94198) <= 1302857;
srom_1(94199) <= 1626766;
srom_1(94200) <= 1982384;
srom_1(94201) <= 2368043;
srom_1(94202) <= 2781934;
srom_1(94203) <= 3222117;
srom_1(94204) <= 3686527;
srom_1(94205) <= 4172987;
srom_1(94206) <= 4679216;
srom_1(94207) <= 5202839;
srom_1(94208) <= 5741401;
srom_1(94209) <= 6292377;
srom_1(94210) <= 6853183;
srom_1(94211) <= 7421189;
srom_1(94212) <= 7993731;
srom_1(94213) <= 8568125;
srom_1(94214) <= 9141678;
srom_1(94215) <= 9711699;
srom_1(94216) <= 10275515;
srom_1(94217) <= 10830483;
srom_1(94218) <= 11374001;
srom_1(94219) <= 11903519;
srom_1(94220) <= 12416554;
srom_1(94221) <= 12910701;
srom_1(94222) <= 13383642;
srom_1(94223) <= 13833159;
srom_1(94224) <= 14257146;
srom_1(94225) <= 14653612;
srom_1(94226) <= 15020700;
srom_1(94227) <= 15356688;
srom_1(94228) <= 15660000;
srom_1(94229) <= 15929214;
srom_1(94230) <= 16163068;
srom_1(94231) <= 16360464;
srom_1(94232) <= 16520478;
srom_1(94233) <= 16642358;
srom_1(94234) <= 16725534;
srom_1(94235) <= 16769615;
srom_1(94236) <= 16774395;
srom_1(94237) <= 16739850;
srom_1(94238) <= 16666144;
srom_1(94239) <= 16553622;
srom_1(94240) <= 16402811;
srom_1(94241) <= 16214419;
srom_1(94242) <= 15989329;
srom_1(94243) <= 15728596;
srom_1(94244) <= 15433444;
srom_1(94245) <= 15105256;
srom_1(94246) <= 14745572;
srom_1(94247) <= 14356077;
srom_1(94248) <= 13938599;
srom_1(94249) <= 13495095;
srom_1(94250) <= 13027645;
srom_1(94251) <= 12538441;
srom_1(94252) <= 12029777;
srom_1(94253) <= 11504038;
srom_1(94254) <= 10963690;
srom_1(94255) <= 10411266;
srom_1(94256) <= 9849358;
srom_1(94257) <= 9280600;
srom_1(94258) <= 8707658;
srom_1(94259) <= 8133221;
srom_1(94260) <= 7559981;
srom_1(94261) <= 6990627;
srom_1(94262) <= 6427828;
srom_1(94263) <= 5874224;
srom_1(94264) <= 5332412;
srom_1(94265) <= 4804930;
srom_1(94266) <= 4294254;
srom_1(94267) <= 3802777;
srom_1(94268) <= 3332805;
srom_1(94269) <= 2886542;
srom_1(94270) <= 2466079;
srom_1(94271) <= 2073389;
srom_1(94272) <= 1710314;
srom_1(94273) <= 1378555;
srom_1(94274) <= 1079669;
srom_1(94275) <= 815057;
srom_1(94276) <= 585960;
srom_1(94277) <= 393452;
srom_1(94278) <= 238436;
srom_1(94279) <= 121639;
srom_1(94280) <= 43609;
srom_1(94281) <= 4712;
srom_1(94282) <= 5129;
srom_1(94283) <= 44859;
srom_1(94284) <= 123716;
srom_1(94285) <= 241330;
srom_1(94286) <= 397150;
srom_1(94287) <= 590444;
srom_1(94288) <= 820306;
srom_1(94289) <= 1085659;
srom_1(94290) <= 1385257;
srom_1(94291) <= 1717697;
srom_1(94292) <= 2081419;
srom_1(94293) <= 2474718;
srom_1(94294) <= 2895748;
srom_1(94295) <= 3342537;
srom_1(94296) <= 3812989;
srom_1(94297) <= 4304897;
srom_1(94298) <= 4815955;
srom_1(94299) <= 5343766;
srom_1(94300) <= 5885856;
srom_1(94301) <= 6439682;
srom_1(94302) <= 7002647;
srom_1(94303) <= 7572111;
srom_1(94304) <= 8145405;
srom_1(94305) <= 8719838;
srom_1(94306) <= 9292719;
srom_1(94307) <= 9861359;
srom_1(94308) <= 10423094;
srom_1(94309) <= 10975288;
srom_1(94310) <= 11515352;
srom_1(94311) <= 12040754;
srom_1(94312) <= 12549030;
srom_1(94313) <= 13037796;
srom_1(94314) <= 13504760;
srom_1(94315) <= 13947733;
srom_1(94316) <= 14364637;
srom_1(94317) <= 14753518;
srom_1(94318) <= 15112551;
srom_1(94319) <= 15440054;
srom_1(94320) <= 15734490;
srom_1(94321) <= 15994478;
srom_1(94322) <= 16218800;
srom_1(94323) <= 16406404;
srom_1(94324) <= 16556409;
srom_1(94325) <= 16668112;
srom_1(94326) <= 16740991;
srom_1(94327) <= 16774702;
srom_1(94328) <= 16769087;
srom_1(94329) <= 16724174;
srom_1(94330) <= 16640173;
srom_1(94331) <= 16517476;
srom_1(94332) <= 16356661;
srom_1(94333) <= 16158481;
srom_1(94334) <= 15923866;
srom_1(94335) <= 15653915;
srom_1(94336) <= 15349894;
srom_1(94337) <= 15013230;
srom_1(94338) <= 14645500;
srom_1(94339) <= 14248430;
srom_1(94340) <= 13823881;
srom_1(94341) <= 13373844;
srom_1(94342) <= 12900429;
srom_1(94343) <= 12405857;
srom_1(94344) <= 11892447;
srom_1(94345) <= 11362606;
srom_1(94346) <= 10818819;
srom_1(94347) <= 10263636;
srom_1(94348) <= 9699661;
srom_1(94349) <= 9129537;
srom_1(94350) <= 8555939;
srom_1(94351) <= 7981556;
srom_1(94352) <= 7409082;
srom_1(94353) <= 6841201;
srom_1(94354) <= 6280577;
srom_1(94355) <= 5729837;
srom_1(94356) <= 5191566;
srom_1(94357) <= 4668287;
srom_1(94358) <= 4162453;
srom_1(94359) <= 3676438;
srom_1(94360) <= 3212519;
srom_1(94361) <= 2772873;
srom_1(94362) <= 2359561;
srom_1(94363) <= 1974522;
srom_1(94364) <= 1619560;
srom_1(94365) <= 1296340;
srom_1(94366) <= 1006379;
srom_1(94367) <= 751035;
srom_1(94368) <= 531507;
srom_1(94369) <= 348823;
srom_1(94370) <= 203841;
srom_1(94371) <= 97239;
srom_1(94372) <= 29519;
srom_1(94373) <= 997;
srom_1(94374) <= 11808;
srom_1(94375) <= 61901;
srom_1(94376) <= 151040;
srom_1(94377) <= 278808;
srom_1(94378) <= 444606;
srom_1(94379) <= 647656;
srom_1(94380) <= 887005;
srom_1(94381) <= 1161533;
srom_1(94382) <= 1469950;
srom_1(94383) <= 1810812;
srom_1(94384) <= 2182519;
srom_1(94385) <= 2583329;
srom_1(94386) <= 3011361;
srom_1(94387) <= 3464609;
srom_1(94388) <= 3940948;
srom_1(94389) <= 4438143;
srom_1(94390) <= 4953863;
srom_1(94391) <= 5485690;
srom_1(94392) <= 6031130;
srom_1(94393) <= 6587625;
srom_1(94394) <= 7152565;
srom_1(94395) <= 7723301;
srom_1(94396) <= 8297158;
srom_1(94397) <= 8871443;
srom_1(94398) <= 9443464;
srom_1(94399) <= 10010538;
srom_1(94400) <= 10570006;
srom_1(94401) <= 11119246;
srom_1(94402) <= 11655680;
srom_1(94403) <= 12176794;
srom_1(94404) <= 12680143;
srom_1(94405) <= 13163369;
srom_1(94406) <= 13624203;
srom_1(94407) <= 14060487;
srom_1(94408) <= 14470173;
srom_1(94409) <= 14851340;
srom_1(94410) <= 15202201;
srom_1(94411) <= 15521111;
srom_1(94412) <= 15806574;
srom_1(94413) <= 16057252;
srom_1(94414) <= 16271969;
srom_1(94415) <= 16449718;
srom_1(94416) <= 16589666;
srom_1(94417) <= 16691156;
srom_1(94418) <= 16753713;
srom_1(94419) <= 16777043;
srom_1(94420) <= 16761036;
srom_1(94421) <= 16705769;
srom_1(94422) <= 16611499;
srom_1(94423) <= 16478670;
srom_1(94424) <= 16307903;
srom_1(94425) <= 16100000;
srom_1(94426) <= 15855936;
srom_1(94427) <= 15576854;
srom_1(94428) <= 15264065;
srom_1(94429) <= 14919034;
srom_1(94430) <= 14543380;
srom_1(94431) <= 14138864;
srom_1(94432) <= 13707383;
srom_1(94433) <= 13250960;
srom_1(94434) <= 12771737;
srom_1(94435) <= 12271959;
srom_1(94436) <= 11753971;
srom_1(94437) <= 11220201;
srom_1(94438) <= 10673153;
srom_1(94439) <= 10115392;
srom_1(94440) <= 9549534;
srom_1(94441) <= 8978232;
srom_1(94442) <= 8404164;
srom_1(94443) <= 7830024;
srom_1(94444) <= 7258503;
srom_1(94445) <= 6692282;
srom_1(94446) <= 6134015;
srom_1(94447) <= 5586321;
srom_1(94448) <= 5051767;
srom_1(94449) <= 4532862;
srom_1(94450) <= 4032037;
srom_1(94451) <= 3551641;
srom_1(94452) <= 3093928;
srom_1(94453) <= 2661044;
srom_1(94454) <= 2255017;
srom_1(94455) <= 1877754;
srom_1(94456) <= 1531022;
srom_1(94457) <= 1216447;
srom_1(94458) <= 935506;
srom_1(94459) <= 689514;
srom_1(94460) <= 479626;
srom_1(94461) <= 306826;
srom_1(94462) <= 171925;
srom_1(94463) <= 75554;
srom_1(94464) <= 18166;
srom_1(94465) <= 29;
srom_1(94466) <= 21230;
srom_1(94467) <= 81668;
srom_1(94468) <= 181061;
srom_1(94469) <= 318941;
srom_1(94470) <= 494663;
srom_1(94471) <= 707402;
srom_1(94472) <= 956161;
srom_1(94473) <= 1239773;
srom_1(94474) <= 1556908;
srom_1(94475) <= 1906080;
srom_1(94476) <= 2285651;
srom_1(94477) <= 2693840;
srom_1(94478) <= 3128734;
srom_1(94479) <= 3588294;
srom_1(94480) <= 4070364;
srom_1(94481) <= 4572683;
srom_1(94482) <= 5092897;
srom_1(94483) <= 5628565;
srom_1(94484) <= 6177176;
srom_1(94485) <= 6736158;
srom_1(94486) <= 7302888;
srom_1(94487) <= 7874709;
srom_1(94488) <= 8448941;
srom_1(94489) <= 9022889;
srom_1(94490) <= 9593863;
srom_1(94491) <= 10159186;
srom_1(94492) <= 10716205;
srom_1(94493) <= 11262309;
srom_1(94494) <= 11794938;
srom_1(94495) <= 12311593;
srom_1(94496) <= 12809852;
srom_1(94497) <= 13287379;
srom_1(94498) <= 13741933;
srom_1(94499) <= 14171383;
srom_1(94500) <= 14573717;
srom_1(94501) <= 14947046;
srom_1(94502) <= 15289620;
srom_1(94503) <= 15599833;
srom_1(94504) <= 15876230;
srom_1(94505) <= 16117515;
srom_1(94506) <= 16322557;
srom_1(94507) <= 16490394;
srom_1(94508) <= 16620238;
srom_1(94509) <= 16711482;
srom_1(94510) <= 16763697;
srom_1(94511) <= 16776638;
srom_1(94512) <= 16750245;
srom_1(94513) <= 16684641;
srom_1(94514) <= 16580134;
srom_1(94515) <= 16437214;
srom_1(94516) <= 16256552;
srom_1(94517) <= 16038994;
srom_1(94518) <= 15785561;
srom_1(94519) <= 15497441;
srom_1(94520) <= 15175985;
srom_1(94521) <= 14822701;
srom_1(94522) <= 14439245;
srom_1(94523) <= 14027416;
srom_1(94524) <= 13589144;
srom_1(94525) <= 13126485;
srom_1(94526) <= 12641609;
srom_1(94527) <= 12136789;
srom_1(94528) <= 11614392;
srom_1(94529) <= 11076869;
srom_1(94530) <= 10526739;
srom_1(94531) <= 9966583;
srom_1(94532) <= 9399027;
srom_1(94533) <= 8826733;
srom_1(94534) <= 8252385;
srom_1(94535) <= 7678675;
srom_1(94536) <= 7108295;
srom_1(94537) <= 6543918;
srom_1(94538) <= 5988192;
srom_1(94539) <= 5443722;
srom_1(94540) <= 4913061;
srom_1(94541) <= 4398699;
srom_1(94542) <= 3903046;
srom_1(94543) <= 3428428;
srom_1(94544) <= 2977070;
srom_1(94545) <= 2551089;
srom_1(94546) <= 2152482;
srom_1(94547) <= 1783118;
srom_1(94548) <= 1444729;
srom_1(94549) <= 1138903;
srom_1(94550) <= 867073;
srom_1(94551) <= 630514;
srom_1(94552) <= 430335;
srom_1(94553) <= 267475;
srom_1(94554) <= 142699;
srom_1(94555) <= 56590;
srom_1(94556) <= 9553;
srom_1(94557) <= 1808;
srom_1(94558) <= 33391;
srom_1(94559) <= 104155;
srom_1(94560) <= 213768;
srom_1(94561) <= 361716;
srom_1(94562) <= 547304;
srom_1(94563) <= 769663;
srom_1(94564) <= 1027749;
srom_1(94565) <= 1320354;
srom_1(94566) <= 1646103;
srom_1(94567) <= 2003471;
srom_1(94568) <= 2390781;
srom_1(94569) <= 2806216;
srom_1(94570) <= 3247829;
srom_1(94571) <= 3713550;
srom_1(94572) <= 4201193;
srom_1(94573) <= 4708472;
srom_1(94574) <= 5233009;
srom_1(94575) <= 5772343;
srom_1(94576) <= 6323946;
srom_1(94577) <= 6885231;
srom_1(94578) <= 7453566;
srom_1(94579) <= 8026286;
srom_1(94580) <= 8600704;
srom_1(94581) <= 9174128;
srom_1(94582) <= 9743868;
srom_1(94583) <= 10307254;
srom_1(94584) <= 10861641;
srom_1(94585) <= 11404432;
srom_1(94586) <= 11933081;
srom_1(94587) <= 12445109;
srom_1(94588) <= 12938114;
srom_1(94589) <= 13409785;
srom_1(94590) <= 13857909;
srom_1(94591) <= 14280387;
srom_1(94592) <= 14675236;
srom_1(94593) <= 15040605;
srom_1(94594) <= 15374780;
srom_1(94595) <= 15676194;
srom_1(94596) <= 15943435;
srom_1(94597) <= 16175248;
srom_1(94598) <= 16370548;
srom_1(94599) <= 16528417;
srom_1(94600) <= 16648116;
srom_1(94601) <= 16729083;
srom_1(94602) <= 16770938;
srom_1(94603) <= 16773486;
srom_1(94604) <= 16736715;
srom_1(94605) <= 16660796;
srom_1(94606) <= 16546087;
srom_1(94607) <= 16393124;
srom_1(94608) <= 16202625;
srom_1(94609) <= 15975483;
srom_1(94610) <= 15712764;
srom_1(94611) <= 15415700;
srom_1(94612) <= 15085683;
srom_1(94613) <= 14724261;
srom_1(94614) <= 14333129;
srom_1(94615) <= 13914121;
srom_1(94616) <= 13469202;
srom_1(94617) <= 13000459;
srom_1(94618) <= 12510089;
srom_1(94619) <= 12000392;
srom_1(94620) <= 11473758;
srom_1(94621) <= 10932656;
srom_1(94622) <= 10379625;
srom_1(94623) <= 9817257;
srom_1(94624) <= 9248190;
srom_1(94625) <= 8675092;
srom_1(94626) <= 8100650;
srom_1(94627) <= 7527559;
srom_1(94628) <= 6958505;
srom_1(94629) <= 6396158;
srom_1(94630) <= 5843154;
srom_1(94631) <= 5302087;
srom_1(94632) <= 4775493;
srom_1(94633) <= 4265842;
srom_1(94634) <= 3775525;
srom_1(94635) <= 3306839;
srom_1(94636) <= 2861984;
srom_1(94637) <= 2443045;
srom_1(94638) <= 2051987;
srom_1(94639) <= 1690644;
srom_1(94640) <= 1360709;
srom_1(94641) <= 1063731;
srom_1(94642) <= 801102;
srom_1(94643) <= 574053;
srom_1(94644) <= 383649;
srom_1(94645) <= 230783;
srom_1(94646) <= 116172;
srom_1(94647) <= 40354;
srom_1(94648) <= 3683;
srom_1(94649) <= 6332;
srom_1(94650) <= 48288;
srom_1(94651) <= 129355;
srom_1(94652) <= 249152;
srom_1(94653) <= 407118;
srom_1(94654) <= 602512;
srom_1(94655) <= 834418;
srom_1(94656) <= 1101748;
srom_1(94657) <= 1403248;
srom_1(94658) <= 1737505;
srom_1(94659) <= 2102952;
srom_1(94660) <= 2497874;
srom_1(94661) <= 2920420;
srom_1(94662) <= 3368608;
srom_1(94663) <= 3840336;
srom_1(94664) <= 4333393;
srom_1(94665) <= 4845466;
srom_1(94666) <= 5374154;
srom_1(94667) <= 5916978;
srom_1(94668) <= 6471393;
srom_1(94669) <= 7034797;
srom_1(94670) <= 7604551;
srom_1(94671) <= 8177980;
srom_1(94672) <= 8752398;
srom_1(94673) <= 9325110;
srom_1(94674) <= 9893430;
srom_1(94675) <= 10454693;
srom_1(94676) <= 11006268;
srom_1(94677) <= 11545568;
srom_1(94678) <= 12070064;
srom_1(94679) <= 12577296;
srom_1(94680) <= 13064886;
srom_1(94681) <= 13530547;
srom_1(94682) <= 13972096;
srom_1(94683) <= 14387462;
srom_1(94684) <= 14774697;
srom_1(94685) <= 15131985;
srom_1(94686) <= 15457652;
srom_1(94687) <= 15750170;
srom_1(94688) <= 16008166;
srom_1(94689) <= 16230432;
srom_1(94690) <= 16415925;
srom_1(94691) <= 16563775;
srom_1(94692) <= 16673289;
srom_1(94693) <= 16743953;
srom_1(94694) <= 16775436;
srom_1(94695) <= 16767590;
srom_1(94696) <= 16720452;
srom_1(94697) <= 16634244;
srom_1(94698) <= 16509369;
srom_1(94699) <= 16346413;
srom_1(94700) <= 16146139;
srom_1(94701) <= 15909489;
srom_1(94702) <= 15637570;
srom_1(94703) <= 15331658;
srom_1(94704) <= 14993188;
srom_1(94705) <= 14623747;
srom_1(94706) <= 14225067;
srom_1(94707) <= 13799018;
srom_1(94708) <= 13347597;
srom_1(94709) <= 12872923;
srom_1(94710) <= 12377219;
srom_1(94711) <= 11862812;
srom_1(94712) <= 11332113;
srom_1(94713) <= 10787611;
srom_1(94714) <= 10231859;
srom_1(94715) <= 9667463;
srom_1(94716) <= 9097071;
srom_1(94717) <= 8523356;
srom_1(94718) <= 7949010;
srom_1(94719) <= 7376724;
srom_1(94720) <= 6809184;
srom_1(94721) <= 6249050;
srom_1(94722) <= 5698950;
srom_1(94723) <= 5161462;
srom_1(94724) <= 4639107;
srom_1(94725) <= 4134335;
srom_1(94726) <= 3649513;
srom_1(94727) <= 3186914;
srom_1(94728) <= 2748708;
srom_1(94729) <= 2336949;
srom_1(94730) <= 1953568;
srom_1(94731) <= 1600363;
srom_1(94732) <= 1278991;
srom_1(94733) <= 990958;
srom_1(94734) <= 737615;
srom_1(94735) <= 520151;
srom_1(94736) <= 339584;
srom_1(94737) <= 196762;
srom_1(94738) <= 92354;
srom_1(94739) <= 26851;
srom_1(94740) <= 558;
srom_1(94741) <= 13600;
srom_1(94742) <= 65915;
srom_1(94743) <= 157258;
srom_1(94744) <= 287201;
srom_1(94745) <= 455134;
srom_1(94746) <= 660270;
srom_1(94747) <= 901646;
srom_1(94748) <= 1178132;
srom_1(94749) <= 1488430;
srom_1(94750) <= 1831085;
srom_1(94751) <= 2204491;
srom_1(94752) <= 2606896;
srom_1(94753) <= 3036414;
srom_1(94754) <= 3491030;
srom_1(94755) <= 3968612;
srom_1(94756) <= 4466921;
srom_1(94757) <= 4983620;
srom_1(94758) <= 5516287;
srom_1(94759) <= 6062422;
srom_1(94760) <= 6619466;
srom_1(94761) <= 7184806;
srom_1(94762) <= 7755792;
srom_1(94763) <= 8329744;
srom_1(94764) <= 8903973;
srom_1(94765) <= 9475785;
srom_1(94766) <= 10042499;
srom_1(94767) <= 10601457;
srom_1(94768) <= 11150038;
srom_1(94769) <= 11685670;
srom_1(94770) <= 12205841;
srom_1(94771) <= 12708111;
srom_1(94772) <= 13190126;
srom_1(94773) <= 13649625;
srom_1(94774) <= 14084454;
srom_1(94775) <= 14492572;
srom_1(94776) <= 14872067;
srom_1(94777) <= 15221159;
srom_1(94778) <= 15538210;
srom_1(94779) <= 15821735;
srom_1(94780) <= 16070403;
srom_1(94781) <= 16283048;
srom_1(94782) <= 16458674;
srom_1(94783) <= 16596457;
srom_1(94784) <= 16695750;
srom_1(94785) <= 16756087;
srom_1(94786) <= 16777187;
srom_1(94787) <= 16758950;
srom_1(94788) <= 16701462;
srom_1(94789) <= 16604992;
srom_1(94790) <= 16469992;
srom_1(94791) <= 16297096;
srom_1(94792) <= 16087114;
srom_1(94793) <= 15841032;
srom_1(94794) <= 15560002;
srom_1(94795) <= 15245343;
srom_1(94796) <= 14898531;
srom_1(94797) <= 14521191;
srom_1(94798) <= 14115094;
srom_1(94799) <= 13682143;
srom_1(94800) <= 13224369;
srom_1(94801) <= 12743918;
srom_1(94802) <= 12243044;
srom_1(94803) <= 11724095;
srom_1(94804) <= 11189505;
srom_1(94805) <= 10641780;
srom_1(94806) <= 10083490;
srom_1(94807) <= 9517251;
srom_1(94808) <= 8945720;
srom_1(94809) <= 8371577;
srom_1(94810) <= 7797513;
srom_1(94811) <= 7226221;
srom_1(94812) <= 6660380;
srom_1(94813) <= 6102643;
srom_1(94814) <= 5555626;
srom_1(94815) <= 5021894;
srom_1(94816) <= 4503949;
srom_1(94817) <= 4004221;
srom_1(94818) <= 3525053;
srom_1(94819) <= 3068692;
srom_1(94820) <= 2637277;
srom_1(94821) <= 2232833;
srom_1(94822) <= 1857255;
srom_1(94823) <= 1512305;
srom_1(94824) <= 1199600;
srom_1(94825) <= 920607;
srom_1(94826) <= 676634;
srom_1(94827) <= 468825;
srom_1(94828) <= 298154;
srom_1(94829) <= 165423;
srom_1(94830) <= 71253;
srom_1(94831) <= 16085;
srom_1(94832) <= 180;
srom_1(94833) <= 23610;
srom_1(94834) <= 86267;
srom_1(94835) <= 187857;
srom_1(94836) <= 327902;
srom_1(94837) <= 505747;
srom_1(94838) <= 720558;
srom_1(94839) <= 971326;
srom_1(94840) <= 1256877;
srom_1(94841) <= 1575871;
srom_1(94842) <= 1926812;
srom_1(94843) <= 2308055;
srom_1(94844) <= 2717811;
srom_1(94845) <= 3154160;
srom_1(94846) <= 3615055;
srom_1(94847) <= 4098334;
srom_1(94848) <= 4601733;
srom_1(94849) <= 5122889;
srom_1(94850) <= 5659359;
srom_1(94851) <= 6208628;
srom_1(94852) <= 6768119;
srom_1(94853) <= 7335210;
srom_1(94854) <= 7907240;
srom_1(94855) <= 8481527;
srom_1(94856) <= 9055379;
srom_1(94857) <= 9626104;
srom_1(94858) <= 10191026;
srom_1(94859) <= 10747496;
srom_1(94860) <= 11292904;
srom_1(94861) <= 11824693;
srom_1(94862) <= 12340368;
srom_1(94863) <= 12837513;
srom_1(94864) <= 13313795;
srom_1(94865) <= 13766982;
srom_1(94866) <= 14194947;
srom_1(94867) <= 14595684;
srom_1(94868) <= 14967315;
srom_1(94869) <= 15308095;
srom_1(94870) <= 15616428;
srom_1(94871) <= 15890866;
srom_1(94872) <= 16130125;
srom_1(94873) <= 16333080;
srom_1(94874) <= 16498781;
srom_1(94875) <= 16626451;
srom_1(94876) <= 16715491;
srom_1(94877) <= 16765483;
srom_1(94878) <= 16776193;
srom_1(94879) <= 16747570;
srom_1(94880) <= 16679750;
srom_1(94881) <= 16573050;
srom_1(94882) <= 16427970;
srom_1(94883) <= 16245190;
srom_1(94884) <= 16025569;
srom_1(94885) <= 15770135;
srom_1(94886) <= 15480086;
srom_1(94887) <= 15156784;
srom_1(94888) <= 14801743;
srom_1(94889) <= 14416628;
srom_1(94890) <= 14003246;
srom_1(94891) <= 13563535;
srom_1(94892) <= 13099557;
srom_1(94893) <= 12613488;
srom_1(94894) <= 12107607;
srom_1(94895) <= 11584286;
srom_1(94896) <= 11045979;
srom_1(94897) <= 10495212;
srom_1(94898) <= 9934565;
srom_1(94899) <= 9366669;
srom_1(94900) <= 8794187;
srom_1(94901) <= 8219803;
srom_1(94902) <= 7646210;
srom_1(94903) <= 7076098;
srom_1(94904) <= 6512142;
srom_1(94905) <= 5956985;
srom_1(94906) <= 5413230;
srom_1(94907) <= 4883428;
srom_1(94908) <= 4370063;
srom_1(94909) <= 3875543;
srom_1(94910) <= 3402185;
srom_1(94911) <= 2952211;
srom_1(94912) <= 2527730;
srom_1(94913) <= 2130733;
srom_1(94914) <= 1763080;
srom_1(94915) <= 1426498;
srom_1(94916) <= 1122563;
srom_1(94917) <= 852701;
srom_1(94918) <= 618177;
srom_1(94919) <= 420091;
srom_1(94920) <= 259373;
srom_1(94921) <= 136776;
srom_1(94922) <= 52874;
srom_1(94923) <= 8061;
srom_1(94924) <= 2547;
srom_1(94925) <= 36359;
srom_1(94926) <= 109337;
srom_1(94927) <= 221140;
srom_1(94928) <= 371242;
srom_1(94929) <= 558941;
srom_1(94930) <= 783356;
srom_1(94931) <= 1043434;
srom_1(94932) <= 1337957;
srom_1(94933) <= 1665542;
srom_1(94934) <= 2024654;
srom_1(94935) <= 2413609;
srom_1(94936) <= 2830583;
srom_1(94937) <= 3273620;
srom_1(94938) <= 3740643;
srom_1(94939) <= 4229462;
srom_1(94940) <= 4737784;
srom_1(94941) <= 5263227;
srom_1(94942) <= 5803325;
srom_1(94943) <= 6355547;
srom_1(94944) <= 6917303;
srom_1(94945) <= 7485958;
srom_1(94946) <= 8058846;
srom_1(94947) <= 8633280;
srom_1(94948) <= 9206567;
srom_1(94949) <= 9776018;
srom_1(94950) <= 10338963;
srom_1(94951) <= 10892762;
srom_1(94952) <= 11434819;
srom_1(94953) <= 11962590;
srom_1(94954) <= 12473602;
srom_1(94955) <= 12965458;
srom_1(94956) <= 13435852;
srom_1(94957) <= 13882577;
srom_1(94958) <= 14303539;
srom_1(94959) <= 14696764;
srom_1(94960) <= 15060408;
srom_1(94961) <= 15392766;
srom_1(94962) <= 15692279;
srom_1(94963) <= 15957542;
srom_1(94964) <= 16187312;
srom_1(94965) <= 16380511;
srom_1(94966) <= 16536233;
srom_1(94967) <= 16653748;
srom_1(94968) <= 16732506;
srom_1(94969) <= 16772135;
srom_1(94970) <= 16772452;
srom_1(94971) <= 16733454;
srom_1(94972) <= 16655324;
srom_1(94973) <= 16538428;
srom_1(94974) <= 16383315;
srom_1(94975) <= 16190713;
srom_1(94976) <= 15961523;
srom_1(94977) <= 15696821;
srom_1(94978) <= 15397849;
srom_1(94979) <= 15066008;
srom_1(94980) <= 14702855;
srom_1(94981) <= 14310091;
srom_1(94982) <= 13889560;
srom_1(94983) <= 13443233;
srom_1(94984) <= 12973203;
srom_1(94985) <= 12481674;
srom_1(94986) <= 11970952;
srom_1(94987) <= 11443431;
srom_1(94988) <= 10901584;
srom_1(94989) <= 10347953;
srom_1(94990) <= 9785135;
srom_1(94991) <= 9215767;
srom_1(94992) <= 8642521;
srom_1(94993) <= 8068084;
srom_1(94994) <= 7495150;
srom_1(94995) <= 6926405;
srom_1(94996) <= 6364518;
srom_1(94997) <= 5812122;
srom_1(94998) <= 5271808;
srom_1(94999) <= 4746110;
srom_1(95000) <= 4237493;
srom_1(95001) <= 3748342;
srom_1(95002) <= 3280950;
srom_1(95003) <= 2837510;
srom_1(95004) <= 2420102;
srom_1(95005) <= 2030681;
srom_1(95006) <= 1671075;
srom_1(95007) <= 1342970;
srom_1(95008) <= 1047904;
srom_1(95009) <= 787261;
srom_1(95010) <= 562264;
srom_1(95011) <= 373967;
srom_1(95012) <= 223254;
srom_1(95013) <= 110830;
srom_1(95014) <= 37224;
srom_1(95015) <= 2780;
srom_1(95016) <= 7661;
srom_1(95017) <= 51842;
srom_1(95018) <= 135118;
srom_1(95019) <= 257097;
srom_1(95020) <= 417207;
srom_1(95021) <= 614698;
srom_1(95022) <= 848644;
srom_1(95023) <= 1117947;
srom_1(95024) <= 1421345;
srom_1(95025) <= 1757414;
srom_1(95026) <= 2124580;
srom_1(95027) <= 2521119;
srom_1(95028) <= 2945174;
srom_1(95029) <= 3394754;
srom_1(95030) <= 3867752;
srom_1(95031) <= 4361951;
srom_1(95032) <= 4875031;
srom_1(95033) <= 5404588;
srom_1(95034) <= 5948138;
srom_1(95035) <= 6503132;
srom_1(95036) <= 7066968;
srom_1(95037) <= 7637002;
srom_1(95038) <= 8210560;
srom_1(95039) <= 8784952;
srom_1(95040) <= 9357487;
srom_1(95041) <= 9925478;
srom_1(95042) <= 10486262;
srom_1(95043) <= 11037209;
srom_1(95044) <= 11575736;
srom_1(95045) <= 12099318;
srom_1(95046) <= 12605498;
srom_1(95047) <= 13091905;
srom_1(95048) <= 13556256;
srom_1(95049) <= 13996374;
srom_1(95050) <= 14410195;
srom_1(95051) <= 14795779;
srom_1(95052) <= 15151318;
srom_1(95053) <= 15475144;
srom_1(95054) <= 15765738;
srom_1(95055) <= 16021739;
srom_1(95056) <= 16241946;
srom_1(95057) <= 16425325;
srom_1(95058) <= 16571018;
srom_1(95059) <= 16678340;
srom_1(95060) <= 16746789;
srom_1(95061) <= 16776043;
srom_1(95062) <= 16765966;
srom_1(95063) <= 16716605;
srom_1(95064) <= 16628191;
srom_1(95065) <= 16501138;
srom_1(95066) <= 16336044;
srom_1(95067) <= 16133680;
srom_1(95068) <= 15894998;
srom_1(95069) <= 15621115;
srom_1(95070) <= 15313317;
srom_1(95071) <= 14973047;
srom_1(95072) <= 14601899;
srom_1(95073) <= 14201616;
srom_1(95074) <= 13774073;
srom_1(95075) <= 13321276;
srom_1(95076) <= 12845348;
srom_1(95077) <= 12348521;
srom_1(95078) <= 11833124;
srom_1(95079) <= 11301575;
srom_1(95080) <= 10756366;
srom_1(95081) <= 10200054;
srom_1(95082) <= 9635247;
srom_1(95083) <= 9064594;
srom_1(95084) <= 8490772;
srom_1(95085) <= 7916470;
srom_1(95086) <= 7344382;
srom_1(95087) <= 6777191;
srom_1(95088) <= 6217557;
srom_1(95089) <= 5668103;
srom_1(95090) <= 5131407;
srom_1(95091) <= 4609984;
srom_1(95092) <= 4106281;
srom_1(95093) <= 3622660;
srom_1(95094) <= 3161387;
srom_1(95095) <= 2724627;
srom_1(95096) <= 2314427;
srom_1(95097) <= 1932711;
srom_1(95098) <= 1581269;
srom_1(95099) <= 1261749;
srom_1(95100) <= 975649;
srom_1(95101) <= 724311;
srom_1(95102) <= 508913;
srom_1(95103) <= 330467;
srom_1(95104) <= 189807;
srom_1(95105) <= 87595;
srom_1(95106) <= 24308;
srom_1(95107) <= 245;
srom_1(95108) <= 15518;
srom_1(95109) <= 70055;
srom_1(95110) <= 163601;
srom_1(95111) <= 295716;
srom_1(95112) <= 465782;
srom_1(95113) <= 673001;
srom_1(95114) <= 916401;
srom_1(95115) <= 1194840;
srom_1(95116) <= 1507014;
srom_1(95117) <= 1851457;
srom_1(95118) <= 2226556;
srom_1(95119) <= 2630551;
srom_1(95120) <= 3061547;
srom_1(95121) <= 3517524;
srom_1(95122) <= 3996342;
srom_1(95123) <= 4495758;
srom_1(95124) <= 5013428;
srom_1(95125) <= 5546926;
srom_1(95126) <= 6093750;
srom_1(95127) <= 6651335;
srom_1(95128) <= 7217066;
srom_1(95129) <= 7788291;
srom_1(95130) <= 8362332;
srom_1(95131) <= 8936495;
srom_1(95132) <= 9508090;
srom_1(95133) <= 10074434;
srom_1(95134) <= 10632873;
srom_1(95135) <= 11180789;
srom_1(95136) <= 11715610;
srom_1(95137) <= 12234830;
srom_1(95138) <= 12736014;
srom_1(95139) <= 13216812;
srom_1(95140) <= 13674968;
srom_1(95141) <= 14108335;
srom_1(95142) <= 14514880;
srom_1(95143) <= 14892696;
srom_1(95144) <= 15240013;
srom_1(95145) <= 15555201;
srom_1(95146) <= 15836783;
srom_1(95147) <= 16083438;
srom_1(95148) <= 16294008;
srom_1(95149) <= 16467508;
srom_1(95150) <= 16603123;
srom_1(95151) <= 16700217;
srom_1(95152) <= 16758336;
srom_1(95153) <= 16777205;
srom_1(95154) <= 16756738;
srom_1(95155) <= 16697030;
srom_1(95156) <= 16598360;
srom_1(95157) <= 16461193;
srom_1(95158) <= 16286170;
srom_1(95159) <= 16074113;
srom_1(95160) <= 15826015;
srom_1(95161) <= 15543041;
srom_1(95162) <= 15226518;
srom_1(95163) <= 14877929;
srom_1(95164) <= 14498910;
srom_1(95165) <= 14091237;
srom_1(95166) <= 13656823;
srom_1(95167) <= 13197704;
srom_1(95168) <= 12716034;
srom_1(95169) <= 12214071;
srom_1(95170) <= 11694169;
srom_1(95171) <= 11158766;
srom_1(95172) <= 10610373;
srom_1(95173) <= 10051561;
srom_1(95174) <= 9484951;
srom_1(95175) <= 8913200;
srom_1(95176) <= 8338989;
srom_1(95177) <= 7765011;
srom_1(95178) <= 7193956;
srom_1(95179) <= 6628504;
srom_1(95180) <= 6071306;
srom_1(95181) <= 5524974;
srom_1(95182) <= 4992071;
srom_1(95183) <= 4475096;
srom_1(95184) <= 3976472;
srom_1(95185) <= 3498538;
srom_1(95186) <= 3043536;
srom_1(95187) <= 2613598;
srom_1(95188) <= 2210741;
srom_1(95189) <= 1836855;
srom_1(95190) <= 1493691;
srom_1(95191) <= 1182861;
srom_1(95192) <= 905821;
srom_1(95193) <= 663870;
srom_1(95194) <= 458143;
srom_1(95195) <= 289604;
srom_1(95196) <= 159045;
srom_1(95197) <= 67077;
srom_1(95198) <= 14131;
srom_1(95199) <= 457;
srom_1(95200) <= 26117;
srom_1(95201) <= 90991;
srom_1(95202) <= 194776;
srom_1(95203) <= 336985;
srom_1(95204) <= 516951;
srom_1(95205) <= 733829;
srom_1(95206) <= 986604;
srom_1(95207) <= 1274088;
srom_1(95208) <= 1594936;
srom_1(95209) <= 1947641;
srom_1(95210) <= 2330550;
srom_1(95211) <= 2741867;
srom_1(95212) <= 3179664;
srom_1(95213) <= 3641888;
srom_1(95214) <= 4126370;
srom_1(95215) <= 4630840;
srom_1(95216) <= 5152931;
srom_1(95217) <= 5690195;
srom_1(95218) <= 6240113;
srom_1(95219) <= 6800106;
srom_1(95220) <= 7367547;
srom_1(95221) <= 7939778;
srom_1(95222) <= 8514112;
srom_1(95223) <= 9087859;
srom_1(95224) <= 9658326;
srom_1(95225) <= 10222839;
srom_1(95226) <= 10778751;
srom_1(95227) <= 11323454;
srom_1(95228) <= 11854395;
srom_1(95229) <= 12369084;
srom_1(95230) <= 12865107;
srom_1(95231) <= 13340138;
srom_1(95232) <= 13791949;
srom_1(95233) <= 14218423;
srom_1(95234) <= 14617558;
srom_1(95235) <= 14987484;
srom_1(95236) <= 15326465;
srom_1(95237) <= 15632913;
srom_1(95238) <= 15905389;
srom_1(95239) <= 16142617;
srom_1(95240) <= 16343483;
srom_1(95241) <= 16507046;
srom_1(95242) <= 16632539;
srom_1(95243) <= 16719374;
srom_1(95244) <= 16767142;
srom_1(95245) <= 16775621;
srom_1(95246) <= 16744770;
srom_1(95247) <= 16674734;
srom_1(95248) <= 16565842;
srom_1(95249) <= 16418604;
srom_1(95250) <= 16233710;
srom_1(95251) <= 16012028;
srom_1(95252) <= 15754598;
srom_1(95253) <= 15462625;
srom_1(95254) <= 15137480;
srom_1(95255) <= 14780688;
srom_1(95256) <= 14393920;
srom_1(95257) <= 13978992;
srom_1(95258) <= 13537848;
srom_1(95259) <= 13072558;
srom_1(95260) <= 12585303;
srom_1(95261) <= 12078368;
srom_1(95262) <= 11554131;
srom_1(95263) <= 11015050;
srom_1(95264) <= 10463652;
srom_1(95265) <= 9902524;
srom_1(95266) <= 9334296;
srom_1(95267) <= 8761634;
srom_1(95268) <= 8187223;
srom_1(95269) <= 7613755;
srom_1(95270) <= 7043922;
srom_1(95271) <= 6480394;
srom_1(95272) <= 5925814;
srom_1(95273) <= 5382784;
srom_1(95274) <= 4853848;
srom_1(95275) <= 4341488;
srom_1(95276) <= 3848107;
srom_1(95277) <= 3376018;
srom_1(95278) <= 2927434;
srom_1(95279) <= 2504460;
srom_1(95280) <= 2109078;
srom_1(95281) <= 1743143;
srom_1(95282) <= 1408371;
srom_1(95283) <= 1106332;
srom_1(95284) <= 838442;
srom_1(95285) <= 605957;
srom_1(95286) <= 409968;
srom_1(95287) <= 251394;
srom_1(95288) <= 130977;
srom_1(95289) <= 49284;
srom_1(95290) <= 6696;
srom_1(95291) <= 3414;
srom_1(95292) <= 39453;
srom_1(95293) <= 114644;
srom_1(95294) <= 228635;
srom_1(95295) <= 380890;
srom_1(95296) <= 570697;
srom_1(95297) <= 797164;
srom_1(95298) <= 1059230;
srom_1(95299) <= 1355666;
srom_1(95300) <= 1685082;
srom_1(95301) <= 2045933;
srom_1(95302) <= 2436527;
srom_1(95303) <= 2855033;
srom_1(95304) <= 3299487;
srom_1(95305) <= 3767806;
srom_1(95306) <= 4257793;
srom_1(95307) <= 4767152;
srom_1(95308) <= 5293492;
srom_1(95309) <= 5834347;
srom_1(95310) <= 6387179;
srom_1(95311) <= 6949397;
srom_1(95312) <= 7518363;
srom_1(95313) <= 8091411;
srom_1(95314) <= 8665852;
srom_1(95315) <= 9238993;
srom_1(95316) <= 9808146;
srom_1(95317) <= 10370643;
srom_1(95318) <= 10923845;
srom_1(95319) <= 11465159;
srom_1(95320) <= 11992045;
srom_1(95321) <= 12502034;
srom_1(95322) <= 12992734;
srom_1(95323) <= 13461843;
srom_1(95324) <= 13907162;
srom_1(95325) <= 14326602;
srom_1(95326) <= 14718198;
srom_1(95327) <= 15080111;
srom_1(95328) <= 15410646;
srom_1(95329) <= 15708253;
srom_1(95330) <= 15971534;
srom_1(95331) <= 16199257;
srom_1(95332) <= 16390353;
srom_1(95333) <= 16543926;
srom_1(95334) <= 16659257;
srom_1(95335) <= 16735803;
srom_1(95336) <= 16773206;
srom_1(95337) <= 16771291;
srom_1(95338) <= 16730067;
srom_1(95339) <= 16649726;
srom_1(95340) <= 16530647;
srom_1(95341) <= 16373386;
srom_1(95342) <= 16178683;
srom_1(95343) <= 15947449;
srom_1(95344) <= 15680769;
srom_1(95345) <= 15379893;
srom_1(95346) <= 15046233;
srom_1(95347) <= 14681353;
srom_1(95348) <= 14286964;
srom_1(95349) <= 13864916;
srom_1(95350) <= 13417187;
srom_1(95351) <= 12945878;
srom_1(95352) <= 12453198;
srom_1(95353) <= 11941458;
srom_1(95354) <= 11413057;
srom_1(95355) <= 10870474;
srom_1(95356) <= 10316252;
srom_1(95357) <= 9752991;
srom_1(95358) <= 9183332;
srom_1(95359) <= 8609946;
srom_1(95360) <= 8035522;
srom_1(95361) <= 7462754;
srom_1(95362) <= 6894328;
srom_1(95363) <= 6332908;
srom_1(95364) <= 5781129;
srom_1(95365) <= 5241577;
srom_1(95366) <= 4716782;
srom_1(95367) <= 4209206;
srom_1(95368) <= 3721229;
srom_1(95369) <= 3255138;
srom_1(95370) <= 2813120;
srom_1(95371) <= 2397248;
srom_1(95372) <= 2009471;
srom_1(95373) <= 1651608;
srom_1(95374) <= 1325337;
srom_1(95375) <= 1032188;
srom_1(95376) <= 773536;
srom_1(95377) <= 550593;
srom_1(95378) <= 364406;
srom_1(95379) <= 215847;
srom_1(95380) <= 105613;
srom_1(95381) <= 34220;
srom_1(95382) <= 2005;
srom_1(95383) <= 9117;
srom_1(95384) <= 55523;
srom_1(95385) <= 141006;
srom_1(95386) <= 265164;
srom_1(95387) <= 427417;
srom_1(95388) <= 627002;
srom_1(95389) <= 862984;
srom_1(95390) <= 1134256;
srom_1(95391) <= 1439546;
srom_1(95392) <= 1777423;
srom_1(95393) <= 2146302;
srom_1(95394) <= 2544453;
srom_1(95395) <= 2970010;
srom_1(95396) <= 3420976;
srom_1(95397) <= 3895237;
srom_1(95398) <= 4390569;
srom_1(95399) <= 4904649;
srom_1(95400) <= 5435067;
srom_1(95401) <= 5979335;
srom_1(95402) <= 6534900;
srom_1(95403) <= 7099159;
srom_1(95404) <= 7669464;
srom_1(95405) <= 8243141;
srom_1(95406) <= 8817501;
srom_1(95407) <= 9389849;
srom_1(95408) <= 9957502;
srom_1(95409) <= 10517798;
srom_1(95410) <= 11068110;
srom_1(95411) <= 11605856;
srom_1(95412) <= 12128516;
srom_1(95413) <= 12633638;
srom_1(95414) <= 13118853;
srom_1(95415) <= 13581887;
srom_1(95416) <= 14020567;
srom_1(95417) <= 14432838;
srom_1(95418) <= 14816765;
srom_1(95419) <= 15170548;
srom_1(95420) <= 15492528;
srom_1(95421) <= 15781196;
srom_1(95422) <= 16035197;
srom_1(95423) <= 16253341;
srom_1(95424) <= 16434604;
srom_1(95425) <= 16578137;
srom_1(95426) <= 16683266;
srom_1(95427) <= 16749499;
srom_1(95428) <= 16776524;
srom_1(95429) <= 16764216;
srom_1(95430) <= 16712632;
srom_1(95431) <= 16622013;
srom_1(95432) <= 16492786;
srom_1(95433) <= 16325555;
srom_1(95434) <= 16121104;
srom_1(95435) <= 15880394;
srom_1(95436) <= 15604552;
srom_1(95437) <= 15294872;
srom_1(95438) <= 14952806;
srom_1(95439) <= 14579958;
srom_1(95440) <= 14178077;
srom_1(95441) <= 13749047;
srom_1(95442) <= 13294880;
srom_1(95443) <= 12817706;
srom_1(95444) <= 12319763;
srom_1(95445) <= 11803384;
srom_1(95446) <= 11270993;
srom_1(95447) <= 10725085;
srom_1(95448) <= 10168221;
srom_1(95449) <= 9603012;
srom_1(95450) <= 9032107;
srom_1(95451) <= 8458186;
srom_1(95452) <= 7883937;
srom_1(95453) <= 7312056;
srom_1(95454) <= 6745222;
srom_1(95455) <= 6186096;
srom_1(95456) <= 5637297;
srom_1(95457) <= 5101400;
srom_1(95458) <= 4580918;
srom_1(95459) <= 4078292;
srom_1(95460) <= 3595878;
srom_1(95461) <= 3135939;
srom_1(95462) <= 2700632;
srom_1(95463) <= 2291997;
srom_1(95464) <= 1911952;
srom_1(95465) <= 1562277;
srom_1(95466) <= 1244614;
srom_1(95467) <= 960452;
srom_1(95468) <= 711122;
srom_1(95469) <= 497795;
srom_1(95470) <= 321471;
srom_1(95471) <= 182976;
srom_1(95472) <= 82960;
srom_1(95473) <= 21892;
srom_1(95474) <= 59;
srom_1(95475) <= 17563;
srom_1(95476) <= 74321;
srom_1(95477) <= 170067;
srom_1(95478) <= 304354;
srom_1(95479) <= 476550;
srom_1(95480) <= 685848;
srom_1(95481) <= 931267;
srom_1(95482) <= 1211657;
srom_1(95483) <= 1525701;
srom_1(95484) <= 1871928;
srom_1(95485) <= 2248714;
srom_1(95486) <= 2654292;
srom_1(95487) <= 3086761;
srom_1(95488) <= 3544091;
srom_1(95489) <= 4024139;
srom_1(95490) <= 4524654;
srom_1(95491) <= 5043287;
srom_1(95492) <= 5577609;
srom_1(95493) <= 6125112;
srom_1(95494) <= 6683229;
srom_1(95495) <= 7249343;
srom_1(95496) <= 7820800;
srom_1(95497) <= 8394919;
srom_1(95498) <= 8969009;
srom_1(95499) <= 9540377;
srom_1(95500) <= 10106344;
srom_1(95501) <= 10664256;
srom_1(95502) <= 11211497;
srom_1(95503) <= 11745500;
srom_1(95504) <= 12263762;
srom_1(95505) <= 12763851;
srom_1(95506) <= 13243424;
srom_1(95507) <= 13700231;
srom_1(95508) <= 14132129;
srom_1(95509) <= 14537095;
srom_1(95510) <= 14913228;
srom_1(95511) <= 15258764;
srom_1(95512) <= 15572084;
srom_1(95513) <= 15851719;
srom_1(95514) <= 16096356;
srom_1(95515) <= 16304849;
srom_1(95516) <= 16476220;
srom_1(95517) <= 16609666;
srom_1(95518) <= 16704560;
srom_1(95519) <= 16760458;
srom_1(95520) <= 16777097;
srom_1(95521) <= 16754399;
srom_1(95522) <= 16692472;
srom_1(95523) <= 16591605;
srom_1(95524) <= 16452271;
srom_1(95525) <= 16275124;
srom_1(95526) <= 16060995;
srom_1(95527) <= 15810887;
srom_1(95528) <= 15525973;
srom_1(95529) <= 15207590;
srom_1(95530) <= 14857230;
srom_1(95531) <= 14476536;
srom_1(95532) <= 14067295;
srom_1(95533) <= 13631424;
srom_1(95534) <= 13170967;
srom_1(95535) <= 12688084;
srom_1(95536) <= 12185040;
srom_1(95537) <= 11664193;
srom_1(95538) <= 11127985;
srom_1(95539) <= 10578932;
srom_1(95540) <= 10019608;
srom_1(95541) <= 9452635;
srom_1(95542) <= 8880672;
srom_1(95543) <= 8306402;
srom_1(95544) <= 7732518;
srom_1(95545) <= 7161710;
srom_1(95546) <= 6596655;
srom_1(95547) <= 6040004;
srom_1(95548) <= 5494366;
srom_1(95549) <= 4962300;
srom_1(95550) <= 4446301;
srom_1(95551) <= 3948789;
srom_1(95552) <= 3472097;
srom_1(95553) <= 3018460;
srom_1(95554) <= 2590006;
srom_1(95555) <= 2188743;
srom_1(95556) <= 1816553;
srom_1(95557) <= 1475182;
srom_1(95558) <= 1166231;
srom_1(95559) <= 891147;
srom_1(95560) <= 651222;
srom_1(95561) <= 447580;
srom_1(95562) <= 281177;
srom_1(95563) <= 152791;
srom_1(95564) <= 63027;
srom_1(95565) <= 12304;
srom_1(95566) <= 860;
srom_1(95567) <= 28749;
srom_1(95568) <= 95841;
srom_1(95569) <= 201820;
srom_1(95570) <= 346190;
srom_1(95571) <= 528273;
srom_1(95572) <= 747216;
srom_1(95573) <= 1001993;
srom_1(95574) <= 1291407;
srom_1(95575) <= 1614103;
srom_1(95576) <= 1968567;
srom_1(95577) <= 2353137;
srom_1(95578) <= 2766009;
srom_1(95579) <= 3205247;
srom_1(95580) <= 3668792;
srom_1(95581) <= 4154470;
srom_1(95582) <= 4660003;
srom_1(95583) <= 5183021;
srom_1(95584) <= 5721071;
srom_1(95585) <= 6271630;
srom_1(95586) <= 6832116;
srom_1(95587) <= 7399901;
srom_1(95588) <= 7972322;
srom_1(95589) <= 8546695;
srom_1(95590) <= 9120328;
srom_1(95591) <= 9690528;
srom_1(95592) <= 10254624;
srom_1(95593) <= 10809969;
srom_1(95594) <= 11353960;
srom_1(95595) <= 11884045;
srom_1(95596) <= 12397739;
srom_1(95597) <= 12892633;
srom_1(95598) <= 13366405;
srom_1(95599) <= 13816836;
srom_1(95600) <= 14241811;
srom_1(95601) <= 14639338;
srom_1(95602) <= 15007554;
srom_1(95603) <= 15344731;
srom_1(95604) <= 15649289;
srom_1(95605) <= 15919799;
srom_1(95606) <= 16154992;
srom_1(95607) <= 16353766;
srom_1(95608) <= 16515189;
srom_1(95609) <= 16638503;
srom_1(95610) <= 16723131;
srom_1(95611) <= 16768675;
srom_1(95612) <= 16774923;
srom_1(95613) <= 16741844;
srom_1(95614) <= 16669594;
srom_1(95615) <= 16558511;
srom_1(95616) <= 16409117;
srom_1(95617) <= 16222112;
srom_1(95618) <= 15998373;
srom_1(95619) <= 15738949;
srom_1(95620) <= 15445057;
srom_1(95621) <= 15118075;
srom_1(95622) <= 14759536;
srom_1(95623) <= 14371122;
srom_1(95624) <= 13954653;
srom_1(95625) <= 13512083;
srom_1(95626) <= 13045488;
srom_1(95627) <= 12557055;
srom_1(95628) <= 12049075;
srom_1(95629) <= 11523929;
srom_1(95630) <= 10984081;
srom_1(95631) <= 10432062;
srom_1(95632) <= 9870460;
srom_1(95633) <= 9301909;
srom_1(95634) <= 8729076;
srom_1(95635) <= 8154646;
srom_1(95636) <= 7581313;
srom_1(95637) <= 7011766;
srom_1(95638) <= 6448675;
srom_1(95639) <= 5894681;
srom_1(95640) <= 5352382;
srom_1(95641) <= 4824321;
srom_1(95642) <= 4312975;
srom_1(95643) <= 3820740;
srom_1(95644) <= 3349925;
srom_1(95645) <= 2902739;
srom_1(95646) <= 2481278;
srom_1(95647) <= 2087518;
srom_1(95648) <= 1723306;
srom_1(95649) <= 1390351;
srom_1(95650) <= 1090212;
srom_1(95651) <= 824298;
srom_1(95652) <= 593856;
srom_1(95653) <= 399965;
srom_1(95654) <= 243537;
srom_1(95655) <= 125303;
srom_1(95656) <= 45819;
srom_1(95657) <= 5457;
srom_1(95658) <= 4407;
srom_1(95659) <= 42673;
srom_1(95660) <= 120076;
srom_1(95661) <= 236253;
srom_1(95662) <= 390659;
srom_1(95663) <= 582570;
srom_1(95664) <= 811086;
srom_1(95665) <= 1075136;
srom_1(95666) <= 1373482;
srom_1(95667) <= 1704723;
srom_1(95668) <= 2067308;
srom_1(95669) <= 2459536;
srom_1(95670) <= 2879566;
srom_1(95671) <= 3325431;
srom_1(95672) <= 3795039;
srom_1(95673) <= 4286187;
srom_1(95674) <= 4796573;
srom_1(95675) <= 5323804;
srom_1(95676) <= 5865406;
srom_1(95677) <= 6418841;
srom_1(95678) <= 6981512;
srom_1(95679) <= 7550782;
srom_1(95680) <= 8123980;
srom_1(95681) <= 8698420;
srom_1(95682) <= 9271406;
srom_1(95683) <= 9840253;
srom_1(95684) <= 10402293;
srom_1(95685) <= 10954890;
srom_1(95686) <= 11495452;
srom_1(95687) <= 12021446;
srom_1(95688) <= 12530404;
srom_1(95689) <= 13019939;
srom_1(95690) <= 13487757;
srom_1(95691) <= 13931663;
srom_1(95692) <= 14349576;
srom_1(95693) <= 14739536;
srom_1(95694) <= 15099714;
srom_1(95695) <= 15428421;
srom_1(95696) <= 15724116;
srom_1(95697) <= 15985413;
srom_1(95698) <= 16211085;
srom_1(95699) <= 16400075;
srom_1(95700) <= 16551497;
srom_1(95701) <= 16664640;
srom_1(95702) <= 16738974;
srom_1(95703) <= 16774150;
srom_1(95704) <= 16770003;
srom_1(95705) <= 16726553;
srom_1(95706) <= 16644004;
srom_1(95707) <= 16522742;
srom_1(95708) <= 16363337;
srom_1(95709) <= 16166535;
srom_1(95710) <= 15933260;
srom_1(95711) <= 15664605;
srom_1(95712) <= 15361831;
srom_1(95713) <= 15026357;
srom_1(95714) <= 14659756;
srom_1(95715) <= 14263748;
srom_1(95716) <= 13840189;
srom_1(95717) <= 13391066;
srom_1(95718) <= 12918484;
srom_1(95719) <= 12424661;
srom_1(95720) <= 11911911;
srom_1(95721) <= 11382639;
srom_1(95722) <= 10839326;
srom_1(95723) <= 10284522;
srom_1(95724) <= 9720827;
srom_1(95725) <= 9150885;
srom_1(95726) <= 8577368;
srom_1(95727) <= 8002966;
srom_1(95728) <= 7430372;
srom_1(95729) <= 6862272;
srom_1(95730) <= 6301330;
srom_1(95731) <= 5750175;
srom_1(95732) <= 5211393;
srom_1(95733) <= 4687510;
srom_1(95734) <= 4180983;
srom_1(95735) <= 3694186;
srom_1(95736) <= 3229404;
srom_1(95737) <= 2788814;
srom_1(95738) <= 2374484;
srom_1(95739) <= 1988356;
srom_1(95740) <= 1632242;
srom_1(95741) <= 1307810;
srom_1(95742) <= 1016582;
srom_1(95743) <= 759925;
srom_1(95744) <= 539041;
srom_1(95745) <= 354966;
srom_1(95746) <= 208564;
srom_1(95747) <= 100520;
srom_1(95748) <= 31343;
srom_1(95749) <= 1355;
srom_1(95750) <= 10699;
srom_1(95751) <= 59329;
srom_1(95752) <= 147018;
srom_1(95753) <= 273354;
srom_1(95754) <= 437746;
srom_1(95755) <= 639422;
srom_1(95756) <= 877437;
srom_1(95757) <= 1150674;
srom_1(95758) <= 1457853;
srom_1(95759) <= 1797532;
srom_1(95760) <= 2168118;
srom_1(95761) <= 2567875;
srom_1(95762) <= 2994927;
srom_1(95763) <= 3447273;
srom_1(95764) <= 3922789;
srom_1(95765) <= 4419248;
srom_1(95766) <= 4934320;
srom_1(95767) <= 5465590;
srom_1(95768) <= 6010568;
srom_1(95769) <= 6566697;
srom_1(95770) <= 7131369;
srom_1(95771) <= 7701937;
srom_1(95772) <= 8275725;
srom_1(95773) <= 8850043;
srom_1(95774) <= 9422196;
srom_1(95775) <= 9989503;
srom_1(95776) <= 10549303;
srom_1(95777) <= 11098970;
srom_1(95778) <= 11635928;
srom_1(95779) <= 12157657;
srom_1(95780) <= 12661713;
srom_1(95781) <= 13145730;
srom_1(95782) <= 13607440;
srom_1(95783) <= 14044676;
srom_1(95784) <= 14455389;
srom_1(95785) <= 14837654;
srom_1(95786) <= 15189676;
srom_1(95787) <= 15509806;
srom_1(95788) <= 15796542;
srom_1(95789) <= 16048539;
srom_1(95790) <= 16264617;
srom_1(95791) <= 16443761;
srom_1(95792) <= 16585132;
srom_1(95793) <= 16688067;
srom_1(95794) <= 16752082;
srom_1(95795) <= 16776879;
srom_1(95796) <= 16762340;
srom_1(95797) <= 16708533;
srom_1(95798) <= 16615712;
srom_1(95799) <= 16484311;
srom_1(95800) <= 16314946;
srom_1(95801) <= 16108412;
srom_1(95802) <= 15865677;
srom_1(95803) <= 15587880;
srom_1(95804) <= 15276322;
srom_1(95805) <= 14932466;
srom_1(95806) <= 14557924;
srom_1(95807) <= 14154451;
srom_1(95808) <= 13723940;
srom_1(95809) <= 13268411;
srom_1(95810) <= 12789998;
srom_1(95811) <= 12290945;
srom_1(95812) <= 11773593;
srom_1(95813) <= 11240368;
srom_1(95814) <= 10693770;
srom_1(95815) <= 10136362;
srom_1(95816) <= 9570758;
srom_1(95817) <= 8999611;
srom_1(95818) <= 8425598;
srom_1(95819) <= 7851412;
srom_1(95820) <= 7279746;
srom_1(95821) <= 6713279;
srom_1(95822) <= 6154668;
srom_1(95823) <= 5606533;
srom_1(95824) <= 5071444;
srom_1(95825) <= 4551910;
srom_1(95826) <= 4050368;
srom_1(95827) <= 3569169;
srom_1(95828) <= 3110571;
srom_1(95829) <= 2676723;
srom_1(95830) <= 2269659;
srom_1(95831) <= 1891290;
srom_1(95832) <= 1543389;
srom_1(95833) <= 1227588;
srom_1(95834) <= 945366;
srom_1(95835) <= 698049;
srom_1(95836) <= 486796;
srom_1(95837) <= 312597;
srom_1(95838) <= 176269;
srom_1(95839) <= 78451;
srom_1(95840) <= 19603;
srom_1(95841) <= 0;
srom_1(95842) <= 19733;
srom_1(95843) <= 78712;
srom_1(95844) <= 176658;
srom_1(95845) <= 313113;
srom_1(95846) <= 487437;
srom_1(95847) <= 698812;
srom_1(95848) <= 946247;
srom_1(95849) <= 1228582;
srom_1(95850) <= 1544493;
srom_1(95851) <= 1892498;
srom_1(95852) <= 2270965;
srom_1(95853) <= 2678121;
srom_1(95854) <= 3112054;
srom_1(95855) <= 3570732;
srom_1(95856) <= 4052002;
srom_1(95857) <= 4553607;
srom_1(95858) <= 5073197;
srom_1(95859) <= 5608333;
srom_1(95860) <= 6156508;
srom_1(95861) <= 6715149;
srom_1(95862) <= 7281638;
srom_1(95863) <= 7853317;
srom_1(95864) <= 8427507;
srom_1(95865) <= 9001514;
srom_1(95866) <= 9572648;
srom_1(95867) <= 10138229;
srom_1(95868) <= 10695605;
srom_1(95869) <= 11242163;
srom_1(95870) <= 11775340;
srom_1(95871) <= 12292635;
srom_1(95872) <= 12791623;
srom_1(95873) <= 13269963;
srom_1(95874) <= 13725413;
srom_1(95875) <= 14155837;
srom_1(95876) <= 14559217;
srom_1(95877) <= 14933660;
srom_1(95878) <= 15277412;
srom_1(95879) <= 15588859;
srom_1(95880) <= 15866542;
srom_1(95881) <= 16109159;
srom_1(95882) <= 16315571;
srom_1(95883) <= 16484810;
srom_1(95884) <= 16616084;
srom_1(95885) <= 16708777;
srom_1(95886) <= 16762453;
srom_1(95887) <= 16776862;
srom_1(95888) <= 16751935;
srom_1(95889) <= 16687789;
srom_1(95890) <= 16584726;
srom_1(95891) <= 16443228;
srom_1(95892) <= 16263960;
srom_1(95893) <= 16047761;
srom_1(95894) <= 15795646;
srom_1(95895) <= 15508797;
srom_1(95896) <= 15188558;
srom_1(95897) <= 14836433;
srom_1(95898) <= 14454071;
srom_1(95899) <= 14043266;
srom_1(95900) <= 13605945;
srom_1(95901) <= 13144158;
srom_1(95902) <= 12660070;
srom_1(95903) <= 12155952;
srom_1(95904) <= 11634168;
srom_1(95905) <= 11097164;
srom_1(95906) <= 10547458;
srom_1(95907) <= 9987629;
srom_1(95908) <= 9420302;
srom_1(95909) <= 8848137;
srom_1(95910) <= 8273817;
srom_1(95911) <= 7700035;
srom_1(95912) <= 7129482;
srom_1(95913) <= 6564833;
srom_1(95914) <= 6008737;
srom_1(95915) <= 5463801;
srom_1(95916) <= 4932580;
srom_1(95917) <= 4417566;
srom_1(95918) <= 3921174;
srom_1(95919) <= 3445730;
srom_1(95920) <= 2993466;
srom_1(95921) <= 2566501;
srom_1(95922) <= 2166838;
srom_1(95923) <= 1796351;
srom_1(95924) <= 1456777;
srom_1(95925) <= 1149710;
srom_1(95926) <= 876587;
srom_1(95927) <= 638692;
srom_1(95928) <= 437138;
srom_1(95929) <= 272871;
srom_1(95930) <= 146662;
srom_1(95931) <= 59102;
srom_1(95932) <= 10603;
srom_1(95933) <= 1390;
srom_1(95934) <= 31508;
srom_1(95935) <= 100815;
srom_1(95936) <= 208987;
srom_1(95937) <= 355516;
srom_1(95938) <= 539714;
srom_1(95939) <= 760719;
srom_1(95940) <= 1017493;
srom_1(95941) <= 1308834;
srom_1(95942) <= 1633373;
srom_1(95943) <= 1989591;
srom_1(95944) <= 2375815;
srom_1(95945) <= 2790236;
srom_1(95946) <= 3230909;
srom_1(95947) <= 3695768;
srom_1(95948) <= 4182634;
srom_1(95949) <= 4689223;
srom_1(95950) <= 5213160;
srom_1(95951) <= 5751987;
srom_1(95952) <= 6303178;
srom_1(95953) <= 6864149;
srom_1(95954) <= 7432269;
srom_1(95955) <= 8004873;
srom_1(95956) <= 8579276;
srom_1(95957) <= 9152786;
srom_1(95958) <= 9722712;
srom_1(95959) <= 10286381;
srom_1(95960) <= 10841152;
srom_1(95961) <= 11384422;
srom_1(95962) <= 11913643;
srom_1(95963) <= 12426334;
srom_1(95964) <= 12920091;
srom_1(95965) <= 13392598;
srom_1(95966) <= 13841640;
srom_1(95967) <= 14265110;
srom_1(95968) <= 14661024;
srom_1(95969) <= 15027524;
srom_1(95970) <= 15362892;
srom_1(95971) <= 15665555;
srom_1(95972) <= 15934094;
srom_1(95973) <= 16167250;
srom_1(95974) <= 16363929;
srom_1(95975) <= 16523209;
srom_1(95976) <= 16644343;
srom_1(95977) <= 16726763;
srom_1(95978) <= 16770082;
srom_1(95979) <= 16774098;
srom_1(95980) <= 16738791;
srom_1(95981) <= 16664328;
srom_1(95982) <= 16551057;
srom_1(95983) <= 16399509;
srom_1(95984) <= 16210395;
srom_1(95985) <= 15984603;
srom_1(95986) <= 15723190;
srom_1(95987) <= 15427383;
srom_1(95988) <= 15098568;
srom_1(95989) <= 14738288;
srom_1(95990) <= 14348233;
srom_1(95991) <= 13930230;
srom_1(95992) <= 13486241;
srom_1(95993) <= 13018348;
srom_1(95994) <= 12528744;
srom_1(95995) <= 12019725;
srom_1(95996) <= 11493679;
srom_1(95997) <= 10953073;
srom_1(95998) <= 10400440;
srom_1(95999) <= 9838373;
srom_1(96000) <= 9269508;
srom_1(96001) <= 8696512;
end Behavioral;